magic
tech sky130A
magscale 1 2
timestamp 1625507855
<< obsli1 >>
rect 1104 2159 153916 155057
<< obsm1 >>
rect 474 8 154270 156732
<< metal2 >>
rect 1398 156455 1454 157255
rect 2778 156455 2834 157255
rect 4158 156455 4214 157255
rect 5078 156455 5134 157255
rect 6458 156455 6514 157255
rect 7838 156455 7894 157255
rect 9218 156455 9274 157255
rect 10138 156455 10194 157255
rect 11518 156455 11574 157255
rect 12898 156455 12954 157255
rect 14278 156455 14334 157255
rect 15198 156455 15254 157255
rect 16578 156455 16634 157255
rect 17958 156455 18014 157255
rect 19338 156455 19394 157255
rect 20718 156455 20774 157255
rect 21638 156455 21694 157255
rect 23018 156455 23074 157255
rect 24398 156455 24454 157255
rect 25778 156455 25834 157255
rect 26698 156455 26754 157255
rect 28078 156455 28134 157255
rect 29458 156455 29514 157255
rect 30838 156455 30894 157255
rect 31758 156455 31814 157255
rect 33138 156455 33194 157255
rect 34518 156455 34574 157255
rect 35898 156455 35954 157255
rect 36818 156455 36874 157255
rect 38198 156455 38254 157255
rect 39578 156455 39634 157255
rect 40958 156455 41014 157255
rect 42338 156455 42394 157255
rect 43258 156455 43314 157255
rect 44638 156455 44694 157255
rect 46018 156455 46074 157255
rect 47398 156455 47454 157255
rect 48318 156455 48374 157255
rect 49698 156455 49754 157255
rect 51078 156455 51134 157255
rect 52458 156455 52514 157255
rect 53378 156455 53434 157255
rect 54758 156455 54814 157255
rect 56138 156455 56194 157255
rect 57518 156455 57574 157255
rect 58898 156455 58954 157255
rect 59818 156455 59874 157255
rect 61198 156455 61254 157255
rect 62578 156455 62634 157255
rect 63958 156455 64014 157255
rect 64878 156455 64934 157255
rect 66258 156455 66314 157255
rect 67638 156455 67694 157255
rect 69018 156455 69074 157255
rect 69938 156455 69994 157255
rect 71318 156455 71374 157255
rect 72698 156455 72754 157255
rect 74078 156455 74134 157255
rect 75458 156455 75514 157255
rect 76378 156455 76434 157255
rect 77758 156455 77814 157255
rect 79138 156455 79194 157255
rect 80518 156455 80574 157255
rect 81438 156455 81494 157255
rect 82818 156455 82874 157255
rect 84198 156455 84254 157255
rect 85578 156455 85634 157255
rect 86498 156455 86554 157255
rect 87878 156455 87934 157255
rect 89258 156455 89314 157255
rect 90638 156455 90694 157255
rect 91558 156455 91614 157255
rect 92938 156455 92994 157255
rect 94318 156455 94374 157255
rect 95698 156455 95754 157255
rect 97078 156455 97134 157255
rect 97998 156455 98054 157255
rect 99378 156455 99434 157255
rect 100758 156455 100814 157255
rect 102138 156455 102194 157255
rect 103058 156455 103114 157255
rect 104438 156455 104494 157255
rect 105818 156455 105874 157255
rect 107198 156455 107254 157255
rect 108118 156455 108174 157255
rect 109498 156455 109554 157255
rect 110878 156455 110934 157255
rect 112258 156455 112314 157255
rect 113638 156455 113694 157255
rect 114558 156455 114614 157255
rect 115938 156455 115994 157255
rect 117318 156455 117374 157255
rect 118698 156455 118754 157255
rect 119618 156455 119674 157255
rect 120998 156455 121054 157255
rect 122378 156455 122434 157255
rect 123758 156455 123814 157255
rect 124678 156455 124734 157255
rect 126058 156455 126114 157255
rect 127438 156455 127494 157255
rect 128818 156455 128874 157255
rect 130198 156455 130254 157255
rect 131118 156455 131174 157255
rect 132498 156455 132554 157255
rect 133878 156455 133934 157255
rect 135258 156455 135314 157255
rect 136178 156455 136234 157255
rect 137558 156455 137614 157255
rect 138938 156455 138994 157255
rect 140318 156455 140374 157255
rect 141238 156455 141294 157255
rect 142618 156455 142674 157255
rect 143998 156455 144054 157255
rect 145378 156455 145434 157255
rect 146758 156455 146814 157255
rect 147678 156455 147734 157255
rect 149058 156455 149114 157255
rect 150438 156455 150494 157255
rect 151818 156455 151874 157255
rect 152738 156455 152794 157255
rect 154118 156455 154174 157255
rect 478 0 534 800
rect 1398 0 1454 800
rect 2778 0 2834 800
rect 4158 0 4214 800
rect 5538 0 5594 800
rect 6458 0 6514 800
rect 7838 0 7894 800
rect 9218 0 9274 800
rect 10598 0 10654 800
rect 11518 0 11574 800
rect 12898 0 12954 800
rect 14278 0 14334 800
rect 15658 0 15714 800
rect 16578 0 16634 800
rect 17958 0 18014 800
rect 19338 0 19394 800
rect 20718 0 20774 800
rect 22098 0 22154 800
rect 23018 0 23074 800
rect 24398 0 24454 800
rect 25778 0 25834 800
rect 27158 0 27214 800
rect 28078 0 28134 800
rect 29458 0 29514 800
rect 30838 0 30894 800
rect 32218 0 32274 800
rect 33138 0 33194 800
rect 34518 0 34574 800
rect 35898 0 35954 800
rect 37278 0 37334 800
rect 38658 0 38714 800
rect 39578 0 39634 800
rect 40958 0 41014 800
rect 42338 0 42394 800
rect 43718 0 43774 800
rect 44638 0 44694 800
rect 46018 0 46074 800
rect 47398 0 47454 800
rect 48778 0 48834 800
rect 49698 0 49754 800
rect 51078 0 51134 800
rect 52458 0 52514 800
rect 53838 0 53894 800
rect 55218 0 55274 800
rect 56138 0 56194 800
rect 57518 0 57574 800
rect 58898 0 58954 800
rect 60278 0 60334 800
rect 61198 0 61254 800
rect 62578 0 62634 800
rect 63958 0 64014 800
rect 65338 0 65394 800
rect 66258 0 66314 800
rect 67638 0 67694 800
rect 69018 0 69074 800
rect 70398 0 70454 800
rect 71318 0 71374 800
rect 72698 0 72754 800
rect 74078 0 74134 800
rect 75458 0 75514 800
rect 76838 0 76894 800
rect 77758 0 77814 800
rect 79138 0 79194 800
rect 80518 0 80574 800
rect 81898 0 81954 800
rect 82818 0 82874 800
rect 84198 0 84254 800
rect 85578 0 85634 800
rect 86958 0 87014 800
rect 87878 0 87934 800
rect 89258 0 89314 800
rect 90638 0 90694 800
rect 92018 0 92074 800
rect 93398 0 93454 800
rect 94318 0 94374 800
rect 95698 0 95754 800
rect 97078 0 97134 800
rect 98458 0 98514 800
rect 99378 0 99434 800
rect 100758 0 100814 800
rect 102138 0 102194 800
rect 103518 0 103574 800
rect 104438 0 104494 800
rect 105818 0 105874 800
rect 107198 0 107254 800
rect 108578 0 108634 800
rect 109958 0 110014 800
rect 110878 0 110934 800
rect 112258 0 112314 800
rect 113638 0 113694 800
rect 115018 0 115074 800
rect 115938 0 115994 800
rect 117318 0 117374 800
rect 118698 0 118754 800
rect 120078 0 120134 800
rect 120998 0 121054 800
rect 122378 0 122434 800
rect 123758 0 123814 800
rect 125138 0 125194 800
rect 126518 0 126574 800
rect 127438 0 127494 800
rect 128818 0 128874 800
rect 130198 0 130254 800
rect 131578 0 131634 800
rect 132498 0 132554 800
rect 133878 0 133934 800
rect 135258 0 135314 800
rect 136638 0 136694 800
rect 137558 0 137614 800
rect 138938 0 138994 800
rect 140318 0 140374 800
rect 141698 0 141754 800
rect 142618 0 142674 800
rect 143998 0 144054 800
rect 145378 0 145434 800
rect 146758 0 146814 800
rect 148138 0 148194 800
rect 149058 0 149114 800
rect 150438 0 150494 800
rect 151818 0 151874 800
rect 153198 0 153254 800
rect 154118 0 154174 800
<< obsm2 >>
rect 480 156399 1342 156738
rect 1510 156399 2722 156738
rect 2890 156399 4102 156738
rect 4270 156399 5022 156738
rect 5190 156399 6402 156738
rect 6570 156399 7782 156738
rect 7950 156399 9162 156738
rect 9330 156399 10082 156738
rect 10250 156399 11462 156738
rect 11630 156399 12842 156738
rect 13010 156399 14222 156738
rect 14390 156399 15142 156738
rect 15310 156399 16522 156738
rect 16690 156399 17902 156738
rect 18070 156399 19282 156738
rect 19450 156399 20662 156738
rect 20830 156399 21582 156738
rect 21750 156399 22962 156738
rect 23130 156399 24342 156738
rect 24510 156399 25722 156738
rect 25890 156399 26642 156738
rect 26810 156399 28022 156738
rect 28190 156399 29402 156738
rect 29570 156399 30782 156738
rect 30950 156399 31702 156738
rect 31870 156399 33082 156738
rect 33250 156399 34462 156738
rect 34630 156399 35842 156738
rect 36010 156399 36762 156738
rect 36930 156399 38142 156738
rect 38310 156399 39522 156738
rect 39690 156399 40902 156738
rect 41070 156399 42282 156738
rect 42450 156399 43202 156738
rect 43370 156399 44582 156738
rect 44750 156399 45962 156738
rect 46130 156399 47342 156738
rect 47510 156399 48262 156738
rect 48430 156399 49642 156738
rect 49810 156399 51022 156738
rect 51190 156399 52402 156738
rect 52570 156399 53322 156738
rect 53490 156399 54702 156738
rect 54870 156399 56082 156738
rect 56250 156399 57462 156738
rect 57630 156399 58842 156738
rect 59010 156399 59762 156738
rect 59930 156399 61142 156738
rect 61310 156399 62522 156738
rect 62690 156399 63902 156738
rect 64070 156399 64822 156738
rect 64990 156399 66202 156738
rect 66370 156399 67582 156738
rect 67750 156399 68962 156738
rect 69130 156399 69882 156738
rect 70050 156399 71262 156738
rect 71430 156399 72642 156738
rect 72810 156399 74022 156738
rect 74190 156399 75402 156738
rect 75570 156399 76322 156738
rect 76490 156399 77702 156738
rect 77870 156399 79082 156738
rect 79250 156399 80462 156738
rect 80630 156399 81382 156738
rect 81550 156399 82762 156738
rect 82930 156399 84142 156738
rect 84310 156399 85522 156738
rect 85690 156399 86442 156738
rect 86610 156399 87822 156738
rect 87990 156399 89202 156738
rect 89370 156399 90582 156738
rect 90750 156399 91502 156738
rect 91670 156399 92882 156738
rect 93050 156399 94262 156738
rect 94430 156399 95642 156738
rect 95810 156399 97022 156738
rect 97190 156399 97942 156738
rect 98110 156399 99322 156738
rect 99490 156399 100702 156738
rect 100870 156399 102082 156738
rect 102250 156399 103002 156738
rect 103170 156399 104382 156738
rect 104550 156399 105762 156738
rect 105930 156399 107142 156738
rect 107310 156399 108062 156738
rect 108230 156399 109442 156738
rect 109610 156399 110822 156738
rect 110990 156399 112202 156738
rect 112370 156399 113582 156738
rect 113750 156399 114502 156738
rect 114670 156399 115882 156738
rect 116050 156399 117262 156738
rect 117430 156399 118642 156738
rect 118810 156399 119562 156738
rect 119730 156399 120942 156738
rect 121110 156399 122322 156738
rect 122490 156399 123702 156738
rect 123870 156399 124622 156738
rect 124790 156399 126002 156738
rect 126170 156399 127382 156738
rect 127550 156399 128762 156738
rect 128930 156399 130142 156738
rect 130310 156399 131062 156738
rect 131230 156399 132442 156738
rect 132610 156399 133822 156738
rect 133990 156399 135202 156738
rect 135370 156399 136122 156738
rect 136290 156399 137502 156738
rect 137670 156399 138882 156738
rect 139050 156399 140262 156738
rect 140430 156399 141182 156738
rect 141350 156399 142562 156738
rect 142730 156399 143942 156738
rect 144110 156399 145322 156738
rect 145490 156399 146702 156738
rect 146870 156399 147622 156738
rect 147790 156399 149002 156738
rect 149170 156399 150382 156738
rect 150550 156399 151762 156738
rect 151930 156399 152682 156738
rect 152850 156399 154062 156738
rect 154230 156399 154264 156738
rect 480 856 154264 156399
rect 590 2 1342 856
rect 1510 2 2722 856
rect 2890 2 4102 856
rect 4270 2 5482 856
rect 5650 2 6402 856
rect 6570 2 7782 856
rect 7950 2 9162 856
rect 9330 2 10542 856
rect 10710 2 11462 856
rect 11630 2 12842 856
rect 13010 2 14222 856
rect 14390 2 15602 856
rect 15770 2 16522 856
rect 16690 2 17902 856
rect 18070 2 19282 856
rect 19450 2 20662 856
rect 20830 2 22042 856
rect 22210 2 22962 856
rect 23130 2 24342 856
rect 24510 2 25722 856
rect 25890 2 27102 856
rect 27270 2 28022 856
rect 28190 2 29402 856
rect 29570 2 30782 856
rect 30950 2 32162 856
rect 32330 2 33082 856
rect 33250 2 34462 856
rect 34630 2 35842 856
rect 36010 2 37222 856
rect 37390 2 38602 856
rect 38770 2 39522 856
rect 39690 2 40902 856
rect 41070 2 42282 856
rect 42450 2 43662 856
rect 43830 2 44582 856
rect 44750 2 45962 856
rect 46130 2 47342 856
rect 47510 2 48722 856
rect 48890 2 49642 856
rect 49810 2 51022 856
rect 51190 2 52402 856
rect 52570 2 53782 856
rect 53950 2 55162 856
rect 55330 2 56082 856
rect 56250 2 57462 856
rect 57630 2 58842 856
rect 59010 2 60222 856
rect 60390 2 61142 856
rect 61310 2 62522 856
rect 62690 2 63902 856
rect 64070 2 65282 856
rect 65450 2 66202 856
rect 66370 2 67582 856
rect 67750 2 68962 856
rect 69130 2 70342 856
rect 70510 2 71262 856
rect 71430 2 72642 856
rect 72810 2 74022 856
rect 74190 2 75402 856
rect 75570 2 76782 856
rect 76950 2 77702 856
rect 77870 2 79082 856
rect 79250 2 80462 856
rect 80630 2 81842 856
rect 82010 2 82762 856
rect 82930 2 84142 856
rect 84310 2 85522 856
rect 85690 2 86902 856
rect 87070 2 87822 856
rect 87990 2 89202 856
rect 89370 2 90582 856
rect 90750 2 91962 856
rect 92130 2 93342 856
rect 93510 2 94262 856
rect 94430 2 95642 856
rect 95810 2 97022 856
rect 97190 2 98402 856
rect 98570 2 99322 856
rect 99490 2 100702 856
rect 100870 2 102082 856
rect 102250 2 103462 856
rect 103630 2 104382 856
rect 104550 2 105762 856
rect 105930 2 107142 856
rect 107310 2 108522 856
rect 108690 2 109902 856
rect 110070 2 110822 856
rect 110990 2 112202 856
rect 112370 2 113582 856
rect 113750 2 114962 856
rect 115130 2 115882 856
rect 116050 2 117262 856
rect 117430 2 118642 856
rect 118810 2 120022 856
rect 120190 2 120942 856
rect 121110 2 122322 856
rect 122490 2 123702 856
rect 123870 2 125082 856
rect 125250 2 126462 856
rect 126630 2 127382 856
rect 127550 2 128762 856
rect 128930 2 130142 856
rect 130310 2 131522 856
rect 131690 2 132442 856
rect 132610 2 133822 856
rect 133990 2 135202 856
rect 135370 2 136582 856
rect 136750 2 137502 856
rect 137670 2 138882 856
rect 139050 2 140262 856
rect 140430 2 141642 856
rect 141810 2 142562 856
rect 142730 2 143942 856
rect 144110 2 145322 856
rect 145490 2 146702 856
rect 146870 2 148082 856
rect 148250 2 149002 856
rect 149170 2 150382 856
rect 150550 2 151762 856
rect 151930 2 153142 856
rect 153310 2 154062 856
rect 154230 2 154264 856
<< metal3 >>
rect 0 156408 800 156528
rect 154311 155728 155111 155848
rect 0 154368 800 154488
rect 154311 153688 155111 153808
rect 0 153008 800 153128
rect 154311 152328 155111 152448
rect 0 150968 800 151088
rect 154311 150288 155111 150408
rect 0 148928 800 149048
rect 154311 148248 155111 148368
rect 0 146888 800 147008
rect 154311 146208 155111 146328
rect 0 145528 800 145648
rect 154311 144848 155111 144968
rect 0 143488 800 143608
rect 154311 142808 155111 142928
rect 0 141448 800 141568
rect 154311 140768 155111 140888
rect 0 139408 800 139528
rect 154311 138728 155111 138848
rect 0 138048 800 138168
rect 154311 136688 155111 136808
rect 0 136008 800 136128
rect 154311 135328 155111 135448
rect 0 133968 800 134088
rect 154311 133288 155111 133408
rect 0 131928 800 132048
rect 154311 131248 155111 131368
rect 0 129888 800 130008
rect 154311 129208 155111 129328
rect 0 128528 800 128648
rect 154311 127848 155111 127968
rect 0 126488 800 126608
rect 154311 125808 155111 125928
rect 0 124448 800 124568
rect 154311 123768 155111 123888
rect 0 122408 800 122528
rect 154311 121728 155111 121848
rect 0 121048 800 121168
rect 154311 120368 155111 120488
rect 0 119008 800 119128
rect 154311 118328 155111 118448
rect 0 116968 800 117088
rect 154311 116288 155111 116408
rect 0 114928 800 115048
rect 154311 114248 155111 114368
rect 0 113568 800 113688
rect 154311 112208 155111 112328
rect 0 111528 800 111648
rect 154311 110848 155111 110968
rect 0 109488 800 109608
rect 154311 108808 155111 108928
rect 0 107448 800 107568
rect 154311 106768 155111 106888
rect 0 105408 800 105528
rect 154311 104728 155111 104848
rect 0 104048 800 104168
rect 154311 103368 155111 103488
rect 0 102008 800 102128
rect 154311 101328 155111 101448
rect 0 99968 800 100088
rect 154311 99288 155111 99408
rect 0 97928 800 98048
rect 154311 97248 155111 97368
rect 0 96568 800 96688
rect 154311 95888 155111 96008
rect 0 94528 800 94648
rect 154311 93848 155111 93968
rect 0 92488 800 92608
rect 154311 91808 155111 91928
rect 0 90448 800 90568
rect 154311 89768 155111 89888
rect 0 89088 800 89208
rect 154311 87728 155111 87848
rect 0 87048 800 87168
rect 154311 86368 155111 86488
rect 0 85008 800 85128
rect 154311 84328 155111 84448
rect 0 82968 800 83088
rect 154311 82288 155111 82408
rect 0 81608 800 81728
rect 154311 80248 155111 80368
rect 0 79568 800 79688
rect 154311 78888 155111 79008
rect 0 77528 800 77648
rect 154311 76848 155111 76968
rect 0 75488 800 75608
rect 154311 74808 155111 74928
rect 0 73448 800 73568
rect 154311 72768 155111 72888
rect 0 72088 800 72208
rect 154311 71408 155111 71528
rect 0 70048 800 70168
rect 154311 69368 155111 69488
rect 0 68008 800 68128
rect 154311 67328 155111 67448
rect 0 65968 800 66088
rect 154311 65288 155111 65408
rect 0 64608 800 64728
rect 154311 63248 155111 63368
rect 0 62568 800 62688
rect 154311 61888 155111 62008
rect 0 60528 800 60648
rect 154311 59848 155111 59968
rect 0 58488 800 58608
rect 154311 57808 155111 57928
rect 0 57128 800 57248
rect 154311 55768 155111 55888
rect 0 55088 800 55208
rect 154311 54408 155111 54528
rect 0 53048 800 53168
rect 154311 52368 155111 52488
rect 0 51008 800 51128
rect 154311 50328 155111 50448
rect 0 48968 800 49088
rect 154311 48288 155111 48408
rect 0 47608 800 47728
rect 154311 46928 155111 47048
rect 0 45568 800 45688
rect 154311 44888 155111 45008
rect 0 43528 800 43648
rect 154311 42848 155111 42968
rect 0 41488 800 41608
rect 154311 40808 155111 40928
rect 0 40128 800 40248
rect 154311 39448 155111 39568
rect 0 38088 800 38208
rect 154311 37408 155111 37528
rect 0 36048 800 36168
rect 154311 35368 155111 35488
rect 0 34008 800 34128
rect 154311 33328 155111 33448
rect 0 32648 800 32768
rect 154311 31288 155111 31408
rect 0 30608 800 30728
rect 154311 29928 155111 30048
rect 0 28568 800 28688
rect 154311 27888 155111 28008
rect 0 26528 800 26648
rect 154311 25848 155111 25968
rect 0 24488 800 24608
rect 154311 23808 155111 23928
rect 0 23128 800 23248
rect 154311 22448 155111 22568
rect 0 21088 800 21208
rect 154311 20408 155111 20528
rect 0 19048 800 19168
rect 154311 18368 155111 18488
rect 0 17008 800 17128
rect 154311 16328 155111 16448
rect 0 15648 800 15768
rect 154311 14968 155111 15088
rect 0 13608 800 13728
rect 154311 12928 155111 13048
rect 0 11568 800 11688
rect 154311 10888 155111 11008
rect 0 9528 800 9648
rect 154311 8848 155111 8968
rect 0 8168 800 8288
rect 154311 6808 155111 6928
rect 0 6128 800 6248
rect 154311 5448 155111 5568
rect 0 4088 800 4208
rect 154311 3408 155111 3528
rect 0 2048 800 2168
rect 154311 1368 155111 1488
<< obsm3 >>
rect 880 156328 154311 156501
rect 800 155928 154311 156328
rect 800 155648 154231 155928
rect 800 154568 154311 155648
rect 880 154288 154311 154568
rect 800 153888 154311 154288
rect 800 153608 154231 153888
rect 800 153208 154311 153608
rect 880 152928 154311 153208
rect 800 152528 154311 152928
rect 800 152248 154231 152528
rect 800 151168 154311 152248
rect 880 150888 154311 151168
rect 800 150488 154311 150888
rect 800 150208 154231 150488
rect 800 149128 154311 150208
rect 880 148848 154311 149128
rect 800 148448 154311 148848
rect 800 148168 154231 148448
rect 800 147088 154311 148168
rect 880 146808 154311 147088
rect 800 146408 154311 146808
rect 800 146128 154231 146408
rect 800 145728 154311 146128
rect 880 145448 154311 145728
rect 800 145048 154311 145448
rect 800 144768 154231 145048
rect 800 143688 154311 144768
rect 880 143408 154311 143688
rect 800 143008 154311 143408
rect 800 142728 154231 143008
rect 800 141648 154311 142728
rect 880 141368 154311 141648
rect 800 140968 154311 141368
rect 800 140688 154231 140968
rect 800 139608 154311 140688
rect 880 139328 154311 139608
rect 800 138928 154311 139328
rect 800 138648 154231 138928
rect 800 138248 154311 138648
rect 880 137968 154311 138248
rect 800 136888 154311 137968
rect 800 136608 154231 136888
rect 800 136208 154311 136608
rect 880 135928 154311 136208
rect 800 135528 154311 135928
rect 800 135248 154231 135528
rect 800 134168 154311 135248
rect 880 133888 154311 134168
rect 800 133488 154311 133888
rect 800 133208 154231 133488
rect 800 132128 154311 133208
rect 880 131848 154311 132128
rect 800 131448 154311 131848
rect 800 131168 154231 131448
rect 800 130088 154311 131168
rect 880 129808 154311 130088
rect 800 129408 154311 129808
rect 800 129128 154231 129408
rect 800 128728 154311 129128
rect 880 128448 154311 128728
rect 800 128048 154311 128448
rect 800 127768 154231 128048
rect 800 126688 154311 127768
rect 880 126408 154311 126688
rect 800 126008 154311 126408
rect 800 125728 154231 126008
rect 800 124648 154311 125728
rect 880 124368 154311 124648
rect 800 123968 154311 124368
rect 800 123688 154231 123968
rect 800 122608 154311 123688
rect 880 122328 154311 122608
rect 800 121928 154311 122328
rect 800 121648 154231 121928
rect 800 121248 154311 121648
rect 880 120968 154311 121248
rect 800 120568 154311 120968
rect 800 120288 154231 120568
rect 800 119208 154311 120288
rect 880 118928 154311 119208
rect 800 118528 154311 118928
rect 800 118248 154231 118528
rect 800 117168 154311 118248
rect 880 116888 154311 117168
rect 800 116488 154311 116888
rect 800 116208 154231 116488
rect 800 115128 154311 116208
rect 880 114848 154311 115128
rect 800 114448 154311 114848
rect 800 114168 154231 114448
rect 800 113768 154311 114168
rect 880 113488 154311 113768
rect 800 112408 154311 113488
rect 800 112128 154231 112408
rect 800 111728 154311 112128
rect 880 111448 154311 111728
rect 800 111048 154311 111448
rect 800 110768 154231 111048
rect 800 109688 154311 110768
rect 880 109408 154311 109688
rect 800 109008 154311 109408
rect 800 108728 154231 109008
rect 800 107648 154311 108728
rect 880 107368 154311 107648
rect 800 106968 154311 107368
rect 800 106688 154231 106968
rect 800 105608 154311 106688
rect 880 105328 154311 105608
rect 800 104928 154311 105328
rect 800 104648 154231 104928
rect 800 104248 154311 104648
rect 880 103968 154311 104248
rect 800 103568 154311 103968
rect 800 103288 154231 103568
rect 800 102208 154311 103288
rect 880 101928 154311 102208
rect 800 101528 154311 101928
rect 800 101248 154231 101528
rect 800 100168 154311 101248
rect 880 99888 154311 100168
rect 800 99488 154311 99888
rect 800 99208 154231 99488
rect 800 98128 154311 99208
rect 880 97848 154311 98128
rect 800 97448 154311 97848
rect 800 97168 154231 97448
rect 800 96768 154311 97168
rect 880 96488 154311 96768
rect 800 96088 154311 96488
rect 800 95808 154231 96088
rect 800 94728 154311 95808
rect 880 94448 154311 94728
rect 800 94048 154311 94448
rect 800 93768 154231 94048
rect 800 92688 154311 93768
rect 880 92408 154311 92688
rect 800 92008 154311 92408
rect 800 91728 154231 92008
rect 800 90648 154311 91728
rect 880 90368 154311 90648
rect 800 89968 154311 90368
rect 800 89688 154231 89968
rect 800 89288 154311 89688
rect 880 89008 154311 89288
rect 800 87928 154311 89008
rect 800 87648 154231 87928
rect 800 87248 154311 87648
rect 880 86968 154311 87248
rect 800 86568 154311 86968
rect 800 86288 154231 86568
rect 800 85208 154311 86288
rect 880 84928 154311 85208
rect 800 84528 154311 84928
rect 800 84248 154231 84528
rect 800 83168 154311 84248
rect 880 82888 154311 83168
rect 800 82488 154311 82888
rect 800 82208 154231 82488
rect 800 81808 154311 82208
rect 880 81528 154311 81808
rect 800 80448 154311 81528
rect 800 80168 154231 80448
rect 800 79768 154311 80168
rect 880 79488 154311 79768
rect 800 79088 154311 79488
rect 800 78808 154231 79088
rect 800 77728 154311 78808
rect 880 77448 154311 77728
rect 800 77048 154311 77448
rect 800 76768 154231 77048
rect 800 75688 154311 76768
rect 880 75408 154311 75688
rect 800 75008 154311 75408
rect 800 74728 154231 75008
rect 800 73648 154311 74728
rect 880 73368 154311 73648
rect 800 72968 154311 73368
rect 800 72688 154231 72968
rect 800 72288 154311 72688
rect 880 72008 154311 72288
rect 800 71608 154311 72008
rect 800 71328 154231 71608
rect 800 70248 154311 71328
rect 880 69968 154311 70248
rect 800 69568 154311 69968
rect 800 69288 154231 69568
rect 800 68208 154311 69288
rect 880 67928 154311 68208
rect 800 67528 154311 67928
rect 800 67248 154231 67528
rect 800 66168 154311 67248
rect 880 65888 154311 66168
rect 800 65488 154311 65888
rect 800 65208 154231 65488
rect 800 64808 154311 65208
rect 880 64528 154311 64808
rect 800 63448 154311 64528
rect 800 63168 154231 63448
rect 800 62768 154311 63168
rect 880 62488 154311 62768
rect 800 62088 154311 62488
rect 800 61808 154231 62088
rect 800 60728 154311 61808
rect 880 60448 154311 60728
rect 800 60048 154311 60448
rect 800 59768 154231 60048
rect 800 58688 154311 59768
rect 880 58408 154311 58688
rect 800 58008 154311 58408
rect 800 57728 154231 58008
rect 800 57328 154311 57728
rect 880 57048 154311 57328
rect 800 55968 154311 57048
rect 800 55688 154231 55968
rect 800 55288 154311 55688
rect 880 55008 154311 55288
rect 800 54608 154311 55008
rect 800 54328 154231 54608
rect 800 53248 154311 54328
rect 880 52968 154311 53248
rect 800 52568 154311 52968
rect 800 52288 154231 52568
rect 800 51208 154311 52288
rect 880 50928 154311 51208
rect 800 50528 154311 50928
rect 800 50248 154231 50528
rect 800 49168 154311 50248
rect 880 48888 154311 49168
rect 800 48488 154311 48888
rect 800 48208 154231 48488
rect 800 47808 154311 48208
rect 880 47528 154311 47808
rect 800 47128 154311 47528
rect 800 46848 154231 47128
rect 800 45768 154311 46848
rect 880 45488 154311 45768
rect 800 45088 154311 45488
rect 800 44808 154231 45088
rect 800 43728 154311 44808
rect 880 43448 154311 43728
rect 800 43048 154311 43448
rect 800 42768 154231 43048
rect 800 41688 154311 42768
rect 880 41408 154311 41688
rect 800 41008 154311 41408
rect 800 40728 154231 41008
rect 800 40328 154311 40728
rect 880 40048 154311 40328
rect 800 39648 154311 40048
rect 800 39368 154231 39648
rect 800 38288 154311 39368
rect 880 38008 154311 38288
rect 800 37608 154311 38008
rect 800 37328 154231 37608
rect 800 36248 154311 37328
rect 880 35968 154311 36248
rect 800 35568 154311 35968
rect 800 35288 154231 35568
rect 800 34208 154311 35288
rect 880 33928 154311 34208
rect 800 33528 154311 33928
rect 800 33248 154231 33528
rect 800 32848 154311 33248
rect 880 32568 154311 32848
rect 800 31488 154311 32568
rect 800 31208 154231 31488
rect 800 30808 154311 31208
rect 880 30528 154311 30808
rect 800 30128 154311 30528
rect 800 29848 154231 30128
rect 800 28768 154311 29848
rect 880 28488 154311 28768
rect 800 28088 154311 28488
rect 800 27808 154231 28088
rect 800 26728 154311 27808
rect 880 26448 154311 26728
rect 800 26048 154311 26448
rect 800 25768 154231 26048
rect 800 24688 154311 25768
rect 880 24408 154311 24688
rect 800 24008 154311 24408
rect 800 23728 154231 24008
rect 800 23328 154311 23728
rect 880 23048 154311 23328
rect 800 22648 154311 23048
rect 800 22368 154231 22648
rect 800 21288 154311 22368
rect 880 21008 154311 21288
rect 800 20608 154311 21008
rect 800 20328 154231 20608
rect 800 19248 154311 20328
rect 880 18968 154311 19248
rect 800 18568 154311 18968
rect 800 18288 154231 18568
rect 800 17208 154311 18288
rect 880 16928 154311 17208
rect 800 16528 154311 16928
rect 800 16248 154231 16528
rect 800 15848 154311 16248
rect 880 15568 154311 15848
rect 800 15168 154311 15568
rect 800 14888 154231 15168
rect 800 13808 154311 14888
rect 880 13528 154311 13808
rect 800 13128 154311 13528
rect 800 12848 154231 13128
rect 800 11768 154311 12848
rect 880 11488 154311 11768
rect 800 11088 154311 11488
rect 800 10808 154231 11088
rect 800 9728 154311 10808
rect 880 9448 154311 9728
rect 800 9048 154311 9448
rect 800 8768 154231 9048
rect 800 8368 154311 8768
rect 880 8088 154311 8368
rect 800 7008 154311 8088
rect 800 6728 154231 7008
rect 800 6328 154311 6728
rect 880 6048 154311 6328
rect 800 5648 154311 6048
rect 800 5368 154231 5648
rect 800 4288 154311 5368
rect 880 4008 154311 4288
rect 800 3608 154311 4008
rect 800 3328 154231 3608
rect 800 2248 154311 3328
rect 880 1968 154311 2248
rect 800 1568 154311 1968
rect 800 1395 154231 1568
<< metal4 >>
rect 4208 2128 4528 155088
rect 19568 2128 19888 155088
rect 34928 2128 35248 155088
rect 50288 2128 50608 155088
rect 65648 2128 65968 155088
rect 81008 2128 81328 155088
rect 96368 2128 96688 155088
rect 111728 2128 112048 155088
rect 127088 2128 127408 155088
rect 142448 2128 142768 155088
<< obsm4 >>
rect 20115 155168 145669 155413
rect 20115 2048 34848 155168
rect 35328 2048 50208 155168
rect 50688 2048 65568 155168
rect 66048 2048 80928 155168
rect 81408 2048 96288 155168
rect 96768 2048 111648 155168
rect 112128 2048 127008 155168
rect 127488 2048 142368 155168
rect 142848 2048 145669 155168
rect 20115 1939 145669 2048
<< metal5 >>
rect 1104 143160 153916 143480
rect 1104 127842 153916 128162
rect 1104 112524 153916 112844
rect 1104 97206 153916 97526
rect 1104 81888 153916 82208
rect 1104 66570 153916 66890
rect 1104 51252 153916 51572
rect 1104 35934 153916 36254
rect 1104 20616 153916 20936
rect 1104 5298 153916 5618
<< obsm5 >>
rect 47956 82528 115068 88220
rect 47956 75660 115068 81568
<< labels >>
rlabel metal2 s 135258 156455 135314 157255 6 clk
port 1 nsew signal input
rlabel metal2 s 47398 156455 47454 157255 6 eoi[0]
port 2 nsew signal output
rlabel metal3 s 154311 48288 155111 48408 6 eoi[10]
port 3 nsew signal output
rlabel metal2 s 17958 156455 18014 157255 6 eoi[11]
port 4 nsew signal output
rlabel metal2 s 44638 156455 44694 157255 6 eoi[12]
port 5 nsew signal output
rlabel metal3 s 154311 89768 155111 89888 6 eoi[13]
port 6 nsew signal output
rlabel metal3 s 0 28568 800 28688 6 eoi[14]
port 7 nsew signal output
rlabel metal2 s 11518 0 11574 800 6 eoi[15]
port 8 nsew signal output
rlabel metal3 s 154311 14968 155111 15088 6 eoi[16]
port 9 nsew signal output
rlabel metal2 s 130198 0 130254 800 6 eoi[17]
port 10 nsew signal output
rlabel metal3 s 0 30608 800 30728 6 eoi[18]
port 11 nsew signal output
rlabel metal3 s 154311 106768 155111 106888 6 eoi[19]
port 12 nsew signal output
rlabel metal3 s 0 15648 800 15768 6 eoi[1]
port 13 nsew signal output
rlabel metal2 s 142618 0 142674 800 6 eoi[20]
port 14 nsew signal output
rlabel metal2 s 107198 156455 107254 157255 6 eoi[21]
port 15 nsew signal output
rlabel metal3 s 0 48968 800 49088 6 eoi[22]
port 16 nsew signal output
rlabel metal2 s 148138 0 148194 800 6 eoi[23]
port 17 nsew signal output
rlabel metal3 s 0 81608 800 81728 6 eoi[24]
port 18 nsew signal output
rlabel metal2 s 14278 0 14334 800 6 eoi[25]
port 19 nsew signal output
rlabel metal3 s 0 96568 800 96688 6 eoi[26]
port 20 nsew signal output
rlabel metal2 s 67638 156455 67694 157255 6 eoi[27]
port 21 nsew signal output
rlabel metal3 s 0 143488 800 143608 6 eoi[28]
port 22 nsew signal output
rlabel metal2 s 21638 156455 21694 157255 6 eoi[29]
port 23 nsew signal output
rlabel metal2 s 153198 0 153254 800 6 eoi[2]
port 24 nsew signal output
rlabel metal2 s 35898 0 35954 800 6 eoi[30]
port 25 nsew signal output
rlabel metal2 s 69018 0 69074 800 6 eoi[31]
port 26 nsew signal output
rlabel metal2 s 115018 0 115074 800 6 eoi[3]
port 27 nsew signal output
rlabel metal3 s 0 104048 800 104168 6 eoi[4]
port 28 nsew signal output
rlabel metal2 s 89258 156455 89314 157255 6 eoi[5]
port 29 nsew signal output
rlabel metal3 s 154311 93848 155111 93968 6 eoi[6]
port 30 nsew signal output
rlabel metal2 s 38658 0 38714 800 6 eoi[7]
port 31 nsew signal output
rlabel metal3 s 0 146888 800 147008 6 eoi[8]
port 32 nsew signal output
rlabel metal2 s 43258 156455 43314 157255 6 eoi[9]
port 33 nsew signal output
rlabel metal3 s 154311 84328 155111 84448 6 irq[0]
port 34 nsew signal input
rlabel metal2 s 140318 156455 140374 157255 6 irq[10]
port 35 nsew signal input
rlabel metal3 s 154311 55768 155111 55888 6 irq[11]
port 36 nsew signal input
rlabel metal2 s 11518 156455 11574 157255 6 irq[12]
port 37 nsew signal input
rlabel metal2 s 77758 156455 77814 157255 6 irq[13]
port 38 nsew signal input
rlabel metal3 s 0 133968 800 134088 6 irq[14]
port 39 nsew signal input
rlabel metal3 s 154311 131248 155111 131368 6 irq[15]
port 40 nsew signal input
rlabel metal2 s 86958 0 87014 800 6 irq[16]
port 41 nsew signal input
rlabel metal2 s 136638 0 136694 800 6 irq[17]
port 42 nsew signal input
rlabel metal3 s 0 23128 800 23248 6 irq[18]
port 43 nsew signal input
rlabel metal3 s 0 34008 800 34128 6 irq[19]
port 44 nsew signal input
rlabel metal2 s 69938 156455 69994 157255 6 irq[1]
port 45 nsew signal input
rlabel metal2 s 123758 156455 123814 157255 6 irq[20]
port 46 nsew signal input
rlabel metal2 s 97078 156455 97134 157255 6 irq[21]
port 47 nsew signal input
rlabel metal2 s 23018 0 23074 800 6 irq[22]
port 48 nsew signal input
rlabel metal2 s 65338 0 65394 800 6 irq[23]
port 49 nsew signal input
rlabel metal2 s 30838 156455 30894 157255 6 irq[24]
port 50 nsew signal input
rlabel metal2 s 107198 0 107254 800 6 irq[25]
port 51 nsew signal input
rlabel metal3 s 0 111528 800 111648 6 irq[26]
port 52 nsew signal input
rlabel metal3 s 154311 148248 155111 148368 6 irq[27]
port 53 nsew signal input
rlabel metal3 s 154311 140768 155111 140888 6 irq[28]
port 54 nsew signal input
rlabel metal3 s 154311 50328 155111 50448 6 irq[29]
port 55 nsew signal input
rlabel metal3 s 154311 40808 155111 40928 6 irq[2]
port 56 nsew signal input
rlabel metal2 s 52458 156455 52514 157255 6 irq[30]
port 57 nsew signal input
rlabel metal3 s 154311 120368 155111 120488 6 irq[31]
port 58 nsew signal input
rlabel metal2 s 39578 156455 39634 157255 6 irq[3]
port 59 nsew signal input
rlabel metal3 s 154311 16328 155111 16448 6 irq[4]
port 60 nsew signal input
rlabel metal2 s 74078 0 74134 800 6 irq[5]
port 61 nsew signal input
rlabel metal3 s 154311 8848 155111 8968 6 irq[6]
port 62 nsew signal input
rlabel metal2 s 147678 156455 147734 157255 6 irq[7]
port 63 nsew signal input
rlabel metal2 s 47398 0 47454 800 6 irq[8]
port 64 nsew signal input
rlabel metal2 s 131578 0 131634 800 6 irq[9]
port 65 nsew signal input
rlabel metal3 s 0 148928 800 149048 6 mem_addr[0]
port 66 nsew signal output
rlabel metal2 s 28078 156455 28134 157255 6 mem_addr[10]
port 67 nsew signal output
rlabel metal2 s 143998 0 144054 800 6 mem_addr[11]
port 68 nsew signal output
rlabel metal3 s 154311 101328 155111 101448 6 mem_addr[12]
port 69 nsew signal output
rlabel metal3 s 154311 67328 155111 67448 6 mem_addr[13]
port 70 nsew signal output
rlabel metal2 s 7838 0 7894 800 6 mem_addr[14]
port 71 nsew signal output
rlabel metal2 s 70398 0 70454 800 6 mem_addr[15]
port 72 nsew signal output
rlabel metal2 s 80518 156455 80574 157255 6 mem_addr[16]
port 73 nsew signal output
rlabel metal3 s 0 126488 800 126608 6 mem_addr[17]
port 74 nsew signal output
rlabel metal2 s 137558 156455 137614 157255 6 mem_addr[18]
port 75 nsew signal output
rlabel metal2 s 51078 0 51134 800 6 mem_addr[19]
port 76 nsew signal output
rlabel metal3 s 0 141448 800 141568 6 mem_addr[1]
port 77 nsew signal output
rlabel metal2 s 113638 156455 113694 157255 6 mem_addr[20]
port 78 nsew signal output
rlabel metal3 s 154311 33328 155111 33448 6 mem_addr[21]
port 79 nsew signal output
rlabel metal2 s 75458 156455 75514 157255 6 mem_addr[22]
port 80 nsew signal output
rlabel metal3 s 0 19048 800 19168 6 mem_addr[23]
port 81 nsew signal output
rlabel metal2 s 4158 0 4214 800 6 mem_addr[24]
port 82 nsew signal output
rlabel metal3 s 154311 82288 155111 82408 6 mem_addr[25]
port 83 nsew signal output
rlabel metal2 s 146758 156455 146814 157255 6 mem_addr[26]
port 84 nsew signal output
rlabel metal2 s 49698 156455 49754 157255 6 mem_addr[27]
port 85 nsew signal output
rlabel metal3 s 154311 12928 155111 13048 6 mem_addr[28]
port 86 nsew signal output
rlabel metal3 s 154311 69368 155111 69488 6 mem_addr[29]
port 87 nsew signal output
rlabel metal2 s 63958 156455 64014 157255 6 mem_addr[2]
port 88 nsew signal output
rlabel metal3 s 0 64608 800 64728 6 mem_addr[30]
port 89 nsew signal output
rlabel metal2 s 115938 0 115994 800 6 mem_addr[31]
port 90 nsew signal output
rlabel metal2 s 92938 156455 92994 157255 6 mem_addr[3]
port 91 nsew signal output
rlabel metal2 s 49698 0 49754 800 6 mem_addr[4]
port 92 nsew signal output
rlabel metal2 s 37278 0 37334 800 6 mem_addr[5]
port 93 nsew signal output
rlabel metal2 s 151818 156455 151874 157255 6 mem_addr[6]
port 94 nsew signal output
rlabel metal2 s 108118 156455 108174 157255 6 mem_addr[7]
port 95 nsew signal output
rlabel metal2 s 98458 0 98514 800 6 mem_addr[8]
port 96 nsew signal output
rlabel metal3 s 0 109488 800 109608 6 mem_addr[9]
port 97 nsew signal output
rlabel metal3 s 0 57128 800 57248 6 mem_instr
port 98 nsew signal output
rlabel metal3 s 154311 127848 155111 127968 6 mem_la_addr[0]
port 99 nsew signal output
rlabel metal2 s 61198 156455 61254 157255 6 mem_la_addr[10]
port 100 nsew signal output
rlabel metal3 s 154311 78888 155111 79008 6 mem_la_addr[11]
port 101 nsew signal output
rlabel metal2 s 85578 0 85634 800 6 mem_la_addr[12]
port 102 nsew signal output
rlabel metal2 s 112258 156455 112314 157255 6 mem_la_addr[13]
port 103 nsew signal output
rlabel metal2 s 151818 0 151874 800 6 mem_la_addr[14]
port 104 nsew signal output
rlabel metal2 s 76838 0 76894 800 6 mem_la_addr[15]
port 105 nsew signal output
rlabel metal3 s 0 136008 800 136128 6 mem_la_addr[16]
port 106 nsew signal output
rlabel metal3 s 0 89088 800 89208 6 mem_la_addr[17]
port 107 nsew signal output
rlabel metal2 s 120078 0 120134 800 6 mem_la_addr[18]
port 108 nsew signal output
rlabel metal2 s 74078 156455 74134 157255 6 mem_la_addr[19]
port 109 nsew signal output
rlabel metal3 s 0 150968 800 151088 6 mem_la_addr[1]
port 110 nsew signal output
rlabel metal2 s 141698 0 141754 800 6 mem_la_addr[20]
port 111 nsew signal output
rlabel metal3 s 0 128528 800 128648 6 mem_la_addr[21]
port 112 nsew signal output
rlabel metal2 s 16578 156455 16634 157255 6 mem_la_addr[22]
port 113 nsew signal output
rlabel metal3 s 154311 39448 155111 39568 6 mem_la_addr[23]
port 114 nsew signal output
rlabel metal2 s 150438 156455 150494 157255 6 mem_la_addr[24]
port 115 nsew signal output
rlabel metal2 s 117318 0 117374 800 6 mem_la_addr[25]
port 116 nsew signal output
rlabel metal2 s 19338 0 19394 800 6 mem_la_addr[26]
port 117 nsew signal output
rlabel metal3 s 0 55088 800 55208 6 mem_la_addr[27]
port 118 nsew signal output
rlabel metal2 s 59818 156455 59874 157255 6 mem_la_addr[28]
port 119 nsew signal output
rlabel metal3 s 154311 144848 155111 144968 6 mem_la_addr[29]
port 120 nsew signal output
rlabel metal2 s 120998 156455 121054 157255 6 mem_la_addr[2]
port 121 nsew signal output
rlabel metal2 s 33138 156455 33194 157255 6 mem_la_addr[30]
port 122 nsew signal output
rlabel metal2 s 104438 0 104494 800 6 mem_la_addr[31]
port 123 nsew signal output
rlabel metal2 s 103518 0 103574 800 6 mem_la_addr[3]
port 124 nsew signal output
rlabel metal3 s 0 139408 800 139528 6 mem_la_addr[4]
port 125 nsew signal output
rlabel metal3 s 154311 76848 155111 76968 6 mem_la_addr[5]
port 126 nsew signal output
rlabel metal2 s 145378 0 145434 800 6 mem_la_addr[6]
port 127 nsew signal output
rlabel metal3 s 154311 22448 155111 22568 6 mem_la_addr[7]
port 128 nsew signal output
rlabel metal3 s 154311 25848 155111 25968 6 mem_la_addr[8]
port 129 nsew signal output
rlabel metal2 s 76378 156455 76434 157255 6 mem_la_addr[9]
port 130 nsew signal output
rlabel metal2 s 126058 156455 126114 157255 6 mem_la_read
port 131 nsew signal output
rlabel metal2 s 95698 0 95754 800 6 mem_la_wdata[0]
port 132 nsew signal output
rlabel metal2 s 112258 0 112314 800 6 mem_la_wdata[10]
port 133 nsew signal output
rlabel metal2 s 100758 156455 100814 157255 6 mem_la_wdata[11]
port 134 nsew signal output
rlabel metal2 s 82818 0 82874 800 6 mem_la_wdata[12]
port 135 nsew signal output
rlabel metal2 s 77758 0 77814 800 6 mem_la_wdata[13]
port 136 nsew signal output
rlabel metal2 s 2778 156455 2834 157255 6 mem_la_wdata[14]
port 137 nsew signal output
rlabel metal3 s 0 94528 800 94648 6 mem_la_wdata[15]
port 138 nsew signal output
rlabel metal3 s 0 153008 800 153128 6 mem_la_wdata[16]
port 139 nsew signal output
rlabel metal3 s 154311 86368 155111 86488 6 mem_la_wdata[17]
port 140 nsew signal output
rlabel metal3 s 0 129888 800 130008 6 mem_la_wdata[18]
port 141 nsew signal output
rlabel metal3 s 154311 95888 155111 96008 6 mem_la_wdata[19]
port 142 nsew signal output
rlabel metal2 s 82818 156455 82874 157255 6 mem_la_wdata[1]
port 143 nsew signal output
rlabel metal2 s 52458 0 52514 800 6 mem_la_wdata[20]
port 144 nsew signal output
rlabel metal3 s 154311 91808 155111 91928 6 mem_la_wdata[21]
port 145 nsew signal output
rlabel metal3 s 154311 110848 155111 110968 6 mem_la_wdata[22]
port 146 nsew signal output
rlabel metal2 s 132498 156455 132554 157255 6 mem_la_wdata[23]
port 147 nsew signal output
rlabel metal3 s 0 77528 800 77648 6 mem_la_wdata[24]
port 148 nsew signal output
rlabel metal2 s 146758 0 146814 800 6 mem_la_wdata[25]
port 149 nsew signal output
rlabel metal3 s 154311 1368 155111 1488 6 mem_la_wdata[26]
port 150 nsew signal output
rlabel metal2 s 32218 0 32274 800 6 mem_la_wdata[27]
port 151 nsew signal output
rlabel metal2 s 48318 156455 48374 157255 6 mem_la_wdata[28]
port 152 nsew signal output
rlabel metal3 s 154311 52368 155111 52488 6 mem_la_wdata[29]
port 153 nsew signal output
rlabel metal2 s 56138 0 56194 800 6 mem_la_wdata[2]
port 154 nsew signal output
rlabel metal3 s 154311 10888 155111 11008 6 mem_la_wdata[30]
port 155 nsew signal output
rlabel metal2 s 58898 156455 58954 157255 6 mem_la_wdata[31]
port 156 nsew signal output
rlabel metal3 s 0 119008 800 119128 6 mem_la_wdata[3]
port 157 nsew signal output
rlabel metal2 s 85578 156455 85634 157255 6 mem_la_wdata[4]
port 158 nsew signal output
rlabel metal3 s 154311 97248 155111 97368 6 mem_la_wdata[5]
port 159 nsew signal output
rlabel metal3 s 0 6128 800 6248 6 mem_la_wdata[6]
port 160 nsew signal output
rlabel metal2 s 136178 156455 136234 157255 6 mem_la_wdata[7]
port 161 nsew signal output
rlabel metal2 s 71318 156455 71374 157255 6 mem_la_wdata[8]
port 162 nsew signal output
rlabel metal2 s 133878 0 133934 800 6 mem_la_wdata[9]
port 163 nsew signal output
rlabel metal2 s 1398 0 1454 800 6 mem_la_write
port 164 nsew signal output
rlabel metal3 s 0 58488 800 58608 6 mem_la_wstrb[0]
port 165 nsew signal output
rlabel metal2 s 109498 156455 109554 157255 6 mem_la_wstrb[1]
port 166 nsew signal output
rlabel metal3 s 0 38088 800 38208 6 mem_la_wstrb[2]
port 167 nsew signal output
rlabel metal2 s 55218 0 55274 800 6 mem_la_wstrb[3]
port 168 nsew signal output
rlabel metal2 s 6458 0 6514 800 6 mem_rdata[0]
port 169 nsew signal input
rlabel metal3 s 0 97928 800 98048 6 mem_rdata[10]
port 170 nsew signal input
rlabel metal2 s 94318 0 94374 800 6 mem_rdata[11]
port 171 nsew signal input
rlabel metal3 s 154311 153688 155111 153808 6 mem_rdata[12]
port 172 nsew signal input
rlabel metal2 s 67638 0 67694 800 6 mem_rdata[13]
port 173 nsew signal input
rlabel metal3 s 0 26528 800 26648 6 mem_rdata[14]
port 174 nsew signal input
rlabel metal3 s 154311 152328 155111 152448 6 mem_rdata[15]
port 175 nsew signal input
rlabel metal2 s 46018 156455 46074 157255 6 mem_rdata[16]
port 176 nsew signal input
rlabel metal2 s 15198 156455 15254 157255 6 mem_rdata[17]
port 177 nsew signal input
rlabel metal2 s 28078 0 28134 800 6 mem_rdata[18]
port 178 nsew signal input
rlabel metal3 s 154311 133288 155111 133408 6 mem_rdata[19]
port 179 nsew signal input
rlabel metal2 s 132498 0 132554 800 6 mem_rdata[1]
port 180 nsew signal input
rlabel metal3 s 154311 5448 155111 5568 6 mem_rdata[20]
port 181 nsew signal input
rlabel metal3 s 0 70048 800 70168 6 mem_rdata[21]
port 182 nsew signal input
rlabel metal2 s 105818 156455 105874 157255 6 mem_rdata[22]
port 183 nsew signal input
rlabel metal3 s 0 73448 800 73568 6 mem_rdata[23]
port 184 nsew signal input
rlabel metal3 s 0 32648 800 32768 6 mem_rdata[24]
port 185 nsew signal input
rlabel metal2 s 102138 156455 102194 157255 6 mem_rdata[25]
port 186 nsew signal input
rlabel metal2 s 24398 156455 24454 157255 6 mem_rdata[26]
port 187 nsew signal input
rlabel metal2 s 102138 0 102194 800 6 mem_rdata[27]
port 188 nsew signal input
rlabel metal3 s 0 53048 800 53168 6 mem_rdata[28]
port 189 nsew signal input
rlabel metal3 s 154311 54408 155111 54528 6 mem_rdata[29]
port 190 nsew signal input
rlabel metal2 s 92018 0 92074 800 6 mem_rdata[2]
port 191 nsew signal input
rlabel metal2 s 143998 156455 144054 157255 6 mem_rdata[30]
port 192 nsew signal input
rlabel metal2 s 108578 0 108634 800 6 mem_rdata[31]
port 193 nsew signal input
rlabel metal3 s 0 4088 800 4208 6 mem_rdata[3]
port 194 nsew signal input
rlabel metal2 s 119618 156455 119674 157255 6 mem_rdata[4]
port 195 nsew signal input
rlabel metal3 s 154311 150288 155111 150408 6 mem_rdata[5]
port 196 nsew signal input
rlabel metal2 s 478 0 534 800 6 mem_rdata[6]
port 197 nsew signal input
rlabel metal2 s 23018 156455 23074 157255 6 mem_rdata[7]
port 198 nsew signal input
rlabel metal2 s 114558 156455 114614 157255 6 mem_rdata[8]
port 199 nsew signal input
rlabel metal3 s 0 102008 800 102128 6 mem_rdata[9]
port 200 nsew signal input
rlabel metal2 s 141238 156455 141294 157255 6 mem_ready
port 201 nsew signal input
rlabel metal3 s 0 45568 800 45688 6 mem_valid
port 202 nsew signal output
rlabel metal3 s 0 47608 800 47728 6 mem_wdata[0]
port 203 nsew signal output
rlabel metal2 s 1398 156455 1454 157255 6 mem_wdata[10]
port 204 nsew signal output
rlabel metal2 s 133878 156455 133934 157255 6 mem_wdata[11]
port 205 nsew signal output
rlabel metal3 s 0 116968 800 117088 6 mem_wdata[12]
port 206 nsew signal output
rlabel metal2 s 53838 0 53894 800 6 mem_wdata[13]
port 207 nsew signal output
rlabel metal2 s 97998 156455 98054 157255 6 mem_wdata[14]
port 208 nsew signal output
rlabel metal3 s 154311 37408 155111 37528 6 mem_wdata[15]
port 209 nsew signal output
rlabel metal3 s 0 68008 800 68128 6 mem_wdata[16]
port 210 nsew signal output
rlabel metal2 s 36818 156455 36874 157255 6 mem_wdata[17]
port 211 nsew signal output
rlabel metal2 s 81898 0 81954 800 6 mem_wdata[18]
port 212 nsew signal output
rlabel metal2 s 127438 0 127494 800 6 mem_wdata[19]
port 213 nsew signal output
rlabel metal2 s 34518 156455 34574 157255 6 mem_wdata[1]
port 214 nsew signal output
rlabel metal3 s 154311 135328 155111 135448 6 mem_wdata[20]
port 215 nsew signal output
rlabel metal2 s 89258 0 89314 800 6 mem_wdata[21]
port 216 nsew signal output
rlabel metal2 s 72698 156455 72754 157255 6 mem_wdata[22]
port 217 nsew signal output
rlabel metal2 s 57518 156455 57574 157255 6 mem_wdata[23]
port 218 nsew signal output
rlabel metal2 s 94318 156455 94374 157255 6 mem_wdata[24]
port 219 nsew signal output
rlabel metal2 s 56138 156455 56194 157255 6 mem_wdata[25]
port 220 nsew signal output
rlabel metal2 s 31758 156455 31814 157255 6 mem_wdata[26]
port 221 nsew signal output
rlabel metal2 s 149058 0 149114 800 6 mem_wdata[27]
port 222 nsew signal output
rlabel metal3 s 154311 103368 155111 103488 6 mem_wdata[28]
port 223 nsew signal output
rlabel metal3 s 0 113568 800 113688 6 mem_wdata[29]
port 224 nsew signal output
rlabel metal3 s 154311 108808 155111 108928 6 mem_wdata[2]
port 225 nsew signal output
rlabel metal3 s 0 145528 800 145648 6 mem_wdata[30]
port 226 nsew signal output
rlabel metal2 s 115938 156455 115994 157255 6 mem_wdata[31]
port 227 nsew signal output
rlabel metal3 s 0 131928 800 132048 6 mem_wdata[3]
port 228 nsew signal output
rlabel metal3 s 154311 57808 155111 57928 6 mem_wdata[4]
port 229 nsew signal output
rlabel metal3 s 0 124448 800 124568 6 mem_wdata[5]
port 230 nsew signal output
rlabel metal2 s 135258 0 135314 800 6 mem_wdata[6]
port 231 nsew signal output
rlabel metal3 s 154311 112208 155111 112328 6 mem_wdata[7]
port 232 nsew signal output
rlabel metal2 s 34518 0 34574 800 6 mem_wdata[8]
port 233 nsew signal output
rlabel metal2 s 72698 0 72754 800 6 mem_wdata[9]
port 234 nsew signal output
rlabel metal2 s 150438 0 150494 800 6 mem_wstrb[0]
port 235 nsew signal output
rlabel metal2 s 127438 156455 127494 157255 6 mem_wstrb[1]
port 236 nsew signal output
rlabel metal2 s 12898 156455 12954 157255 6 mem_wstrb[2]
port 237 nsew signal output
rlabel metal2 s 40958 0 41014 800 6 mem_wstrb[3]
port 238 nsew signal output
rlabel metal2 s 126518 0 126574 800 6 pcpi_insn[0]
port 239 nsew signal output
rlabel metal2 s 42338 156455 42394 157255 6 pcpi_insn[10]
port 240 nsew signal output
rlabel metal2 s 29458 156455 29514 157255 6 pcpi_insn[11]
port 241 nsew signal output
rlabel metal3 s 0 51008 800 51128 6 pcpi_insn[12]
port 242 nsew signal output
rlabel metal2 s 124678 156455 124734 157255 6 pcpi_insn[13]
port 243 nsew signal output
rlabel metal3 s 154311 121728 155111 121848 6 pcpi_insn[14]
port 244 nsew signal output
rlabel metal3 s 154311 3408 155111 3528 6 pcpi_insn[15]
port 245 nsew signal output
rlabel metal2 s 46018 0 46074 800 6 pcpi_insn[16]
port 246 nsew signal output
rlabel metal3 s 154311 61888 155111 62008 6 pcpi_insn[17]
port 247 nsew signal output
rlabel metal2 s 90638 156455 90694 157255 6 pcpi_insn[18]
port 248 nsew signal output
rlabel metal3 s 0 107448 800 107568 6 pcpi_insn[19]
port 249 nsew signal output
rlabel metal2 s 60278 0 60334 800 6 pcpi_insn[1]
port 250 nsew signal output
rlabel metal3 s 154311 104728 155111 104848 6 pcpi_insn[20]
port 251 nsew signal output
rlabel metal2 s 71318 0 71374 800 6 pcpi_insn[21]
port 252 nsew signal output
rlabel metal3 s 0 121048 800 121168 6 pcpi_insn[22]
port 253 nsew signal output
rlabel metal2 s 7838 156455 7894 157255 6 pcpi_insn[23]
port 254 nsew signal output
rlabel metal2 s 38198 156455 38254 157255 6 pcpi_insn[24]
port 255 nsew signal output
rlabel metal3 s 0 13608 800 13728 6 pcpi_insn[25]
port 256 nsew signal output
rlabel metal3 s 0 85008 800 85128 6 pcpi_insn[26]
port 257 nsew signal output
rlabel metal3 s 154311 42848 155111 42968 6 pcpi_insn[27]
port 258 nsew signal output
rlabel metal3 s 0 8168 800 8288 6 pcpi_insn[28]
port 259 nsew signal output
rlabel metal3 s 154311 46928 155111 47048 6 pcpi_insn[29]
port 260 nsew signal output
rlabel metal2 s 69018 156455 69074 157255 6 pcpi_insn[2]
port 261 nsew signal output
rlabel metal3 s 0 82968 800 83088 6 pcpi_insn[30]
port 262 nsew signal output
rlabel metal2 s 5538 0 5594 800 6 pcpi_insn[31]
port 263 nsew signal output
rlabel metal2 s 87878 156455 87934 157255 6 pcpi_insn[3]
port 264 nsew signal output
rlabel metal2 s 12898 0 12954 800 6 pcpi_insn[4]
port 265 nsew signal output
rlabel metal3 s 154311 63248 155111 63368 6 pcpi_insn[5]
port 266 nsew signal output
rlabel metal2 s 24398 0 24454 800 6 pcpi_insn[6]
port 267 nsew signal output
rlabel metal3 s 154311 123768 155111 123888 6 pcpi_insn[7]
port 268 nsew signal output
rlabel metal3 s 0 72088 800 72208 6 pcpi_insn[8]
port 269 nsew signal output
rlabel metal2 s 84198 156455 84254 157255 6 pcpi_insn[9]
port 270 nsew signal output
rlabel metal3 s 0 114928 800 115048 6 pcpi_rd[0]
port 271 nsew signal input
rlabel metal3 s 154311 44888 155111 45008 6 pcpi_rd[10]
port 272 nsew signal input
rlabel metal2 s 118698 0 118754 800 6 pcpi_rd[11]
port 273 nsew signal input
rlabel metal3 s 154311 23808 155111 23928 6 pcpi_rd[12]
port 274 nsew signal input
rlabel metal2 s 62578 156455 62634 157255 6 pcpi_rd[13]
port 275 nsew signal input
rlabel metal3 s 0 41488 800 41608 6 pcpi_rd[14]
port 276 nsew signal input
rlabel metal3 s 0 17008 800 17128 6 pcpi_rd[15]
port 277 nsew signal input
rlabel metal2 s 6458 156455 6514 157255 6 pcpi_rd[16]
port 278 nsew signal input
rlabel metal3 s 154311 20408 155111 20528 6 pcpi_rd[17]
port 279 nsew signal input
rlabel metal2 s 97078 0 97134 800 6 pcpi_rd[18]
port 280 nsew signal input
rlabel metal3 s 154311 129208 155111 129328 6 pcpi_rd[19]
port 281 nsew signal input
rlabel metal3 s 0 75488 800 75608 6 pcpi_rd[1]
port 282 nsew signal input
rlabel metal2 s 20718 0 20774 800 6 pcpi_rd[20]
port 283 nsew signal input
rlabel metal2 s 33138 0 33194 800 6 pcpi_rd[21]
port 284 nsew signal input
rlabel metal2 s 66258 0 66314 800 6 pcpi_rd[22]
port 285 nsew signal input
rlabel metal2 s 138938 0 138994 800 6 pcpi_rd[23]
port 286 nsew signal input
rlabel metal3 s 0 99968 800 100088 6 pcpi_rd[24]
port 287 nsew signal input
rlabel metal3 s 0 40128 800 40248 6 pcpi_rd[25]
port 288 nsew signal input
rlabel metal3 s 154311 31288 155111 31408 6 pcpi_rd[26]
port 289 nsew signal input
rlabel metal2 s 19338 156455 19394 157255 6 pcpi_rd[27]
port 290 nsew signal input
rlabel metal3 s 154311 125808 155111 125928 6 pcpi_rd[28]
port 291 nsew signal input
rlabel metal3 s 0 36048 800 36168 6 pcpi_rd[29]
port 292 nsew signal input
rlabel metal2 s 9218 156455 9274 157255 6 pcpi_rd[2]
port 293 nsew signal input
rlabel metal2 s 51078 156455 51134 157255 6 pcpi_rd[30]
port 294 nsew signal input
rlabel metal2 s 90638 0 90694 800 6 pcpi_rd[31]
port 295 nsew signal input
rlabel metal2 s 61198 0 61254 800 6 pcpi_rd[3]
port 296 nsew signal input
rlabel metal2 s 20718 156455 20774 157255 6 pcpi_rd[4]
port 297 nsew signal input
rlabel metal2 s 5078 156455 5134 157255 6 pcpi_rd[5]
port 298 nsew signal input
rlabel metal3 s 154311 114248 155111 114368 6 pcpi_rd[6]
port 299 nsew signal input
rlabel metal2 s 80518 0 80574 800 6 pcpi_rd[7]
port 300 nsew signal input
rlabel metal3 s 154311 35368 155111 35488 6 pcpi_rd[8]
port 301 nsew signal input
rlabel metal3 s 0 43528 800 43648 6 pcpi_rd[9]
port 302 nsew signal input
rlabel metal2 s 81438 156455 81494 157255 6 pcpi_ready
port 303 nsew signal input
rlabel metal3 s 154311 87728 155111 87848 6 pcpi_rs1[0]
port 304 nsew signal output
rlabel metal2 s 103058 156455 103114 157255 6 pcpi_rs1[10]
port 305 nsew signal output
rlabel metal2 s 16578 0 16634 800 6 pcpi_rs1[11]
port 306 nsew signal output
rlabel metal2 s 27158 0 27214 800 6 pcpi_rs1[12]
port 307 nsew signal output
rlabel metal3 s 154311 118328 155111 118448 6 pcpi_rs1[13]
port 308 nsew signal output
rlabel metal3 s 0 92488 800 92608 6 pcpi_rs1[14]
port 309 nsew signal output
rlabel metal2 s 120998 0 121054 800 6 pcpi_rs1[15]
port 310 nsew signal output
rlabel metal2 s 100758 0 100814 800 6 pcpi_rs1[16]
port 311 nsew signal output
rlabel metal3 s 154311 18368 155111 18488 6 pcpi_rs1[17]
port 312 nsew signal output
rlabel metal3 s 0 79568 800 79688 6 pcpi_rs1[18]
port 313 nsew signal output
rlabel metal2 s 54758 156455 54814 157255 6 pcpi_rs1[19]
port 314 nsew signal output
rlabel metal3 s 0 105408 800 105528 6 pcpi_rs1[1]
port 315 nsew signal output
rlabel metal2 s 99378 0 99434 800 6 pcpi_rs1[20]
port 316 nsew signal output
rlabel metal2 s 26698 156455 26754 157255 6 pcpi_rs1[21]
port 317 nsew signal output
rlabel metal3 s 154311 142808 155111 142928 6 pcpi_rs1[22]
port 318 nsew signal output
rlabel metal3 s 154311 27888 155111 28008 6 pcpi_rs1[23]
port 319 nsew signal output
rlabel metal2 s 130198 156455 130254 157255 6 pcpi_rs1[24]
port 320 nsew signal output
rlabel metal2 s 113638 0 113694 800 6 pcpi_rs1[25]
port 321 nsew signal output
rlabel metal2 s 84198 0 84254 800 6 pcpi_rs1[26]
port 322 nsew signal output
rlabel metal2 s 99378 156455 99434 157255 6 pcpi_rs1[27]
port 323 nsew signal output
rlabel metal2 s 110878 0 110934 800 6 pcpi_rs1[28]
port 324 nsew signal output
rlabel metal2 s 25778 0 25834 800 6 pcpi_rs1[29]
port 325 nsew signal output
rlabel metal2 s 9218 0 9274 800 6 pcpi_rs1[2]
port 326 nsew signal output
rlabel metal2 s 42338 0 42394 800 6 pcpi_rs1[30]
port 327 nsew signal output
rlabel metal2 s 95698 156455 95754 157255 6 pcpi_rs1[31]
port 328 nsew signal output
rlabel metal3 s 154311 116288 155111 116408 6 pcpi_rs1[3]
port 329 nsew signal output
rlabel metal3 s 154311 71408 155111 71528 6 pcpi_rs1[4]
port 330 nsew signal output
rlabel metal3 s 0 156408 800 156528 6 pcpi_rs1[5]
port 331 nsew signal output
rlabel metal2 s 93398 0 93454 800 6 pcpi_rs1[6]
port 332 nsew signal output
rlabel metal3 s 154311 74808 155111 74928 6 pcpi_rs1[7]
port 333 nsew signal output
rlabel metal3 s 154311 6808 155111 6928 6 pcpi_rs1[8]
port 334 nsew signal output
rlabel metal2 s 39578 0 39634 800 6 pcpi_rs1[9]
port 335 nsew signal output
rlabel metal2 s 86498 156455 86554 157255 6 pcpi_rs2[0]
port 336 nsew signal output
rlabel metal2 s 22098 0 22154 800 6 pcpi_rs2[10]
port 337 nsew signal output
rlabel metal3 s 154311 59848 155111 59968 6 pcpi_rs2[11]
port 338 nsew signal output
rlabel metal3 s 154311 99288 155111 99408 6 pcpi_rs2[12]
port 339 nsew signal output
rlabel metal2 s 138938 156455 138994 157255 6 pcpi_rs2[13]
port 340 nsew signal output
rlabel metal2 s 152738 156455 152794 157255 6 pcpi_rs2[14]
port 341 nsew signal output
rlabel metal3 s 154311 138728 155111 138848 6 pcpi_rs2[15]
port 342 nsew signal output
rlabel metal2 s 131118 156455 131174 157255 6 pcpi_rs2[16]
port 343 nsew signal output
rlabel metal2 s 79138 156455 79194 157255 6 pcpi_rs2[17]
port 344 nsew signal output
rlabel metal2 s 10598 0 10654 800 6 pcpi_rs2[18]
port 345 nsew signal output
rlabel metal3 s 0 65968 800 66088 6 pcpi_rs2[19]
port 346 nsew signal output
rlabel metal2 s 91558 156455 91614 157255 6 pcpi_rs2[1]
port 347 nsew signal output
rlabel metal2 s 14278 156455 14334 157255 6 pcpi_rs2[20]
port 348 nsew signal output
rlabel metal2 s 10138 156455 10194 157255 6 pcpi_rs2[21]
port 349 nsew signal output
rlabel metal2 s 63958 0 64014 800 6 pcpi_rs2[22]
port 350 nsew signal output
rlabel metal3 s 154311 72768 155111 72888 6 pcpi_rs2[23]
port 351 nsew signal output
rlabel metal2 s 105818 0 105874 800 6 pcpi_rs2[24]
port 352 nsew signal output
rlabel metal2 s 140318 0 140374 800 6 pcpi_rs2[25]
port 353 nsew signal output
rlabel metal3 s 0 87048 800 87168 6 pcpi_rs2[26]
port 354 nsew signal output
rlabel metal3 s 0 122408 800 122528 6 pcpi_rs2[27]
port 355 nsew signal output
rlabel metal3 s 154311 80248 155111 80368 6 pcpi_rs2[28]
port 356 nsew signal output
rlabel metal2 s 17958 0 18014 800 6 pcpi_rs2[29]
port 357 nsew signal output
rlabel metal3 s 154311 155728 155111 155848 6 pcpi_rs2[2]
port 358 nsew signal output
rlabel metal2 s 128818 156455 128874 157255 6 pcpi_rs2[30]
port 359 nsew signal output
rlabel metal2 s 117318 156455 117374 157255 6 pcpi_rs2[31]
port 360 nsew signal output
rlabel metal2 s 149058 156455 149114 157255 6 pcpi_rs2[3]
port 361 nsew signal output
rlabel metal3 s 0 11568 800 11688 6 pcpi_rs2[4]
port 362 nsew signal output
rlabel metal2 s 142618 156455 142674 157255 6 pcpi_rs2[5]
port 363 nsew signal output
rlabel metal3 s 0 9528 800 9648 6 pcpi_rs2[6]
port 364 nsew signal output
rlabel metal2 s 58898 0 58954 800 6 pcpi_rs2[7]
port 365 nsew signal output
rlabel metal2 s 62578 0 62634 800 6 pcpi_rs2[8]
port 366 nsew signal output
rlabel metal2 s 122378 156455 122434 157255 6 pcpi_rs2[9]
port 367 nsew signal output
rlabel metal2 s 25778 156455 25834 157255 6 pcpi_valid
port 368 nsew signal output
rlabel metal3 s 0 154368 800 154488 6 pcpi_wait
port 369 nsew signal input
rlabel metal2 s 75458 0 75514 800 6 pcpi_wr
port 370 nsew signal input
rlabel metal2 s 48778 0 48834 800 6 resetn
port 371 nsew signal input
rlabel metal2 s 122378 0 122434 800 6 trace_data[0]
port 372 nsew signal output
rlabel metal2 s 79138 0 79194 800 6 trace_data[10]
port 373 nsew signal output
rlabel metal2 s 87878 0 87934 800 6 trace_data[11]
port 374 nsew signal output
rlabel metal2 s 154118 0 154174 800 6 trace_data[12]
port 375 nsew signal output
rlabel metal3 s 0 21088 800 21208 6 trace_data[13]
port 376 nsew signal output
rlabel metal2 s 4158 156455 4214 157255 6 trace_data[14]
port 377 nsew signal output
rlabel metal2 s 64878 156455 64934 157255 6 trace_data[15]
port 378 nsew signal output
rlabel metal2 s 145378 156455 145434 157255 6 trace_data[16]
port 379 nsew signal output
rlabel metal2 s 57518 0 57574 800 6 trace_data[17]
port 380 nsew signal output
rlabel metal2 s 66258 156455 66314 157255 6 trace_data[18]
port 381 nsew signal output
rlabel metal2 s 125138 0 125194 800 6 trace_data[19]
port 382 nsew signal output
rlabel metal3 s 154311 65288 155111 65408 6 trace_data[1]
port 383 nsew signal output
rlabel metal2 s 43718 0 43774 800 6 trace_data[20]
port 384 nsew signal output
rlabel metal2 s 110878 156455 110934 157255 6 trace_data[21]
port 385 nsew signal output
rlabel metal3 s 0 138048 800 138168 6 trace_data[22]
port 386 nsew signal output
rlabel metal2 s 40958 156455 41014 157255 6 trace_data[23]
port 387 nsew signal output
rlabel metal3 s 0 62568 800 62688 6 trace_data[24]
port 388 nsew signal output
rlabel metal2 s 104438 156455 104494 157255 6 trace_data[25]
port 389 nsew signal output
rlabel metal3 s 0 2048 800 2168 6 trace_data[26]
port 390 nsew signal output
rlabel metal3 s 0 60528 800 60648 6 trace_data[27]
port 391 nsew signal output
rlabel metal3 s 0 90448 800 90568 6 trace_data[28]
port 392 nsew signal output
rlabel metal2 s 2778 0 2834 800 6 trace_data[29]
port 393 nsew signal output
rlabel metal2 s 118698 156455 118754 157255 6 trace_data[2]
port 394 nsew signal output
rlabel metal3 s 154311 146208 155111 146328 6 trace_data[30]
port 395 nsew signal output
rlabel metal2 s 109958 0 110014 800 6 trace_data[31]
port 396 nsew signal output
rlabel metal2 s 137558 0 137614 800 6 trace_data[32]
port 397 nsew signal output
rlabel metal2 s 53378 156455 53434 157255 6 trace_data[33]
port 398 nsew signal output
rlabel metal2 s 30838 0 30894 800 6 trace_data[34]
port 399 nsew signal output
rlabel metal2 s 128818 0 128874 800 6 trace_data[35]
port 400 nsew signal output
rlabel metal2 s 15658 0 15714 800 6 trace_data[3]
port 401 nsew signal output
rlabel metal3 s 154311 136688 155111 136808 6 trace_data[4]
port 402 nsew signal output
rlabel metal3 s 154311 29928 155111 30048 6 trace_data[5]
port 403 nsew signal output
rlabel metal2 s 29458 0 29514 800 6 trace_data[6]
port 404 nsew signal output
rlabel metal2 s 44638 0 44694 800 6 trace_data[7]
port 405 nsew signal output
rlabel metal2 s 123758 0 123814 800 6 trace_data[8]
port 406 nsew signal output
rlabel metal2 s 154118 156455 154174 157255 6 trace_data[9]
port 407 nsew signal output
rlabel metal2 s 35898 156455 35954 157255 6 trace_valid
port 408 nsew signal output
rlabel metal3 s 0 24488 800 24608 6 trap
port 409 nsew signal output
rlabel metal4 s 127088 2128 127408 155088 6 VPWR
port 410 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 155088 6 VPWR
port 411 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 155088 6 VPWR
port 412 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 155088 6 VPWR
port 413 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 155088 6 VPWR
port 414 nsew power bidirectional
rlabel metal5 s 1104 127842 153916 128162 6 VPWR
port 415 nsew power bidirectional
rlabel metal5 s 1104 97206 153916 97526 6 VPWR
port 416 nsew power bidirectional
rlabel metal5 s 1104 66570 153916 66890 6 VPWR
port 417 nsew power bidirectional
rlabel metal5 s 1104 35934 153916 36254 6 VPWR
port 418 nsew power bidirectional
rlabel metal5 s 1104 5298 153916 5618 6 VPWR
port 419 nsew power bidirectional
rlabel metal4 s 142448 2128 142768 155088 6 VGND
port 420 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 155088 6 VGND
port 421 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 155088 6 VGND
port 422 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 155088 6 VGND
port 423 nsew ground bidirectional
rlabel metal4 s 19568 2128 19888 155088 6 VGND
port 424 nsew ground bidirectional
rlabel metal5 s 1104 143160 153916 143480 6 VGND
port 425 nsew ground bidirectional
rlabel metal5 s 1104 112524 153916 112844 6 VGND
port 426 nsew ground bidirectional
rlabel metal5 s 1104 81888 153916 82208 6 VGND
port 427 nsew ground bidirectional
rlabel metal5 s 1104 51252 153916 51572 6 VGND
port 428 nsew ground bidirectional
rlabel metal5 s 1104 20616 153916 20936 6 VGND
port 429 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 155111 157255
string LEFview TRUE
string GDS_FILE /openLANE_flow/designs/picorv32a/runs/05-07_15-00/results/magic/picorv32a.gds
string GDS_END 66454588
string GDS_START 577774
<< end >>

