module picorv32a (clk,
    mem_instr,
    mem_la_read,
    mem_la_write,
    mem_ready,
    mem_valid,
    pcpi_ready,
    pcpi_valid,
    pcpi_wait,
    pcpi_wr,
    resetn,
    trace_valid,
    trap,
    eoi,
    irq,
    mem_addr,
    mem_la_addr,
    mem_la_wdata,
    mem_la_wstrb,
    mem_rdata,
    mem_wdata,
    mem_wstrb,
    pcpi_insn,
    pcpi_rd,
    pcpi_rs1,
    pcpi_rs2,
    trace_data);
 input clk;
 output mem_instr;
 output mem_la_read;
 output mem_la_write;
 input mem_ready;
 output mem_valid;
 input pcpi_ready;
 output pcpi_valid;
 input pcpi_wait;
 input pcpi_wr;
 input resetn;
 output trace_valid;
 output trap;
 output [31:0] eoi;
 input [31:0] irq;
 output [31:0] mem_addr;
 output [31:0] mem_la_addr;
 output [31:0] mem_la_wdata;
 output [3:0] mem_la_wstrb;
 input [31:0] mem_rdata;
 output [31:0] mem_wdata;
 output [3:0] mem_wstrb;
 output [31:0] pcpi_insn;
 input [31:0] pcpi_rd;
 output [31:0] pcpi_rs1;
 output [31:0] pcpi_rs2;
 output [35:0] trace_data;

 sky130_fd_sc_hd__inv_2 _20671_ (.A(mem_valid),
    .Y(_18005_));
 sky130_fd_sc_hd__inv_2 _20672_ (.A(mem_ready),
    .Y(_18006_));
 sky130_fd_sc_hd__nor2_2 _20673_ (.A(_18005_),
    .B(_18006_),
    .Y(_18007_));
 sky130_fd_sc_hd__inv_2 _20674_ (.A(_18007_),
    .Y(_18008_));
 sky130_fd_sc_hd__nand2_2 _20675_ (.A(\mem_state[1] ),
    .B(\mem_state[0] ),
    .Y(_18009_));
 sky130_fd_sc_hd__nor2_2 _20676_ (.A(\mem_state[1] ),
    .B(\mem_state[0] ),
    .Y(_00290_));
 sky130_fd_sc_hd__a21oi_2 _20677_ (.A1(_18008_),
    .A2(_18009_),
    .B1(_00290_),
    .Y(_18010_));
 sky130_fd_sc_hd__nor2_2 _20678_ (.A(mem_do_wdata),
    .B(mem_do_rdata),
    .Y(_18011_));
 sky130_fd_sc_hd__inv_2 _20679_ (.A(mem_do_rinst),
    .Y(_18012_));
 sky130_fd_sc_hd__o21ai_2 _20680_ (.A1(_18011_),
    .A2(_18008_),
    .B1(_18012_),
    .Y(_18013_));
 sky130_fd_sc_hd__nand2_2 _20681_ (.A(_18010_),
    .B(_18013_),
    .Y(_18014_));
 sky130_fd_sc_hd__buf_1 _20682_ (.A(mem_do_prefetch),
    .X(_18015_));
 sky130_fd_sc_hd__inv_2 _20683_ (.A(resetn),
    .Y(_18016_));
 sky130_fd_sc_hd__buf_1 _20684_ (.A(_18016_),
    .X(_18017_));
 sky130_fd_sc_hd__a21oi_2 _20685_ (.A1(_18014_),
    .A2(_18015_),
    .B1(_18017_),
    .Y(_18018_));
 sky130_fd_sc_hd__inv_2 _20686_ (.A(mem_do_rdata),
    .Y(_18019_));
 sky130_fd_sc_hd__inv_2 _20687_ (.A(\cpu_state[6] ),
    .Y(_18020_));
 sky130_fd_sc_hd__nor2_2 _20688_ (.A(_18019_),
    .B(_18020_),
    .Y(_00319_));
 sky130_fd_sc_hd__nand2_2 _20689_ (.A(_18018_),
    .B(_00319_),
    .Y(_18021_));
 sky130_fd_sc_hd__inv_2 _20690_ (.A(_18021_),
    .Y(_18022_));
 sky130_fd_sc_hd__nor2_2 _20691_ (.A(_00332_),
    .B(_18022_),
    .Y(_18023_));
 sky130_fd_sc_hd__buf_1 _20692_ (.A(resetn),
    .X(_18024_));
 sky130_fd_sc_hd__buf_1 _20693_ (.A(_18024_),
    .X(_18025_));
 sky130_fd_sc_hd__buf_1 _20694_ (.A(_18025_),
    .X(_18026_));
 sky130_fd_sc_hd__buf_1 _20695_ (.A(_18026_),
    .X(_18027_));
 sky130_fd_sc_hd__buf_1 _20696_ (.A(_18027_),
    .X(_18028_));
 sky130_fd_sc_hd__buf_1 _20697_ (.A(\cpu_state[6] ),
    .X(_18029_));
 sky130_fd_sc_hd__inv_2 _20698_ (.A(_18023_),
    .Y(_18030_));
 sky130_fd_sc_hd__a21o_2 _20699_ (.A1(instr_lb),
    .A2(_18029_),
    .B1(_18030_),
    .X(_18031_));
 sky130_fd_sc_hd__o211a_2 _20700_ (.A1(latched_is_lb),
    .A2(_18023_),
    .B1(_18028_),
    .C1(_18031_),
    .X(_04071_));
 sky130_fd_sc_hd__a21o_2 _20701_ (.A1(instr_lh),
    .A2(_18029_),
    .B1(_18030_),
    .X(_18032_));
 sky130_fd_sc_hd__o211a_2 _20702_ (.A1(latched_is_lh),
    .A2(_18023_),
    .B1(_18028_),
    .C1(_18032_),
    .X(_04070_));
 sky130_fd_sc_hd__inv_2 _20703_ (.A(instr_retirq),
    .Y(_18033_));
 sky130_fd_sc_hd__nand2_2 _20704_ (.A(_18033_),
    .B(\cpu_state[2] ),
    .Y(_18034_));
 sky130_fd_sc_hd__inv_2 _20705_ (.A(_00331_),
    .Y(_18035_));
 sky130_fd_sc_hd__nand2_2 _20706_ (.A(_18034_),
    .B(_18035_),
    .Y(_18036_));
 sky130_fd_sc_hd__inv_2 _20707_ (.A(latched_branch),
    .Y(_18037_));
 sky130_fd_sc_hd__nand2_2 _20708_ (.A(_18036_),
    .B(_18037_),
    .Y(_18038_));
 sky130_fd_sc_hd__o211a_2 _20709_ (.A1(_20620_),
    .A2(_18036_),
    .B1(_18028_),
    .C1(_18038_),
    .X(_04069_));
 sky130_fd_sc_hd__inv_2 _20710_ (.A(\mem_state[0] ),
    .Y(_18039_));
 sky130_fd_sc_hd__inv_2 _20711_ (.A(\mem_state[1] ),
    .Y(_18040_));
 sky130_fd_sc_hd__nor2_2 _20712_ (.A(_18039_),
    .B(_18012_),
    .Y(_18041_));
 sky130_fd_sc_hd__a211o_2 _20713_ (.A1(_18007_),
    .A2(_18039_),
    .B1(_18040_),
    .C1(_18041_),
    .X(_18042_));
 sky130_fd_sc_hd__nor2_2 _20714_ (.A(mem_do_rinst),
    .B(mem_do_prefetch),
    .Y(_18043_));
 sky130_fd_sc_hd__nand2_2 _20715_ (.A(_18011_),
    .B(_18043_),
    .Y(_18044_));
 sky130_fd_sc_hd__inv_2 _20716_ (.A(_00290_),
    .Y(_18045_));
 sky130_fd_sc_hd__or2_2 _20717_ (.A(_18044_),
    .B(_18045_),
    .X(_18046_));
 sky130_fd_sc_hd__inv_2 _20718_ (.A(trap),
    .Y(_18047_));
 sky130_fd_sc_hd__buf_1 _20719_ (.A(_18017_),
    .X(_18048_));
 sky130_fd_sc_hd__a31o_2 _20720_ (.A1(_18042_),
    .A2(_18046_),
    .A3(_18047_),
    .B1(_18048_),
    .X(_18049_));
 sky130_fd_sc_hd__and2_2 _20721_ (.A(_18049_),
    .B(_00300_),
    .X(_18050_));
 sky130_fd_sc_hd__buf_1 _20722_ (.A(_18017_),
    .X(_18051_));
 sky130_fd_sc_hd__nor2_2 _20723_ (.A(trap),
    .B(_18051_),
    .Y(_18052_));
 sky130_fd_sc_hd__buf_1 _20724_ (.A(_18052_),
    .X(_18053_));
 sky130_fd_sc_hd__nor2_2 _20725_ (.A(_18040_),
    .B(_18050_),
    .Y(_18054_));
 sky130_fd_sc_hd__a31o_2 _20726_ (.A1(_20585_),
    .A2(_18050_),
    .A3(_18053_),
    .B1(_18054_),
    .X(_04068_));
 sky130_fd_sc_hd__nor2_2 _20727_ (.A(_18039_),
    .B(_18050_),
    .Y(_18055_));
 sky130_fd_sc_hd__a31o_2 _20728_ (.A1(_20584_),
    .A2(_18050_),
    .A3(_18053_),
    .B1(_18055_),
    .X(_04067_));
 sky130_fd_sc_hd__nor2_2 _20729_ (.A(_18016_),
    .B(_18014_),
    .Y(_18056_));
 sky130_fd_sc_hd__inv_2 _20730_ (.A(_18056_),
    .Y(_18057_));
 sky130_fd_sc_hd__nor2_2 _20731_ (.A(_18012_),
    .B(_18057_),
    .Y(_18058_));
 sky130_fd_sc_hd__buf_1 _20732_ (.A(_18058_),
    .X(_18059_));
 sky130_fd_sc_hd__buf_1 _20733_ (.A(_18059_),
    .X(_20587_));
 sky130_fd_sc_hd__inv_2 _20734_ (.A(\decoded_rs1[4] ),
    .Y(_00366_));
 sky130_fd_sc_hd__buf_1 _20735_ (.A(_18058_),
    .X(_18060_));
 sky130_fd_sc_hd__buf_1 _20736_ (.A(_18060_),
    .X(_18061_));
 sky130_fd_sc_hd__and3b_2 _20737_ (.A_N(_00326_),
    .B(_00325_),
    .C(_00324_),
    .X(_18062_));
 sky130_fd_sc_hd__inv_2 _20738_ (.A(_00330_),
    .Y(_18063_));
 sky130_fd_sc_hd__inv_2 _20739_ (.A(_00327_),
    .Y(_18064_));
 sky130_fd_sc_hd__nor2_2 _20740_ (.A(\mem_rdata_latched[28] ),
    .B(_18064_),
    .Y(_18065_));
 sky130_fd_sc_hd__nor2_2 _20741_ (.A(_00329_),
    .B(_00328_),
    .Y(_18066_));
 sky130_fd_sc_hd__and4_2 _20742_ (.A(_18062_),
    .B(_18063_),
    .C(_18065_),
    .D(_18066_),
    .X(_18067_));
 sky130_fd_sc_hd__inv_2 _20743_ (.A(\mem_rdata_latched[27] ),
    .Y(_18068_));
 sky130_fd_sc_hd__nor3_2 _20744_ (.A(\mem_rdata_latched[31] ),
    .B(\mem_rdata_latched[30] ),
    .C(\mem_rdata_latched[29] ),
    .Y(_18069_));
 sky130_fd_sc_hd__inv_2 _20745_ (.A(\mem_rdata_latched[25] ),
    .Y(_18070_));
 sky130_fd_sc_hd__and3_2 _20746_ (.A(_18069_),
    .B(\mem_rdata_latched[26] ),
    .C(_18070_),
    .X(_18071_));
 sky130_fd_sc_hd__and3_2 _20747_ (.A(_18067_),
    .B(_18068_),
    .C(_18071_),
    .X(_18072_));
 sky130_fd_sc_hd__buf_1 _20748_ (.A(_18072_),
    .X(_18073_));
 sky130_fd_sc_hd__nand2_2 _20749_ (.A(_18059_),
    .B(_18073_),
    .Y(_18074_));
 sky130_fd_sc_hd__and3b_2 _20750_ (.A_N(\mem_rdata_latched[26] ),
    .B(_18069_),
    .C(_18070_),
    .X(_18075_));
 sky130_fd_sc_hd__and3_2 _20751_ (.A(_18067_),
    .B(_18068_),
    .C(_18075_),
    .X(_18076_));
 sky130_fd_sc_hd__buf_1 _20752_ (.A(_18059_),
    .X(_18077_));
 sky130_fd_sc_hd__o21ai_2 _20753_ (.A1(\mem_rdata_latched[19] ),
    .A2(_18076_),
    .B1(_18077_),
    .Y(_18078_));
 sky130_fd_sc_hd__o211ai_2 _20754_ (.A1(_00366_),
    .A2(_18061_),
    .B1(_18074_),
    .C1(_18078_),
    .Y(_04066_));
 sky130_fd_sc_hd__nand2_2 _20755_ (.A(\cpu_state[1] ),
    .B(decoder_trigger),
    .Y(_18079_));
 sky130_fd_sc_hd__inv_2 _20756_ (.A(decoder_trigger),
    .Y(_18080_));
 sky130_fd_sc_hd__inv_2 _20757_ (.A(\irq_mask[2] ),
    .Y(_18081_));
 sky130_fd_sc_hd__inv_2 _20758_ (.A(\irq_pending[0] ),
    .Y(_18082_));
 sky130_fd_sc_hd__nor2_2 _20759_ (.A(\irq_mask[0] ),
    .B(_18082_),
    .Y(_18083_));
 sky130_fd_sc_hd__inv_2 _20760_ (.A(\irq_pending[1] ),
    .Y(_18084_));
 sky130_fd_sc_hd__nor2_2 _20761_ (.A(\irq_mask[1] ),
    .B(_18084_),
    .Y(_18085_));
 sky130_fd_sc_hd__inv_2 _20762_ (.A(\irq_mask[3] ),
    .Y(_18086_));
 sky130_fd_sc_hd__and2_2 _20763_ (.A(_18086_),
    .B(\irq_pending[3] ),
    .X(_18087_));
 sky130_fd_sc_hd__a2111o_2 _20764_ (.A1(_18081_),
    .A2(\irq_pending[2] ),
    .B1(_18083_),
    .C1(_18085_),
    .D1(_18087_),
    .X(_18088_));
 sky130_fd_sc_hd__inv_2 _20765_ (.A(\irq_mask[17] ),
    .Y(_18089_));
 sky130_fd_sc_hd__inv_2 _20766_ (.A(\irq_pending[16] ),
    .Y(_18090_));
 sky130_fd_sc_hd__nor2_2 _20767_ (.A(\irq_mask[16] ),
    .B(_18090_),
    .Y(_18091_));
 sky130_fd_sc_hd__inv_2 _20768_ (.A(\irq_mask[19] ),
    .Y(_18092_));
 sky130_fd_sc_hd__and2_2 _20769_ (.A(_18092_),
    .B(\irq_pending[19] ),
    .X(_18093_));
 sky130_fd_sc_hd__inv_2 _20770_ (.A(\irq_mask[18] ),
    .Y(_18094_));
 sky130_fd_sc_hd__and2_2 _20771_ (.A(_18094_),
    .B(\irq_pending[18] ),
    .X(_18095_));
 sky130_fd_sc_hd__a2111o_2 _20772_ (.A1(_18089_),
    .A2(\irq_pending[17] ),
    .B1(_18091_),
    .C1(_18093_),
    .D1(_18095_),
    .X(_18096_));
 sky130_fd_sc_hd__and2b_2 _20773_ (.A_N(\irq_mask[27] ),
    .B(\irq_pending[27] ),
    .X(_18097_));
 sky130_fd_sc_hd__and2b_2 _20774_ (.A_N(\irq_mask[26] ),
    .B(\irq_pending[26] ),
    .X(_18098_));
 sky130_fd_sc_hd__inv_2 _20775_ (.A(\irq_mask[25] ),
    .Y(_18099_));
 sky130_fd_sc_hd__inv_2 _20776_ (.A(\irq_mask[24] ),
    .Y(_18100_));
 sky130_fd_sc_hd__a22o_2 _20777_ (.A1(_18099_),
    .A2(\irq_pending[25] ),
    .B1(_18100_),
    .B2(\irq_pending[24] ),
    .X(_18101_));
 sky130_fd_sc_hd__or3_2 _20778_ (.A(_18097_),
    .B(_18098_),
    .C(_18101_),
    .X(_18102_));
 sky130_fd_sc_hd__inv_2 _20779_ (.A(\irq_mask[23] ),
    .Y(_18103_));
 sky130_fd_sc_hd__and2_2 _20780_ (.A(_18103_),
    .B(\irq_pending[23] ),
    .X(_18104_));
 sky130_fd_sc_hd__inv_2 _20781_ (.A(\irq_mask[22] ),
    .Y(_18105_));
 sky130_fd_sc_hd__and2_2 _20782_ (.A(_18105_),
    .B(\irq_pending[22] ),
    .X(_18106_));
 sky130_fd_sc_hd__inv_2 _20783_ (.A(\irq_mask[21] ),
    .Y(_18107_));
 sky130_fd_sc_hd__inv_2 _20784_ (.A(\irq_mask[20] ),
    .Y(_18108_));
 sky130_fd_sc_hd__a22o_2 _20785_ (.A1(_18107_),
    .A2(\irq_pending[21] ),
    .B1(_18108_),
    .B2(\irq_pending[20] ),
    .X(_18109_));
 sky130_fd_sc_hd__or3_2 _20786_ (.A(_18104_),
    .B(_18106_),
    .C(_18109_),
    .X(_18110_));
 sky130_fd_sc_hd__or4_2 _20787_ (.A(_18088_),
    .B(_18096_),
    .C(_18102_),
    .D(_18110_),
    .X(_18111_));
 sky130_fd_sc_hd__and2b_2 _20788_ (.A_N(\irq_mask[11] ),
    .B(\irq_pending[11] ),
    .X(_18112_));
 sky130_fd_sc_hd__and2b_2 _20789_ (.A_N(\irq_mask[10] ),
    .B(\irq_pending[10] ),
    .X(_18113_));
 sky130_fd_sc_hd__inv_2 _20790_ (.A(\irq_mask[9] ),
    .Y(_18114_));
 sky130_fd_sc_hd__inv_2 _20791_ (.A(\irq_mask[8] ),
    .Y(_18115_));
 sky130_fd_sc_hd__a22o_2 _20792_ (.A1(_18114_),
    .A2(\irq_pending[9] ),
    .B1(_18115_),
    .B2(\irq_pending[8] ),
    .X(_18116_));
 sky130_fd_sc_hd__or3_2 _20793_ (.A(_18112_),
    .B(_18113_),
    .C(_18116_),
    .X(_18117_));
 sky130_fd_sc_hd__inv_2 _20794_ (.A(\irq_mask[7] ),
    .Y(_18118_));
 sky130_fd_sc_hd__and2_2 _20795_ (.A(_18118_),
    .B(\irq_pending[7] ),
    .X(_18119_));
 sky130_fd_sc_hd__inv_2 _20796_ (.A(\irq_mask[6] ),
    .Y(_18120_));
 sky130_fd_sc_hd__and2_2 _20797_ (.A(_18120_),
    .B(\irq_pending[6] ),
    .X(_18121_));
 sky130_fd_sc_hd__inv_2 _20798_ (.A(\irq_mask[5] ),
    .Y(_18122_));
 sky130_fd_sc_hd__inv_2 _20799_ (.A(\irq_mask[4] ),
    .Y(_18123_));
 sky130_fd_sc_hd__a22o_2 _20800_ (.A1(_18122_),
    .A2(\irq_pending[5] ),
    .B1(_18123_),
    .B2(\irq_pending[4] ),
    .X(_18124_));
 sky130_fd_sc_hd__or3_2 _20801_ (.A(_18119_),
    .B(_18121_),
    .C(_18124_),
    .X(_18125_));
 sky130_fd_sc_hd__inv_2 _20802_ (.A(\irq_mask[29] ),
    .Y(_18126_));
 sky130_fd_sc_hd__inv_2 _20803_ (.A(\irq_mask[28] ),
    .Y(_18127_));
 sky130_fd_sc_hd__and2_2 _20804_ (.A(_18127_),
    .B(\irq_pending[28] ),
    .X(_18128_));
 sky130_fd_sc_hd__inv_2 _20805_ (.A(\irq_mask[31] ),
    .Y(_18129_));
 sky130_fd_sc_hd__and2_2 _20806_ (.A(_18129_),
    .B(\irq_pending[31] ),
    .X(_18130_));
 sky130_fd_sc_hd__inv_2 _20807_ (.A(\irq_mask[30] ),
    .Y(_18131_));
 sky130_fd_sc_hd__and2_2 _20808_ (.A(_18131_),
    .B(\irq_pending[30] ),
    .X(_18132_));
 sky130_fd_sc_hd__a2111o_2 _20809_ (.A1(_18126_),
    .A2(\irq_pending[29] ),
    .B1(_18128_),
    .C1(_18130_),
    .D1(_18132_),
    .X(_18133_));
 sky130_fd_sc_hd__inv_2 _20810_ (.A(\irq_mask[13] ),
    .Y(_18134_));
 sky130_fd_sc_hd__inv_2 _20811_ (.A(\irq_mask[12] ),
    .Y(_18135_));
 sky130_fd_sc_hd__and2_2 _20812_ (.A(_18135_),
    .B(\irq_pending[12] ),
    .X(_18136_));
 sky130_fd_sc_hd__inv_2 _20813_ (.A(\irq_mask[15] ),
    .Y(_18137_));
 sky130_fd_sc_hd__and2_2 _20814_ (.A(_18137_),
    .B(\irq_pending[15] ),
    .X(_18138_));
 sky130_fd_sc_hd__inv_2 _20815_ (.A(\irq_mask[14] ),
    .Y(_18139_));
 sky130_fd_sc_hd__and2_2 _20816_ (.A(_18139_),
    .B(\irq_pending[14] ),
    .X(_18140_));
 sky130_fd_sc_hd__a2111o_2 _20817_ (.A1(_18134_),
    .A2(\irq_pending[13] ),
    .B1(_18136_),
    .C1(_18138_),
    .D1(_18140_),
    .X(_18141_));
 sky130_fd_sc_hd__or4_2 _20818_ (.A(_18117_),
    .B(_18125_),
    .C(_18133_),
    .D(_18141_),
    .X(_18142_));
 sky130_fd_sc_hd__nor2_2 _20819_ (.A(_18111_),
    .B(_18142_),
    .Y(_18143_));
 sky130_fd_sc_hd__or4_2 _20820_ (.A(irq_active),
    .B(irq_delay),
    .C(_18080_),
    .D(_18143_),
    .X(_18144_));
 sky130_fd_sc_hd__nor2_2 _20821_ (.A(\irq_state[1] ),
    .B(\irq_state[0] ),
    .Y(_18145_));
 sky130_fd_sc_hd__nand2_2 _20822_ (.A(_18144_),
    .B(_18145_),
    .Y(_18146_));
 sky130_fd_sc_hd__inv_2 _20823_ (.A(_18146_),
    .Y(_18147_));
 sky130_fd_sc_hd__inv_2 _20824_ (.A(instr_waitirq),
    .Y(_18148_));
 sky130_fd_sc_hd__nor2_2 _20825_ (.A(decoder_trigger),
    .B(do_waitirq),
    .Y(_18149_));
 sky130_fd_sc_hd__nor2_2 _20826_ (.A(_18148_),
    .B(_18149_),
    .Y(_00309_));
 sky130_fd_sc_hd__inv_2 _20827_ (.A(_00309_),
    .Y(_18150_));
 sky130_fd_sc_hd__nand2_2 _20828_ (.A(_18147_),
    .B(_18150_),
    .Y(_18151_));
 sky130_fd_sc_hd__or2_2 _20829_ (.A(_18079_),
    .B(_18151_),
    .X(_18152_));
 sky130_fd_sc_hd__inv_2 _20830_ (.A(_18152_),
    .Y(_18153_));
 sky130_fd_sc_hd__inv_2 _20831_ (.A(irq_active),
    .Y(_18154_));
 sky130_fd_sc_hd__nand2_2 _20832_ (.A(_18153_),
    .B(_18154_),
    .Y(_18155_));
 sky130_fd_sc_hd__o211a_2 _20833_ (.A1(irq_delay),
    .A2(_18153_),
    .B1(_18028_),
    .C1(_18155_),
    .X(_04065_));
 sky130_fd_sc_hd__buf_1 _20834_ (.A(\pcpi_mul.rs1[32] ),
    .X(_18156_));
 sky130_fd_sc_hd__buf_1 _20835_ (.A(_18156_),
    .X(_18157_));
 sky130_fd_sc_hd__buf_1 _20836_ (.A(_18157_),
    .X(_18158_));
 sky130_fd_sc_hd__nand2_2 _20837_ (.A(_18024_),
    .B(pcpi_valid),
    .Y(_18159_));
 sky130_fd_sc_hd__or4_2 _20838_ (.A(pcpi_insn[31]),
    .B(pcpi_insn[30]),
    .C(pcpi_insn[29]),
    .D(pcpi_insn[28]),
    .X(_18160_));
 sky130_fd_sc_hd__nor2_2 _20839_ (.A(_18159_),
    .B(_18160_),
    .Y(_18161_));
 sky130_fd_sc_hd__inv_2 _20840_ (.A(\pcpi_mul.active[0] ),
    .Y(_18162_));
 sky130_fd_sc_hd__inv_2 _20841_ (.A(\pcpi_mul.active[1] ),
    .Y(_18163_));
 sky130_fd_sc_hd__and3_2 _20842_ (.A(_18161_),
    .B(_18162_),
    .C(_18163_),
    .X(_18164_));
 sky130_fd_sc_hd__or3_2 _20843_ (.A(pcpi_insn[27]),
    .B(pcpi_insn[26]),
    .C(pcpi_insn[14]),
    .X(_18165_));
 sky130_fd_sc_hd__nor3b_2 _20844_ (.A(pcpi_insn[6]),
    .B(pcpi_insn[3]),
    .C_N(pcpi_insn[4]),
    .Y(_18166_));
 sky130_fd_sc_hd__and2_2 _20845_ (.A(_18166_),
    .B(pcpi_insn[5]),
    .X(_18167_));
 sky130_fd_sc_hd__and3b_2 _20846_ (.A_N(pcpi_insn[2]),
    .B(pcpi_insn[1]),
    .C(pcpi_insn[0]),
    .X(_18168_));
 sky130_fd_sc_hd__and4b_2 _20847_ (.A_N(_18165_),
    .B(_18167_),
    .C(pcpi_insn[25]),
    .D(_18168_),
    .X(_18169_));
 sky130_fd_sc_hd__nand2_2 _20848_ (.A(_18164_),
    .B(_18169_),
    .Y(_18170_));
 sky130_fd_sc_hd__buf_1 _20849_ (.A(_18170_),
    .X(_18171_));
 sky130_fd_sc_hd__buf_1 _20850_ (.A(_18171_),
    .X(_18172_));
 sky130_fd_sc_hd__inv_2 _20851_ (.A(pcpi_rs1[31]),
    .Y(_18173_));
 sky130_fd_sc_hd__buf_1 _20852_ (.A(_18170_),
    .X(_18174_));
 sky130_fd_sc_hd__buf_1 _20853_ (.A(_18174_),
    .X(_18175_));
 sky130_fd_sc_hd__nor2_2 _20854_ (.A(_18173_),
    .B(_18175_),
    .Y(_18176_));
 sky130_fd_sc_hd__nor2_2 _20855_ (.A(pcpi_insn[13]),
    .B(pcpi_insn[12]),
    .Y(_18177_));
 sky130_fd_sc_hd__and2_2 _20856_ (.A(pcpi_insn[13]),
    .B(pcpi_insn[12]),
    .X(_18178_));
 sky130_fd_sc_hd__nor2_2 _20857_ (.A(_18177_),
    .B(_18178_),
    .Y(_18179_));
 sky130_fd_sc_hd__a22o_2 _20858_ (.A1(_18158_),
    .A2(_18172_),
    .B1(_18176_),
    .B2(_18179_),
    .X(_04064_));
 sky130_fd_sc_hd__inv_2 _20859_ (.A(_18171_),
    .Y(_03728_));
 sky130_fd_sc_hd__and2b_2 _20860_ (.A_N(pcpi_insn[13]),
    .B(pcpi_insn[12]),
    .X(_18180_));
 sky130_fd_sc_hd__inv_2 _20861_ (.A(\pcpi_mul.rs2[32] ),
    .Y(_18181_));
 sky130_fd_sc_hd__buf_1 _20862_ (.A(_18181_),
    .X(_18182_));
 sky130_fd_sc_hd__buf_1 _20863_ (.A(_18182_),
    .X(_18183_));
 sky130_fd_sc_hd__buf_1 _20864_ (.A(_18183_),
    .X(_18184_));
 sky130_fd_sc_hd__nor2_2 _20865_ (.A(_18184_),
    .B(_03728_),
    .Y(_18185_));
 sky130_fd_sc_hd__a31o_2 _20866_ (.A1(pcpi_rs2[31]),
    .A2(_03728_),
    .A3(_18180_),
    .B1(_18185_),
    .X(_04063_));
 sky130_fd_sc_hd__inv_2 _20867_ (.A(\cpu_state[4] ),
    .Y(_18186_));
 sky130_fd_sc_hd__buf_1 _20868_ (.A(_18186_),
    .X(_18187_));
 sky130_fd_sc_hd__buf_1 _20869_ (.A(_18187_),
    .X(_18188_));
 sky130_fd_sc_hd__buf_1 _20870_ (.A(_18051_),
    .X(_18189_));
 sky130_fd_sc_hd__buf_1 _20871_ (.A(_18189_),
    .X(_18190_));
 sky130_fd_sc_hd__inv_2 _20872_ (.A(alu_wait),
    .Y(_00302_));
 sky130_fd_sc_hd__nand2_2 _20873_ (.A(_00302_),
    .B(is_beq_bne_blt_bge_bltu_bgeu),
    .Y(_18191_));
 sky130_fd_sc_hd__a21oi_2 _20874_ (.A1(_18191_),
    .A2(_00333_),
    .B1(latched_stalu),
    .Y(_18192_));
 sky130_fd_sc_hd__a211oi_2 _20875_ (.A1(_18188_),
    .A2(_00333_),
    .B1(_18190_),
    .C1(_18192_),
    .Y(_04062_));
 sky130_fd_sc_hd__inv_2 _20876_ (.A(\cpu_state[2] ),
    .Y(_18193_));
 sky130_fd_sc_hd__buf_1 _20877_ (.A(_18193_),
    .X(_18194_));
 sky130_fd_sc_hd__or4_2 _20878_ (.A(instr_rdinstrh),
    .B(instr_rdinstr),
    .C(instr_rdcycleh),
    .D(instr_rdcycle),
    .X(_18195_));
 sky130_fd_sc_hd__nor2_2 _20879_ (.A(instr_setq),
    .B(instr_getq),
    .Y(_18196_));
 sky130_fd_sc_hd__inv_2 _20880_ (.A(instr_timer),
    .Y(_18197_));
 sky130_fd_sc_hd__buf_1 _20881_ (.A(instr_maskirq),
    .X(_18198_));
 sky130_fd_sc_hd__inv_2 _20882_ (.A(_18198_),
    .Y(_18199_));
 sky130_fd_sc_hd__and4_2 _20883_ (.A(_18196_),
    .B(_18197_),
    .C(_18199_),
    .D(_18033_),
    .X(_01717_));
 sky130_fd_sc_hd__or2b_2 _20884_ (.A(_18195_),
    .B_N(_01717_),
    .X(_18200_));
 sky130_fd_sc_hd__nor2_2 _20885_ (.A(_18194_),
    .B(_18200_),
    .Y(_18201_));
 sky130_fd_sc_hd__nor2_2 _20886_ (.A(\cpu_state[4] ),
    .B(\cpu_state[2] ),
    .Y(_18202_));
 sky130_fd_sc_hd__inv_2 _20887_ (.A(_18202_),
    .Y(_02542_));
 sky130_fd_sc_hd__nor2_2 _20888_ (.A(\cpu_state[3] ),
    .B(_02542_),
    .Y(_00354_));
 sky130_fd_sc_hd__inv_2 _20889_ (.A(\cpu_state[1] ),
    .Y(_18203_));
 sky130_fd_sc_hd__buf_1 _20890_ (.A(_18203_),
    .X(_18204_));
 sky130_fd_sc_hd__buf_1 _20891_ (.A(_18020_),
    .X(_18205_));
 sky130_fd_sc_hd__buf_1 _20892_ (.A(\cpu_state[4] ),
    .X(_18206_));
 sky130_fd_sc_hd__a32o_2 _20893_ (.A1(_00354_),
    .A2(_18204_),
    .A3(_18205_),
    .B1(_18206_),
    .B2(alu_wait),
    .X(_18207_));
 sky130_fd_sc_hd__nand2_2 _20894_ (.A(_18196_),
    .B(_18033_),
    .Y(_18208_));
 sky130_fd_sc_hd__or4_2 _20895_ (.A(instr_xor),
    .B(instr_sltu),
    .C(instr_maskirq),
    .D(_18208_),
    .X(_18209_));
 sky130_fd_sc_hd__nor2_2 _20896_ (.A(instr_bgeu),
    .B(instr_bge),
    .Y(_18210_));
 sky130_fd_sc_hd__nor2_2 _20897_ (.A(instr_sltiu),
    .B(instr_slti),
    .Y(_18211_));
 sky130_fd_sc_hd__inv_2 _20898_ (.A(instr_and),
    .Y(_18212_));
 sky130_fd_sc_hd__inv_2 _20899_ (.A(instr_or),
    .Y(_18213_));
 sky130_fd_sc_hd__and4_2 _20900_ (.A(_18210_),
    .B(_18211_),
    .C(_18212_),
    .D(_18213_),
    .X(_18214_));
 sky130_fd_sc_hd__or3b_2 _20901_ (.A(_18195_),
    .B(_18209_),
    .C_N(_18214_),
    .X(_18215_));
 sky130_fd_sc_hd__or4_2 _20902_ (.A(instr_bltu),
    .B(instr_blt),
    .C(instr_bne),
    .D(instr_beq),
    .X(_18216_));
 sky130_fd_sc_hd__or4_2 _20903_ (.A(instr_sh),
    .B(instr_sb),
    .C(instr_lhu),
    .D(instr_lbu),
    .X(_18217_));
 sky130_fd_sc_hd__nor2_2 _20904_ (.A(instr_auipc),
    .B(instr_lui),
    .Y(_18218_));
 sky130_fd_sc_hd__inv_2 _20905_ (.A(instr_jal),
    .Y(_00323_));
 sky130_fd_sc_hd__nand2_2 _20906_ (.A(_18218_),
    .B(_00323_),
    .Y(_00005_));
 sky130_fd_sc_hd__or4_2 _20907_ (.A(instr_lw),
    .B(instr_lh),
    .C(instr_lb),
    .D(instr_jalr),
    .X(_18219_));
 sky130_fd_sc_hd__or4_2 _20908_ (.A(instr_sra),
    .B(instr_srl),
    .C(instr_srai),
    .D(instr_srli),
    .X(_18220_));
 sky130_fd_sc_hd__or3_2 _20909_ (.A(_00005_),
    .B(_18219_),
    .C(_18220_),
    .X(_18221_));
 sky130_fd_sc_hd__or4_2 _20910_ (.A(instr_andi),
    .B(instr_ori),
    .C(instr_xori),
    .D(instr_addi),
    .X(_18222_));
 sky130_fd_sc_hd__or4_2 _20911_ (.A(instr_slt),
    .B(instr_sll),
    .C(instr_sub),
    .D(instr_add),
    .X(_18223_));
 sky130_fd_sc_hd__or4_2 _20912_ (.A(instr_timer),
    .B(instr_waitirq),
    .C(instr_slli),
    .D(instr_sw),
    .X(_18224_));
 sky130_fd_sc_hd__or3_2 _20913_ (.A(_18222_),
    .B(_18223_),
    .C(_18224_),
    .X(_18225_));
 sky130_fd_sc_hd__or4_2 _20914_ (.A(_18216_),
    .B(_18217_),
    .C(_18221_),
    .D(_18225_),
    .X(_18226_));
 sky130_fd_sc_hd__nor2_2 _20915_ (.A(_18215_),
    .B(_18226_),
    .Y(_00310_));
 sky130_fd_sc_hd__inv_2 _20916_ (.A(\cpu_state[3] ),
    .Y(_18227_));
 sky130_fd_sc_hd__a21o_2 _20917_ (.A1(_00310_),
    .A2(\pcpi_mul.active[1] ),
    .B1(_18227_),
    .X(_18228_));
 sky130_fd_sc_hd__or3b_2 _20918_ (.A(_18201_),
    .B(_18207_),
    .C_N(_18228_),
    .X(_18229_));
 sky130_fd_sc_hd__inv_2 _20919_ (.A(latched_store),
    .Y(_18230_));
 sky130_fd_sc_hd__nand2_2 _20920_ (.A(_18229_),
    .B(_18230_),
    .Y(_18231_));
 sky130_fd_sc_hd__o211a_2 _20921_ (.A1(_20621_),
    .A2(_18229_),
    .B1(_18028_),
    .C1(_18231_),
    .X(_04061_));
 sky130_fd_sc_hd__inv_2 _20922_ (.A(\irq_state[0] ),
    .Y(_18232_));
 sky130_fd_sc_hd__or2_2 _20923_ (.A(\irq_state[1] ),
    .B(_18204_),
    .X(_18233_));
 sky130_fd_sc_hd__or2_2 _20924_ (.A(_18232_),
    .B(_18233_),
    .X(_18234_));
 sky130_fd_sc_hd__buf_1 _20925_ (.A(_18204_),
    .X(_18235_));
 sky130_fd_sc_hd__buf_1 _20926_ (.A(\irq_state[1] ),
    .X(_18236_));
 sky130_fd_sc_hd__nand2_2 _20927_ (.A(_18235_),
    .B(_18236_),
    .Y(_18237_));
 sky130_fd_sc_hd__buf_1 _20928_ (.A(_18051_),
    .X(_18238_));
 sky130_fd_sc_hd__buf_1 _20929_ (.A(_18238_),
    .X(_18239_));
 sky130_fd_sc_hd__a21oi_2 _20930_ (.A1(_18234_),
    .A2(_18237_),
    .B1(_18239_),
    .Y(_04060_));
 sky130_fd_sc_hd__buf_1 _20931_ (.A(\irq_state[0] ),
    .X(_18240_));
 sky130_fd_sc_hd__buf_1 _20932_ (.A(_18204_),
    .X(_18241_));
 sky130_fd_sc_hd__or4_2 _20933_ (.A(_18236_),
    .B(_18240_),
    .C(_18241_),
    .D(_18144_),
    .X(_18242_));
 sky130_fd_sc_hd__buf_1 _20934_ (.A(_18240_),
    .X(_18243_));
 sky130_fd_sc_hd__nand2_2 _20935_ (.A(_18235_),
    .B(_18243_),
    .Y(_18244_));
 sky130_fd_sc_hd__buf_1 _20936_ (.A(_18238_),
    .X(_18245_));
 sky130_fd_sc_hd__a21oi_2 _20937_ (.A1(_18242_),
    .A2(_18244_),
    .B1(_18245_),
    .Y(_04059_));
 sky130_fd_sc_hd__inv_2 _20938_ (.A(_00310_),
    .Y(_18246_));
 sky130_fd_sc_hd__a21o_2 _20939_ (.A1(is_sb_sh_sw),
    .A2(_18246_),
    .B1(_18228_),
    .X(_18247_));
 sky130_fd_sc_hd__nand2_2 _20940_ (.A(_00354_),
    .B(_18204_),
    .Y(_18248_));
 sky130_fd_sc_hd__nand2_2 _20941_ (.A(_18246_),
    .B(is_lb_lh_lw_lbu_lhu),
    .Y(_18249_));
 sky130_fd_sc_hd__buf_1 _20942_ (.A(\cpu_state[2] ),
    .X(_18250_));
 sky130_fd_sc_hd__nand2_2 _20943_ (.A(_18249_),
    .B(_18250_),
    .Y(_18251_));
 sky130_fd_sc_hd__nand2_2 _20944_ (.A(_00302_),
    .B(\cpu_state[4] ),
    .Y(_18252_));
 sky130_fd_sc_hd__and4_2 _20945_ (.A(_18247_),
    .B(_18248_),
    .C(_18251_),
    .D(_18252_),
    .X(_18253_));
 sky130_fd_sc_hd__nand2_2 _20946_ (.A(_18014_),
    .B(_18025_),
    .Y(_18254_));
 sky130_fd_sc_hd__nor2_2 _20947_ (.A(\cpu_state[6] ),
    .B(\cpu_state[5] ),
    .Y(_00297_));
 sky130_fd_sc_hd__inv_2 _20948_ (.A(_00297_),
    .Y(_18255_));
 sky130_fd_sc_hd__or2_2 _20949_ (.A(_18048_),
    .B(_18191_),
    .X(_18256_));
 sky130_fd_sc_hd__buf_1 _20950_ (.A(\cpu_state[3] ),
    .X(_18257_));
 sky130_fd_sc_hd__nor2_2 _20951_ (.A(\cpu_state[1] ),
    .B(\cpu_state[2] ),
    .Y(_00315_));
 sky130_fd_sc_hd__inv_2 _20952_ (.A(_00315_),
    .Y(_18258_));
 sky130_fd_sc_hd__or3_2 _20953_ (.A(\cpu_state[0] ),
    .B(_18257_),
    .C(_18258_),
    .X(_18259_));
 sky130_fd_sc_hd__or4_2 _20954_ (.A(_00343_),
    .B(_18255_),
    .C(_18256_),
    .D(_18259_),
    .X(_18260_));
 sky130_fd_sc_hd__or3b_2 _20955_ (.A(_00356_),
    .B(_18254_),
    .C_N(_18253_),
    .X(_18261_));
 sky130_fd_sc_hd__o311ai_2 _20956_ (.A1(_18012_),
    .A2(_18253_),
    .A3(_18254_),
    .B1(_18260_),
    .C1(_18261_),
    .Y(_04058_));
 sky130_fd_sc_hd__inv_2 _20957_ (.A(instr_jalr),
    .Y(_02063_));
 sky130_fd_sc_hd__buf_1 _20958_ (.A(instr_jal),
    .X(_18262_));
 sky130_fd_sc_hd__buf_1 _20959_ (.A(_18262_),
    .X(_18263_));
 sky130_fd_sc_hd__a211o_2 _20960_ (.A1(_18033_),
    .A2(_02063_),
    .B1(_18263_),
    .C1(_18079_),
    .X(_18264_));
 sky130_fd_sc_hd__nor2_2 _20961_ (.A(_18263_),
    .B(_18152_),
    .Y(_18265_));
 sky130_fd_sc_hd__inv_2 _20962_ (.A(_18254_),
    .Y(_18266_));
 sky130_fd_sc_hd__o221a_2 _20963_ (.A1(_18151_),
    .A2(_18264_),
    .B1(_18015_),
    .B2(_18265_),
    .C1(_18266_),
    .X(_04057_));
 sky130_fd_sc_hd__nor2_2 _20964_ (.A(_00358_),
    .B(_00357_),
    .Y(_18267_));
 sky130_fd_sc_hd__nor2_2 _20965_ (.A(_00362_),
    .B(_00360_),
    .Y(_18268_));
 sky130_fd_sc_hd__and3_2 _20966_ (.A(_18267_),
    .B(_18268_),
    .C(_00368_),
    .X(_18269_));
 sky130_fd_sc_hd__buf_1 _20967_ (.A(_18269_),
    .X(_18270_));
 sky130_fd_sc_hd__buf_1 _20968_ (.A(_18270_),
    .X(_18271_));
 sky130_fd_sc_hd__nor2_2 _20969_ (.A(_01207_),
    .B(_18271_),
    .Y(\cpuregs_rs1[31] ));
 sky130_fd_sc_hd__nor2_2 _20970_ (.A(_18199_),
    .B(_18193_),
    .Y(_18272_));
 sky130_fd_sc_hd__buf_1 _20971_ (.A(_18272_),
    .X(_18273_));
 sky130_fd_sc_hd__buf_1 _20972_ (.A(_18273_),
    .X(_18274_));
 sky130_fd_sc_hd__buf_1 _20973_ (.A(_18272_),
    .X(_18275_));
 sky130_fd_sc_hd__buf_1 _20974_ (.A(_18275_),
    .X(_18276_));
 sky130_fd_sc_hd__nor2_2 _20975_ (.A(_18129_),
    .B(_18276_),
    .Y(_18277_));
 sky130_fd_sc_hd__a211o_2 _20976_ (.A1(\cpuregs_rs1[31] ),
    .A2(_18274_),
    .B1(_18190_),
    .C1(_18277_),
    .X(_04056_));
 sky130_fd_sc_hd__nor2_2 _20977_ (.A(_01180_),
    .B(_18271_),
    .Y(\cpuregs_rs1[30] ));
 sky130_fd_sc_hd__buf_1 _20978_ (.A(_18051_),
    .X(_18278_));
 sky130_fd_sc_hd__buf_1 _20979_ (.A(_18278_),
    .X(_18279_));
 sky130_fd_sc_hd__nor2_2 _20980_ (.A(_18131_),
    .B(_18276_),
    .Y(_18280_));
 sky130_fd_sc_hd__a211o_2 _20981_ (.A1(\cpuregs_rs1[30] ),
    .A2(_18274_),
    .B1(_18279_),
    .C1(_18280_),
    .X(_04055_));
 sky130_fd_sc_hd__buf_1 _20982_ (.A(_18270_),
    .X(_18281_));
 sky130_fd_sc_hd__nor2_2 _20983_ (.A(_01153_),
    .B(_18281_),
    .Y(\cpuregs_rs1[29] ));
 sky130_fd_sc_hd__nor2_2 _20984_ (.A(_18126_),
    .B(_18276_),
    .Y(_18282_));
 sky130_fd_sc_hd__a211o_2 _20985_ (.A1(\cpuregs_rs1[29] ),
    .A2(_18274_),
    .B1(_18279_),
    .C1(_18282_),
    .X(_04054_));
 sky130_fd_sc_hd__nor2_2 _20986_ (.A(_01126_),
    .B(_18271_),
    .Y(\cpuregs_rs1[28] ));
 sky130_fd_sc_hd__nor2_2 _20987_ (.A(_18127_),
    .B(_18276_),
    .Y(_18283_));
 sky130_fd_sc_hd__a211o_2 _20988_ (.A1(\cpuregs_rs1[28] ),
    .A2(_18274_),
    .B1(_18279_),
    .C1(_18283_),
    .X(_04053_));
 sky130_fd_sc_hd__nor2_2 _20989_ (.A(_01099_),
    .B(_18281_),
    .Y(\cpuregs_rs1[27] ));
 sky130_fd_sc_hd__and2b_2 _20990_ (.A_N(_18273_),
    .B(\irq_mask[27] ),
    .X(_18284_));
 sky130_fd_sc_hd__a211o_2 _20991_ (.A1(\cpuregs_rs1[27] ),
    .A2(_18274_),
    .B1(_18279_),
    .C1(_18284_),
    .X(_04052_));
 sky130_fd_sc_hd__nor2_2 _20992_ (.A(_01072_),
    .B(_18281_),
    .Y(\cpuregs_rs1[26] ));
 sky130_fd_sc_hd__and2b_2 _20993_ (.A_N(_18273_),
    .B(\irq_mask[26] ),
    .X(_18285_));
 sky130_fd_sc_hd__a211o_2 _20994_ (.A1(\cpuregs_rs1[26] ),
    .A2(_18274_),
    .B1(_18279_),
    .C1(_18285_),
    .X(_04051_));
 sky130_fd_sc_hd__nor2_2 _20995_ (.A(_01045_),
    .B(_18281_),
    .Y(\cpuregs_rs1[25] ));
 sky130_fd_sc_hd__buf_1 _20996_ (.A(_18273_),
    .X(_18286_));
 sky130_fd_sc_hd__buf_1 _20997_ (.A(_18275_),
    .X(_18287_));
 sky130_fd_sc_hd__nor2_2 _20998_ (.A(_18099_),
    .B(_18287_),
    .Y(_18288_));
 sky130_fd_sc_hd__a211o_2 _20999_ (.A1(\cpuregs_rs1[25] ),
    .A2(_18286_),
    .B1(_18279_),
    .C1(_18288_),
    .X(_04050_));
 sky130_fd_sc_hd__nor2_2 _21000_ (.A(_01018_),
    .B(_18271_),
    .Y(\cpuregs_rs1[24] ));
 sky130_fd_sc_hd__buf_1 _21001_ (.A(_18278_),
    .X(_18289_));
 sky130_fd_sc_hd__nor2_2 _21002_ (.A(_18100_),
    .B(_18287_),
    .Y(_18290_));
 sky130_fd_sc_hd__a211o_2 _21003_ (.A1(\cpuregs_rs1[24] ),
    .A2(_18286_),
    .B1(_18289_),
    .C1(_18290_),
    .X(_04049_));
 sky130_fd_sc_hd__nor2_2 _21004_ (.A(_00991_),
    .B(_18281_),
    .Y(\cpuregs_rs1[23] ));
 sky130_fd_sc_hd__nor2_2 _21005_ (.A(_18103_),
    .B(_18287_),
    .Y(_18291_));
 sky130_fd_sc_hd__a211o_2 _21006_ (.A1(\cpuregs_rs1[23] ),
    .A2(_18286_),
    .B1(_18289_),
    .C1(_18291_),
    .X(_04048_));
 sky130_fd_sc_hd__nor2_2 _21007_ (.A(_00964_),
    .B(_18281_),
    .Y(\cpuregs_rs1[22] ));
 sky130_fd_sc_hd__nor2_2 _21008_ (.A(_18105_),
    .B(_18287_),
    .Y(_18292_));
 sky130_fd_sc_hd__a211o_2 _21009_ (.A1(\cpuregs_rs1[22] ),
    .A2(_18286_),
    .B1(_18289_),
    .C1(_18292_),
    .X(_04047_));
 sky130_fd_sc_hd__buf_1 _21010_ (.A(_18270_),
    .X(_18293_));
 sky130_fd_sc_hd__nor2_2 _21011_ (.A(_00937_),
    .B(_18293_),
    .Y(\cpuregs_rs1[21] ));
 sky130_fd_sc_hd__nor2_2 _21012_ (.A(_18107_),
    .B(_18287_),
    .Y(_18294_));
 sky130_fd_sc_hd__a211o_2 _21013_ (.A1(\cpuregs_rs1[21] ),
    .A2(_18286_),
    .B1(_18289_),
    .C1(_18294_),
    .X(_04046_));
 sky130_fd_sc_hd__nor2_2 _21014_ (.A(_00910_),
    .B(_18293_),
    .Y(\cpuregs_rs1[20] ));
 sky130_fd_sc_hd__nor2_2 _21015_ (.A(_18108_),
    .B(_18287_),
    .Y(_18295_));
 sky130_fd_sc_hd__a211o_2 _21016_ (.A1(\cpuregs_rs1[20] ),
    .A2(_18286_),
    .B1(_18289_),
    .C1(_18295_),
    .X(_04045_));
 sky130_fd_sc_hd__nor2_2 _21017_ (.A(_00883_),
    .B(_18271_),
    .Y(\cpuregs_rs1[19] ));
 sky130_fd_sc_hd__buf_1 _21018_ (.A(_18275_),
    .X(_18296_));
 sky130_fd_sc_hd__buf_1 _21019_ (.A(_18275_),
    .X(_18297_));
 sky130_fd_sc_hd__nor2_2 _21020_ (.A(_18092_),
    .B(_18297_),
    .Y(_18298_));
 sky130_fd_sc_hd__a211o_2 _21021_ (.A1(\cpuregs_rs1[19] ),
    .A2(_18296_),
    .B1(_18289_),
    .C1(_18298_),
    .X(_04044_));
 sky130_fd_sc_hd__buf_1 _21022_ (.A(_18270_),
    .X(_18299_));
 sky130_fd_sc_hd__nor2_2 _21023_ (.A(_00856_),
    .B(_18299_),
    .Y(\cpuregs_rs1[18] ));
 sky130_fd_sc_hd__buf_1 _21024_ (.A(_18048_),
    .X(_18300_));
 sky130_fd_sc_hd__buf_1 _21025_ (.A(_18300_),
    .X(_18301_));
 sky130_fd_sc_hd__nor2_2 _21026_ (.A(_18094_),
    .B(_18297_),
    .Y(_18302_));
 sky130_fd_sc_hd__a211o_2 _21027_ (.A1(\cpuregs_rs1[18] ),
    .A2(_18296_),
    .B1(_18301_),
    .C1(_18302_),
    .X(_04043_));
 sky130_fd_sc_hd__nor2_2 _21028_ (.A(_00829_),
    .B(_18293_),
    .Y(\cpuregs_rs1[17] ));
 sky130_fd_sc_hd__nor2_2 _21029_ (.A(_18089_),
    .B(_18297_),
    .Y(_18303_));
 sky130_fd_sc_hd__a211o_2 _21030_ (.A1(\cpuregs_rs1[17] ),
    .A2(_18296_),
    .B1(_18301_),
    .C1(_18303_),
    .X(_04042_));
 sky130_fd_sc_hd__nor2_2 _21031_ (.A(_00802_),
    .B(_18299_),
    .Y(\cpuregs_rs1[16] ));
 sky130_fd_sc_hd__inv_2 _21032_ (.A(\irq_mask[16] ),
    .Y(_18304_));
 sky130_fd_sc_hd__nor2_2 _21033_ (.A(_18304_),
    .B(_18297_),
    .Y(_18305_));
 sky130_fd_sc_hd__a211o_2 _21034_ (.A1(\cpuregs_rs1[16] ),
    .A2(_18296_),
    .B1(_18301_),
    .C1(_18305_),
    .X(_04041_));
 sky130_fd_sc_hd__nor2_2 _21035_ (.A(_00775_),
    .B(_18293_),
    .Y(\cpuregs_rs1[15] ));
 sky130_fd_sc_hd__nor2_2 _21036_ (.A(_18137_),
    .B(_18297_),
    .Y(_18306_));
 sky130_fd_sc_hd__a211o_2 _21037_ (.A1(\cpuregs_rs1[15] ),
    .A2(_18296_),
    .B1(_18301_),
    .C1(_18306_),
    .X(_04040_));
 sky130_fd_sc_hd__nor2_2 _21038_ (.A(_00748_),
    .B(_18299_),
    .Y(\cpuregs_rs1[14] ));
 sky130_fd_sc_hd__nor2_2 _21039_ (.A(_18139_),
    .B(_18297_),
    .Y(_18307_));
 sky130_fd_sc_hd__a211o_2 _21040_ (.A1(\cpuregs_rs1[14] ),
    .A2(_18296_),
    .B1(_18301_),
    .C1(_18307_),
    .X(_04039_));
 sky130_fd_sc_hd__nor2_2 _21041_ (.A(_00721_),
    .B(_18293_),
    .Y(\cpuregs_rs1[13] ));
 sky130_fd_sc_hd__buf_1 _21042_ (.A(_18275_),
    .X(_18308_));
 sky130_fd_sc_hd__buf_1 _21043_ (.A(_18272_),
    .X(_18309_));
 sky130_fd_sc_hd__nor2_2 _21044_ (.A(_18134_),
    .B(_18309_),
    .Y(_18310_));
 sky130_fd_sc_hd__a211o_2 _21045_ (.A1(\cpuregs_rs1[13] ),
    .A2(_18308_),
    .B1(_18301_),
    .C1(_18310_),
    .X(_04038_));
 sky130_fd_sc_hd__nor2_2 _21046_ (.A(_00694_),
    .B(_18293_),
    .Y(\cpuregs_rs1[12] ));
 sky130_fd_sc_hd__buf_1 _21047_ (.A(_18300_),
    .X(_18311_));
 sky130_fd_sc_hd__nor2_2 _21048_ (.A(_18135_),
    .B(_18309_),
    .Y(_18312_));
 sky130_fd_sc_hd__a211o_2 _21049_ (.A1(\cpuregs_rs1[12] ),
    .A2(_18308_),
    .B1(_18311_),
    .C1(_18312_),
    .X(_04037_));
 sky130_fd_sc_hd__buf_1 _21050_ (.A(_18270_),
    .X(_18313_));
 sky130_fd_sc_hd__nor2_2 _21051_ (.A(_00667_),
    .B(_18313_),
    .Y(\cpuregs_rs1[11] ));
 sky130_fd_sc_hd__and2b_2 _21052_ (.A_N(_18273_),
    .B(\irq_mask[11] ),
    .X(_18314_));
 sky130_fd_sc_hd__a211o_2 _21053_ (.A1(\cpuregs_rs1[11] ),
    .A2(_18308_),
    .B1(_18311_),
    .C1(_18314_),
    .X(_04036_));
 sky130_fd_sc_hd__nor2_2 _21054_ (.A(_00640_),
    .B(_18313_),
    .Y(\cpuregs_rs1[10] ));
 sky130_fd_sc_hd__and2b_2 _21055_ (.A_N(_18273_),
    .B(\irq_mask[10] ),
    .X(_18315_));
 sky130_fd_sc_hd__a211o_2 _21056_ (.A1(\cpuregs_rs1[10] ),
    .A2(_18308_),
    .B1(_18311_),
    .C1(_18315_),
    .X(_04035_));
 sky130_fd_sc_hd__nor2_2 _21057_ (.A(_00613_),
    .B(_18313_),
    .Y(\cpuregs_rs1[9] ));
 sky130_fd_sc_hd__nor2_2 _21058_ (.A(_18114_),
    .B(_18309_),
    .Y(_18316_));
 sky130_fd_sc_hd__a211o_2 _21059_ (.A1(\cpuregs_rs1[9] ),
    .A2(_18308_),
    .B1(_18311_),
    .C1(_18316_),
    .X(_04034_));
 sky130_fd_sc_hd__nor2_2 _21060_ (.A(_00586_),
    .B(_18299_),
    .Y(\cpuregs_rs1[8] ));
 sky130_fd_sc_hd__nor2_2 _21061_ (.A(_18115_),
    .B(_18309_),
    .Y(_18317_));
 sky130_fd_sc_hd__a211o_2 _21062_ (.A1(\cpuregs_rs1[8] ),
    .A2(_18308_),
    .B1(_18311_),
    .C1(_18317_),
    .X(_04033_));
 sky130_fd_sc_hd__nor2_2 _21063_ (.A(_00559_),
    .B(_18299_),
    .Y(\cpuregs_rs1[7] ));
 sky130_fd_sc_hd__buf_1 _21064_ (.A(_18275_),
    .X(_18318_));
 sky130_fd_sc_hd__nor2_2 _21065_ (.A(_18118_),
    .B(_18309_),
    .Y(_18319_));
 sky130_fd_sc_hd__a211o_2 _21066_ (.A1(\cpuregs_rs1[7] ),
    .A2(_18318_),
    .B1(_18311_),
    .C1(_18319_),
    .X(_04032_));
 sky130_fd_sc_hd__nor2_2 _21067_ (.A(_00532_),
    .B(_18313_),
    .Y(\cpuregs_rs1[6] ));
 sky130_fd_sc_hd__buf_1 _21068_ (.A(_18300_),
    .X(_18320_));
 sky130_fd_sc_hd__nor2_2 _21069_ (.A(_18120_),
    .B(_18309_),
    .Y(_18321_));
 sky130_fd_sc_hd__a211o_2 _21070_ (.A1(\cpuregs_rs1[6] ),
    .A2(_18318_),
    .B1(_18320_),
    .C1(_18321_),
    .X(_04031_));
 sky130_fd_sc_hd__nor2_2 _21071_ (.A(_00505_),
    .B(_18313_),
    .Y(\cpuregs_rs1[5] ));
 sky130_fd_sc_hd__buf_1 _21072_ (.A(_18272_),
    .X(_18322_));
 sky130_fd_sc_hd__nor2_2 _21073_ (.A(_18122_),
    .B(_18322_),
    .Y(_18323_));
 sky130_fd_sc_hd__a211o_2 _21074_ (.A1(\cpuregs_rs1[5] ),
    .A2(_18318_),
    .B1(_18320_),
    .C1(_18323_),
    .X(_04030_));
 sky130_fd_sc_hd__nor2_2 _21075_ (.A(_00478_),
    .B(_18313_),
    .Y(\cpuregs_rs1[4] ));
 sky130_fd_sc_hd__nor2_2 _21076_ (.A(_18123_),
    .B(_18322_),
    .Y(_18324_));
 sky130_fd_sc_hd__a211o_2 _21077_ (.A1(\cpuregs_rs1[4] ),
    .A2(_18318_),
    .B1(_18320_),
    .C1(_18324_),
    .X(_04029_));
 sky130_fd_sc_hd__nor2_2 _21078_ (.A(_00451_),
    .B(_18299_),
    .Y(\cpuregs_rs1[3] ));
 sky130_fd_sc_hd__nor2_2 _21079_ (.A(_18086_),
    .B(_18322_),
    .Y(_18325_));
 sky130_fd_sc_hd__a211o_2 _21080_ (.A1(\cpuregs_rs1[3] ),
    .A2(_18318_),
    .B1(_18320_),
    .C1(_18325_),
    .X(_04028_));
 sky130_fd_sc_hd__nor2_2 _21081_ (.A(_00424_),
    .B(_18271_),
    .Y(\cpuregs_rs1[2] ));
 sky130_fd_sc_hd__nor2_2 _21082_ (.A(_18081_),
    .B(_18322_),
    .Y(_18326_));
 sky130_fd_sc_hd__a211o_2 _21083_ (.A1(\cpuregs_rs1[2] ),
    .A2(_18318_),
    .B1(_18320_),
    .C1(_18326_),
    .X(_04027_));
 sky130_fd_sc_hd__nor2_2 _21084_ (.A(_00397_),
    .B(_18270_),
    .Y(\cpuregs_rs1[1] ));
 sky130_fd_sc_hd__inv_2 _21085_ (.A(\irq_mask[1] ),
    .Y(_18327_));
 sky130_fd_sc_hd__nor2_2 _21086_ (.A(_18327_),
    .B(_18322_),
    .Y(_18328_));
 sky130_fd_sc_hd__a211o_2 _21087_ (.A1(\cpuregs_rs1[1] ),
    .A2(_18276_),
    .B1(_18320_),
    .C1(_18328_),
    .X(_04026_));
 sky130_fd_sc_hd__inv_2 _21088_ (.A(_18269_),
    .Y(_18329_));
 sky130_fd_sc_hd__nand2_2 _21089_ (.A(_18329_),
    .B(_00370_),
    .Y(_18330_));
 sky130_fd_sc_hd__inv_2 _21090_ (.A(_18330_),
    .Y(\cpuregs_rs1[0] ));
 sky130_fd_sc_hd__buf_1 _21091_ (.A(_18300_),
    .X(_18331_));
 sky130_fd_sc_hd__inv_2 _21092_ (.A(\irq_mask[0] ),
    .Y(_18332_));
 sky130_fd_sc_hd__nor2_2 _21093_ (.A(_18332_),
    .B(_18322_),
    .Y(_18333_));
 sky130_fd_sc_hd__a211o_2 _21094_ (.A1(\cpuregs_rs1[0] ),
    .A2(_18276_),
    .B1(_18331_),
    .C1(_18333_),
    .X(_04025_));
 sky130_fd_sc_hd__buf_1 _21095_ (.A(_18043_),
    .X(_00301_));
 sky130_fd_sc_hd__nor2_2 _21096_ (.A(mem_do_wdata),
    .B(_00301_),
    .Y(_18334_));
 sky130_fd_sc_hd__and2_2 _21097_ (.A(_18044_),
    .B(_00290_),
    .X(_18335_));
 sky130_fd_sc_hd__nand2_2 _21098_ (.A(_18335_),
    .B(_18024_),
    .Y(_00316_));
 sky130_fd_sc_hd__nor2_2 _21099_ (.A(trap),
    .B(_00316_),
    .Y(_18336_));
 sky130_fd_sc_hd__buf_1 _21100_ (.A(_18336_),
    .X(_18337_));
 sky130_fd_sc_hd__mux2_2 _21101_ (.A0(mem_instr),
    .A1(_18334_),
    .S(_18337_),
    .X(_04024_));
 sky130_fd_sc_hd__buf_1 _21102_ (.A(is_beq_bne_blt_bge_bltu_bgeu),
    .X(_18338_));
 sky130_fd_sc_hd__buf_1 _21103_ (.A(_18026_),
    .X(_18339_));
 sky130_fd_sc_hd__buf_1 _21104_ (.A(_18339_),
    .X(_18340_));
 sky130_fd_sc_hd__inv_2 _21105_ (.A(_00328_),
    .Y(_18341_));
 sky130_fd_sc_hd__and3_2 _21106_ (.A(_18341_),
    .B(_00329_),
    .C(_00330_),
    .X(_18342_));
 sky130_fd_sc_hd__inv_2 _21107_ (.A(_18060_),
    .Y(_18343_));
 sky130_fd_sc_hd__a31o_2 _21108_ (.A1(_18064_),
    .A2(_18062_),
    .A3(_18342_),
    .B1(_18343_),
    .X(_18344_));
 sky130_fd_sc_hd__o211a_2 _21109_ (.A1(_18338_),
    .A2(_18061_),
    .B1(_18340_),
    .C1(_18344_),
    .X(_04023_));
 sky130_fd_sc_hd__nand2_2 _21110_ (.A(_18061_),
    .B(\mem_rdata_latched[18] ),
    .Y(_18345_));
 sky130_fd_sc_hd__buf_1 _21111_ (.A(_18343_),
    .X(_00337_));
 sky130_fd_sc_hd__a2bb2o_2 _21112_ (.A1_N(_18073_),
    .A2_N(_18345_),
    .B1(\decoded_rs1[3] ),
    .B2(_00337_),
    .X(_04022_));
 sky130_fd_sc_hd__nand2_2 _21113_ (.A(_18077_),
    .B(\mem_rdata_latched[17] ),
    .Y(_18346_));
 sky130_fd_sc_hd__a2bb2o_2 _21114_ (.A1_N(_18073_),
    .A2_N(_18346_),
    .B1(\decoded_rs1[2] ),
    .B2(_00337_),
    .X(_04021_));
 sky130_fd_sc_hd__nand2_2 _21115_ (.A(_18077_),
    .B(\mem_rdata_latched[16] ),
    .Y(_18347_));
 sky130_fd_sc_hd__a2bb2o_2 _21116_ (.A1_N(_18073_),
    .A2_N(_18347_),
    .B1(\decoded_rs1[1] ),
    .B2(_00337_),
    .X(_04020_));
 sky130_fd_sc_hd__nand2_2 _21117_ (.A(_18077_),
    .B(\mem_rdata_latched[15] ),
    .Y(_18348_));
 sky130_fd_sc_hd__a2bb2o_2 _21118_ (.A1_N(_18073_),
    .A2_N(_18348_),
    .B1(\decoded_rs1[0] ),
    .B2(_00337_),
    .X(_04019_));
 sky130_fd_sc_hd__buf_1 _21119_ (.A(_18300_),
    .X(_18349_));
 sky130_fd_sc_hd__buf_1 _21120_ (.A(_18349_),
    .X(_18350_));
 sky130_fd_sc_hd__nor2_2 _21121_ (.A(decoder_pseudo_trigger),
    .B(_18080_),
    .Y(_18351_));
 sky130_fd_sc_hd__buf_1 _21122_ (.A(_18351_),
    .X(_18352_));
 sky130_fd_sc_hd__buf_1 _21123_ (.A(_18352_),
    .X(_18353_));
 sky130_fd_sc_hd__inv_2 _21124_ (.A(\mem_rdata_q[14] ),
    .Y(_00334_));
 sky130_fd_sc_hd__inv_2 _21125_ (.A(\mem_rdata_q[13] ),
    .Y(_18354_));
 sky130_fd_sc_hd__buf_1 _21126_ (.A(_18354_),
    .X(_18355_));
 sky130_fd_sc_hd__inv_2 _21127_ (.A(\mem_rdata_q[12] ),
    .Y(_18356_));
 sky130_fd_sc_hd__or3_2 _21128_ (.A(_00334_),
    .B(_18355_),
    .C(_18356_),
    .X(_18357_));
 sky130_fd_sc_hd__inv_2 _21129_ (.A(is_alu_reg_reg),
    .Y(_18358_));
 sky130_fd_sc_hd__nor2_2 _21130_ (.A(\mem_rdata_q[28] ),
    .B(\mem_rdata_q[26] ),
    .Y(_18359_));
 sky130_fd_sc_hd__inv_2 _21131_ (.A(\mem_rdata_q[27] ),
    .Y(_18360_));
 sky130_fd_sc_hd__inv_2 _21132_ (.A(\mem_rdata_q[25] ),
    .Y(_18361_));
 sky130_fd_sc_hd__and3_2 _21133_ (.A(_18359_),
    .B(_18360_),
    .C(_18361_),
    .X(_18362_));
 sky130_fd_sc_hd__inv_2 _21134_ (.A(\mem_rdata_q[31] ),
    .Y(_18363_));
 sky130_fd_sc_hd__inv_2 _21135_ (.A(\mem_rdata_q[30] ),
    .Y(_18364_));
 sky130_fd_sc_hd__inv_2 _21136_ (.A(\mem_rdata_q[29] ),
    .Y(_18365_));
 sky130_fd_sc_hd__and3_2 _21137_ (.A(_18363_),
    .B(_18364_),
    .C(_18365_),
    .X(_18366_));
 sky130_fd_sc_hd__and3_2 _21138_ (.A(_18362_),
    .B(_18366_),
    .C(_18351_),
    .X(_18367_));
 sky130_fd_sc_hd__inv_2 _21139_ (.A(_18367_),
    .Y(_18368_));
 sky130_fd_sc_hd__nor2_2 _21140_ (.A(_18358_),
    .B(_18368_),
    .Y(_18369_));
 sky130_fd_sc_hd__inv_2 _21141_ (.A(_18369_),
    .Y(_18370_));
 sky130_fd_sc_hd__o22a_2 _21142_ (.A1(_18212_),
    .A2(_18353_),
    .B1(_18357_),
    .B2(_18370_),
    .X(_18371_));
 sky130_fd_sc_hd__nor2_2 _21143_ (.A(_18350_),
    .B(_18371_),
    .Y(_04018_));
 sky130_fd_sc_hd__or3_2 _21144_ (.A(\mem_rdata_q[12] ),
    .B(_00334_),
    .C(_18355_),
    .X(_18372_));
 sky130_fd_sc_hd__o22a_2 _21145_ (.A1(_18213_),
    .A2(_18353_),
    .B1(_18372_),
    .B2(_18370_),
    .X(_18373_));
 sky130_fd_sc_hd__nor2_2 _21146_ (.A(_18350_),
    .B(_18373_),
    .Y(_04017_));
 sky130_fd_sc_hd__and3_2 _21147_ (.A(_18362_),
    .B(_18363_),
    .C(\mem_rdata_q[30] ),
    .X(_18374_));
 sky130_fd_sc_hd__inv_2 _21148_ (.A(decoder_pseudo_trigger),
    .Y(_18375_));
 sky130_fd_sc_hd__and3_2 _21149_ (.A(_18365_),
    .B(_18375_),
    .C(decoder_trigger),
    .X(_18376_));
 sky130_fd_sc_hd__nand2_2 _21150_ (.A(_18374_),
    .B(_18376_),
    .Y(_18377_));
 sky130_fd_sc_hd__inv_2 _21151_ (.A(_18377_),
    .Y(_18378_));
 sky130_fd_sc_hd__buf_1 _21152_ (.A(\mem_rdata_q[14] ),
    .X(_18379_));
 sky130_fd_sc_hd__and3_2 _21153_ (.A(_18355_),
    .B(_18379_),
    .C(\mem_rdata_q[12] ),
    .X(_18380_));
 sky130_fd_sc_hd__inv_2 _21154_ (.A(_18380_),
    .Y(_18381_));
 sky130_fd_sc_hd__nor2_2 _21155_ (.A(_18358_),
    .B(_18381_),
    .Y(_18382_));
 sky130_fd_sc_hd__nand2_2 _21156_ (.A(_18378_),
    .B(_18382_),
    .Y(_18383_));
 sky130_fd_sc_hd__inv_2 _21157_ (.A(_18351_),
    .Y(_18384_));
 sky130_fd_sc_hd__buf_1 _21158_ (.A(_18384_),
    .X(_18385_));
 sky130_fd_sc_hd__buf_1 _21159_ (.A(_18385_),
    .X(_18386_));
 sky130_fd_sc_hd__nand2_2 _21160_ (.A(_18386_),
    .B(instr_sra),
    .Y(_18387_));
 sky130_fd_sc_hd__a21oi_2 _21161_ (.A1(_18383_),
    .A2(_18387_),
    .B1(_18245_),
    .Y(_04016_));
 sky130_fd_sc_hd__buf_1 _21162_ (.A(_18367_),
    .X(_18388_));
 sky130_fd_sc_hd__nand2_2 _21163_ (.A(_18388_),
    .B(_18382_),
    .Y(_18389_));
 sky130_fd_sc_hd__nand2_2 _21164_ (.A(_18386_),
    .B(instr_srl),
    .Y(_18390_));
 sky130_fd_sc_hd__a21oi_2 _21165_ (.A1(_18389_),
    .A2(_18390_),
    .B1(_18245_),
    .Y(_04015_));
 sky130_fd_sc_hd__buf_1 _21166_ (.A(_18384_),
    .X(_18391_));
 sky130_fd_sc_hd__buf_1 _21167_ (.A(_18391_),
    .X(_18392_));
 sky130_fd_sc_hd__and3_2 _21168_ (.A(_18355_),
    .B(_18356_),
    .C(_18379_),
    .X(_18393_));
 sky130_fd_sc_hd__a22o_2 _21169_ (.A1(instr_xor),
    .A2(_18392_),
    .B1(_18369_),
    .B2(_18393_),
    .X(_18394_));
 sky130_fd_sc_hd__buf_1 _21170_ (.A(_18026_),
    .X(_18395_));
 sky130_fd_sc_hd__buf_1 _21171_ (.A(_18395_),
    .X(_18396_));
 sky130_fd_sc_hd__and2_2 _21172_ (.A(_18394_),
    .B(_18396_),
    .X(_04014_));
 sky130_fd_sc_hd__nor2_2 _21173_ (.A(\mem_rdata_q[14] ),
    .B(_18354_),
    .Y(_18397_));
 sky130_fd_sc_hd__buf_1 _21174_ (.A(\mem_rdata_q[12] ),
    .X(_18398_));
 sky130_fd_sc_hd__nand2_2 _21175_ (.A(_18397_),
    .B(_18398_),
    .Y(_18399_));
 sky130_fd_sc_hd__or2_2 _21176_ (.A(_18399_),
    .B(_18370_),
    .X(_18400_));
 sky130_fd_sc_hd__nand2_2 _21177_ (.A(_18386_),
    .B(instr_sltu),
    .Y(_18401_));
 sky130_fd_sc_hd__a21oi_2 _21178_ (.A1(_18400_),
    .A2(_18401_),
    .B1(_18245_),
    .Y(_04013_));
 sky130_fd_sc_hd__nand2_2 _21179_ (.A(_18397_),
    .B(_18356_),
    .Y(_18402_));
 sky130_fd_sc_hd__inv_2 _21180_ (.A(_18402_),
    .Y(_18403_));
 sky130_fd_sc_hd__a22o_2 _21181_ (.A1(instr_slt),
    .A2(_18392_),
    .B1(_18369_),
    .B2(_18403_),
    .X(_18404_));
 sky130_fd_sc_hd__and2_2 _21182_ (.A(_18404_),
    .B(_18396_),
    .X(_04012_));
 sky130_fd_sc_hd__and3_2 _21183_ (.A(_00334_),
    .B(_18355_),
    .C(_18398_),
    .X(_18405_));
 sky130_fd_sc_hd__a22o_2 _21184_ (.A1(instr_sll),
    .A2(_18392_),
    .B1(_18369_),
    .B2(_18405_),
    .X(_18406_));
 sky130_fd_sc_hd__buf_1 _21185_ (.A(_18339_),
    .X(_18407_));
 sky130_fd_sc_hd__and2_2 _21186_ (.A(_18406_),
    .B(_18407_),
    .X(_04011_));
 sky130_fd_sc_hd__and3_2 _21187_ (.A(_00334_),
    .B(_18354_),
    .C(_18356_),
    .X(_18408_));
 sky130_fd_sc_hd__inv_2 _21188_ (.A(_18408_),
    .Y(_18409_));
 sky130_fd_sc_hd__or3_2 _21189_ (.A(_18358_),
    .B(_18409_),
    .C(_18377_),
    .X(_18410_));
 sky130_fd_sc_hd__nand2_2 _21190_ (.A(_18386_),
    .B(instr_sub),
    .Y(_18411_));
 sky130_fd_sc_hd__a21oi_2 _21191_ (.A1(_18410_),
    .A2(_18411_),
    .B1(_18245_),
    .Y(_04010_));
 sky130_fd_sc_hd__a32o_2 _21192_ (.A1(_18388_),
    .A2(is_alu_reg_reg),
    .A3(_18408_),
    .B1(instr_add),
    .B2(_18392_),
    .X(_18412_));
 sky130_fd_sc_hd__and2_2 _21193_ (.A(_18412_),
    .B(_18407_),
    .X(_04009_));
 sky130_fd_sc_hd__buf_1 _21194_ (.A(_18391_),
    .X(_18413_));
 sky130_fd_sc_hd__nand2_2 _21195_ (.A(_18352_),
    .B(is_alu_reg_imm),
    .Y(_18414_));
 sky130_fd_sc_hd__buf_1 _21196_ (.A(_18414_),
    .X(_18415_));
 sky130_fd_sc_hd__o2bb2a_2 _21197_ (.A1_N(instr_andi),
    .A2_N(_18413_),
    .B1(_18415_),
    .B2(_18357_),
    .X(_18416_));
 sky130_fd_sc_hd__nor2_2 _21198_ (.A(_18350_),
    .B(_18416_),
    .Y(_04008_));
 sky130_fd_sc_hd__o2bb2a_2 _21199_ (.A1_N(instr_ori),
    .A2_N(_18413_),
    .B1(_18415_),
    .B2(_18372_),
    .X(_18417_));
 sky130_fd_sc_hd__nor2_2 _21200_ (.A(_18350_),
    .B(_18417_),
    .Y(_04007_));
 sky130_fd_sc_hd__inv_2 _21201_ (.A(_18393_),
    .Y(_18418_));
 sky130_fd_sc_hd__o2bb2a_2 _21202_ (.A1_N(instr_xori),
    .A2_N(_18413_),
    .B1(_18415_),
    .B2(_18418_),
    .X(_18419_));
 sky130_fd_sc_hd__nor2_2 _21203_ (.A(_18350_),
    .B(_18419_),
    .Y(_04006_));
 sky130_fd_sc_hd__buf_1 _21204_ (.A(_18349_),
    .X(_18420_));
 sky130_fd_sc_hd__o2bb2a_2 _21205_ (.A1_N(instr_sltiu),
    .A2_N(_18413_),
    .B1(_18399_),
    .B2(_18415_),
    .X(_18421_));
 sky130_fd_sc_hd__nor2_2 _21206_ (.A(_18420_),
    .B(_18421_),
    .Y(_04005_));
 sky130_fd_sc_hd__o2bb2a_2 _21207_ (.A1_N(instr_slti),
    .A2_N(_18413_),
    .B1(_18402_),
    .B2(_18414_),
    .X(_18422_));
 sky130_fd_sc_hd__nor2_2 _21208_ (.A(_18420_),
    .B(_18422_),
    .Y(_04004_));
 sky130_fd_sc_hd__o2bb2a_2 _21209_ (.A1_N(instr_addi),
    .A2_N(_18413_),
    .B1(_18415_),
    .B2(_18409_),
    .X(_18423_));
 sky130_fd_sc_hd__nor2_2 _21210_ (.A(_18420_),
    .B(_18423_),
    .Y(_04003_));
 sky130_fd_sc_hd__inv_2 _21211_ (.A(instr_bgeu),
    .Y(_18424_));
 sky130_fd_sc_hd__nand2_2 _21212_ (.A(_18352_),
    .B(_18338_),
    .Y(_18425_));
 sky130_fd_sc_hd__o22a_2 _21213_ (.A1(_18424_),
    .A2(_18353_),
    .B1(_18425_),
    .B2(_18357_),
    .X(_18426_));
 sky130_fd_sc_hd__nor2_2 _21214_ (.A(_18420_),
    .B(_18426_),
    .Y(_04002_));
 sky130_fd_sc_hd__buf_1 _21215_ (.A(_18391_),
    .X(_18427_));
 sky130_fd_sc_hd__o2bb2a_2 _21216_ (.A1_N(instr_bltu),
    .A2_N(_18427_),
    .B1(_18425_),
    .B2(_18372_),
    .X(_18428_));
 sky130_fd_sc_hd__nor2_2 _21217_ (.A(_18420_),
    .B(_18428_),
    .Y(_04001_));
 sky130_fd_sc_hd__o2bb2a_2 _21218_ (.A1_N(instr_bge),
    .A2_N(_18427_),
    .B1(_18425_),
    .B2(_18381_),
    .X(_18429_));
 sky130_fd_sc_hd__nor2_2 _21219_ (.A(_18420_),
    .B(_18429_),
    .Y(_04000_));
 sky130_fd_sc_hd__o2bb2a_2 _21220_ (.A1_N(instr_blt),
    .A2_N(_18427_),
    .B1(_18425_),
    .B2(_18418_),
    .X(_18430_));
 sky130_fd_sc_hd__nor2_2 _21221_ (.A(_18239_),
    .B(_18430_),
    .Y(_03999_));
 sky130_fd_sc_hd__nand2_2 _21222_ (.A(_00334_),
    .B(_18355_),
    .Y(_18431_));
 sky130_fd_sc_hd__inv_2 _21223_ (.A(instr_bne),
    .Y(_18432_));
 sky130_fd_sc_hd__o32a_2 _21224_ (.A1(_18356_),
    .A2(_18431_),
    .A3(_18425_),
    .B1(_18432_),
    .B2(_18353_),
    .X(_18433_));
 sky130_fd_sc_hd__nor2_2 _21225_ (.A(_18239_),
    .B(_18433_),
    .Y(_03998_));
 sky130_fd_sc_hd__o2bb2a_2 _21226_ (.A1_N(instr_beq),
    .A2_N(_18427_),
    .B1(_18425_),
    .B2(_18409_),
    .X(_18434_));
 sky130_fd_sc_hd__nor2_2 _21227_ (.A(_18239_),
    .B(_18434_),
    .Y(_03997_));
 sky130_fd_sc_hd__nor2_2 _21228_ (.A(\pcpi_timeout_counter[1] ),
    .B(\pcpi_timeout_counter[0] ),
    .Y(_18435_));
 sky130_fd_sc_hd__inv_2 _21229_ (.A(\pcpi_timeout_counter[2] ),
    .Y(_18436_));
 sky130_fd_sc_hd__nand2_2 _21230_ (.A(_18435_),
    .B(_18436_),
    .Y(_18437_));
 sky130_fd_sc_hd__a21o_2 _21231_ (.A1(_18437_),
    .A2(\pcpi_timeout_counter[3] ),
    .B1(_18159_),
    .X(_03996_));
 sky130_fd_sc_hd__nor2_2 _21232_ (.A(_18436_),
    .B(_18435_),
    .Y(_18438_));
 sky130_fd_sc_hd__inv_2 _21233_ (.A(\pcpi_timeout_counter[3] ),
    .Y(_18439_));
 sky130_fd_sc_hd__nor2_2 _21234_ (.A(_18439_),
    .B(_18437_),
    .Y(_18440_));
 sky130_fd_sc_hd__or3_2 _21235_ (.A(_18159_),
    .B(_18438_),
    .C(_18440_),
    .X(_03995_));
 sky130_fd_sc_hd__o21a_2 _21236_ (.A1(\pcpi_timeout_counter[3] ),
    .A2(\pcpi_timeout_counter[2] ),
    .B1(_18435_),
    .X(_18441_));
 sky130_fd_sc_hd__a211o_2 _21237_ (.A1(\pcpi_timeout_counter[1] ),
    .A2(\pcpi_timeout_counter[0] ),
    .B1(_18159_),
    .C1(_18441_),
    .X(_03994_));
 sky130_fd_sc_hd__and3_2 _21238_ (.A(_18435_),
    .B(_18439_),
    .C(_18436_),
    .X(_18442_));
 sky130_fd_sc_hd__o21bai_2 _21239_ (.A1(\pcpi_timeout_counter[0] ),
    .A2(_18442_),
    .B1_N(_18159_),
    .Y(_03993_));
 sky130_fd_sc_hd__nor2_2 _21240_ (.A(_18250_),
    .B(_18257_),
    .Y(_18443_));
 sky130_fd_sc_hd__buf_1 _21241_ (.A(_18205_),
    .X(_18444_));
 sky130_fd_sc_hd__and3_2 _21242_ (.A(_18443_),
    .B(_18186_),
    .C(_18444_),
    .X(_01706_));
 sky130_fd_sc_hd__inv_2 _21243_ (.A(mem_do_wdata),
    .Y(_00291_));
 sky130_fd_sc_hd__inv_2 _21244_ (.A(\cpu_state[0] ),
    .Y(_18445_));
 sky130_fd_sc_hd__and3_2 _21245_ (.A(_00291_),
    .B(_18241_),
    .C(_18445_),
    .X(_18446_));
 sky130_fd_sc_hd__a32o_2 _21246_ (.A1(_18018_),
    .A2(_01706_),
    .A3(_18446_),
    .B1(_18266_),
    .B2(mem_do_wdata),
    .X(_03992_));
 sky130_fd_sc_hd__inv_2 _21247_ (.A(_18015_),
    .Y(_18447_));
 sky130_fd_sc_hd__nor2_2 _21248_ (.A(_18447_),
    .B(_18056_),
    .Y(_00296_));
 sky130_fd_sc_hd__inv_2 _21249_ (.A(_00296_),
    .Y(_18448_));
 sky130_fd_sc_hd__and3_2 _21250_ (.A(_18019_),
    .B(_18025_),
    .C(\cpu_state[6] ),
    .X(_18449_));
 sky130_fd_sc_hd__a22o_2 _21251_ (.A1(mem_do_rdata),
    .A2(_18266_),
    .B1(_18448_),
    .B2(_18449_),
    .X(_03991_));
 sky130_fd_sc_hd__buf_1 _21252_ (.A(_18241_),
    .X(_18450_));
 sky130_fd_sc_hd__buf_1 _21253_ (.A(\cpu_state[1] ),
    .X(_18451_));
 sky130_fd_sc_hd__buf_1 _21254_ (.A(_18451_),
    .X(_18452_));
 sky130_fd_sc_hd__or2_2 _21255_ (.A(\reg_next_pc[31] ),
    .B(_18452_),
    .X(_18453_));
 sky130_fd_sc_hd__o211a_2 _21256_ (.A1(_02530_),
    .A2(_18450_),
    .B1(_18340_),
    .C1(_18453_),
    .X(_03990_));
 sky130_fd_sc_hd__buf_1 _21257_ (.A(_18235_),
    .X(_00322_));
 sky130_fd_sc_hd__buf_1 _21258_ (.A(_18451_),
    .X(_18454_));
 sky130_fd_sc_hd__or2_2 _21259_ (.A(_18454_),
    .B(\reg_next_pc[30] ),
    .X(_18455_));
 sky130_fd_sc_hd__o211a_2 _21260_ (.A1(_00322_),
    .A2(_02529_),
    .B1(_18340_),
    .C1(_18455_),
    .X(_03989_));
 sky130_fd_sc_hd__or2_2 _21261_ (.A(_18454_),
    .B(\reg_next_pc[29] ),
    .X(_18456_));
 sky130_fd_sc_hd__o211a_2 _21262_ (.A1(_00322_),
    .A2(_02527_),
    .B1(_18340_),
    .C1(_18456_),
    .X(_03988_));
 sky130_fd_sc_hd__or2_2 _21263_ (.A(_18454_),
    .B(\reg_next_pc[28] ),
    .X(_18457_));
 sky130_fd_sc_hd__o211a_2 _21264_ (.A1(_00322_),
    .A2(_02526_),
    .B1(_18340_),
    .C1(_18457_),
    .X(_03987_));
 sky130_fd_sc_hd__or2_2 _21265_ (.A(_18454_),
    .B(\reg_next_pc[27] ),
    .X(_18458_));
 sky130_fd_sc_hd__o211a_2 _21266_ (.A1(_00322_),
    .A2(_02525_),
    .B1(_18340_),
    .C1(_18458_),
    .X(_03986_));
 sky130_fd_sc_hd__buf_1 _21267_ (.A(_18339_),
    .X(_18459_));
 sky130_fd_sc_hd__or2_2 _21268_ (.A(_18454_),
    .B(\reg_next_pc[26] ),
    .X(_18460_));
 sky130_fd_sc_hd__o211a_2 _21269_ (.A1(_00322_),
    .A2(_02524_),
    .B1(_18459_),
    .C1(_18460_),
    .X(_03985_));
 sky130_fd_sc_hd__buf_1 _21270_ (.A(_18235_),
    .X(_18461_));
 sky130_fd_sc_hd__buf_1 _21271_ (.A(\cpu_state[1] ),
    .X(_18462_));
 sky130_fd_sc_hd__buf_1 _21272_ (.A(_18462_),
    .X(_18463_));
 sky130_fd_sc_hd__or2_2 _21273_ (.A(_18463_),
    .B(\reg_next_pc[25] ),
    .X(_18464_));
 sky130_fd_sc_hd__o211a_2 _21274_ (.A1(_18461_),
    .A2(_02523_),
    .B1(_18459_),
    .C1(_18464_),
    .X(_03984_));
 sky130_fd_sc_hd__or2_2 _21275_ (.A(_18463_),
    .B(\reg_next_pc[24] ),
    .X(_18465_));
 sky130_fd_sc_hd__o211a_2 _21276_ (.A1(_18461_),
    .A2(_02522_),
    .B1(_18459_),
    .C1(_18465_),
    .X(_03983_));
 sky130_fd_sc_hd__or2_2 _21277_ (.A(_18463_),
    .B(\reg_next_pc[23] ),
    .X(_18466_));
 sky130_fd_sc_hd__o211a_2 _21278_ (.A1(_18461_),
    .A2(_02521_),
    .B1(_18459_),
    .C1(_18466_),
    .X(_03982_));
 sky130_fd_sc_hd__or2_2 _21279_ (.A(_18463_),
    .B(\reg_next_pc[22] ),
    .X(_18467_));
 sky130_fd_sc_hd__o211a_2 _21280_ (.A1(_18461_),
    .A2(_02520_),
    .B1(_18459_),
    .C1(_18467_),
    .X(_03981_));
 sky130_fd_sc_hd__or2_2 _21281_ (.A(_18463_),
    .B(\reg_next_pc[21] ),
    .X(_18468_));
 sky130_fd_sc_hd__o211a_2 _21282_ (.A1(_18461_),
    .A2(_02519_),
    .B1(_18459_),
    .C1(_18468_),
    .X(_03980_));
 sky130_fd_sc_hd__buf_1 _21283_ (.A(_18339_),
    .X(_18469_));
 sky130_fd_sc_hd__or2_2 _21284_ (.A(_18463_),
    .B(\reg_next_pc[20] ),
    .X(_18470_));
 sky130_fd_sc_hd__o211a_2 _21285_ (.A1(_18461_),
    .A2(_02518_),
    .B1(_18469_),
    .C1(_18470_),
    .X(_03979_));
 sky130_fd_sc_hd__buf_1 _21286_ (.A(_18235_),
    .X(_18471_));
 sky130_fd_sc_hd__buf_1 _21287_ (.A(_18451_),
    .X(_18472_));
 sky130_fd_sc_hd__or2_2 _21288_ (.A(_18472_),
    .B(\reg_next_pc[19] ),
    .X(_18473_));
 sky130_fd_sc_hd__o211a_2 _21289_ (.A1(_18471_),
    .A2(_02516_),
    .B1(_18469_),
    .C1(_18473_),
    .X(_03978_));
 sky130_fd_sc_hd__or2_2 _21290_ (.A(_18472_),
    .B(\reg_next_pc[18] ),
    .X(_18474_));
 sky130_fd_sc_hd__o211a_2 _21291_ (.A1(_18471_),
    .A2(_02515_),
    .B1(_18469_),
    .C1(_18474_),
    .X(_03977_));
 sky130_fd_sc_hd__or2_2 _21292_ (.A(_18472_),
    .B(\reg_next_pc[17] ),
    .X(_18475_));
 sky130_fd_sc_hd__o211a_2 _21293_ (.A1(_18471_),
    .A2(_02514_),
    .B1(_18469_),
    .C1(_18475_),
    .X(_03976_));
 sky130_fd_sc_hd__or2_2 _21294_ (.A(_18472_),
    .B(\reg_next_pc[16] ),
    .X(_18476_));
 sky130_fd_sc_hd__o211a_2 _21295_ (.A1(_18471_),
    .A2(_02513_),
    .B1(_18469_),
    .C1(_18476_),
    .X(_03975_));
 sky130_fd_sc_hd__or2_2 _21296_ (.A(_18472_),
    .B(\reg_next_pc[15] ),
    .X(_18477_));
 sky130_fd_sc_hd__o211a_2 _21297_ (.A1(_18471_),
    .A2(_02512_),
    .B1(_18469_),
    .C1(_18477_),
    .X(_03974_));
 sky130_fd_sc_hd__buf_1 _21298_ (.A(_18339_),
    .X(_18478_));
 sky130_fd_sc_hd__or2_2 _21299_ (.A(_18472_),
    .B(\reg_next_pc[14] ),
    .X(_18479_));
 sky130_fd_sc_hd__o211a_2 _21300_ (.A1(_18471_),
    .A2(_02511_),
    .B1(_18478_),
    .C1(_18479_),
    .X(_03973_));
 sky130_fd_sc_hd__buf_1 _21301_ (.A(_18235_),
    .X(_18480_));
 sky130_fd_sc_hd__buf_1 _21302_ (.A(_18451_),
    .X(_18481_));
 sky130_fd_sc_hd__or2_2 _21303_ (.A(_18481_),
    .B(\reg_next_pc[13] ),
    .X(_18482_));
 sky130_fd_sc_hd__o211a_2 _21304_ (.A1(_18480_),
    .A2(_02510_),
    .B1(_18478_),
    .C1(_18482_),
    .X(_03972_));
 sky130_fd_sc_hd__or2_2 _21305_ (.A(_18481_),
    .B(\reg_next_pc[12] ),
    .X(_18483_));
 sky130_fd_sc_hd__o211a_2 _21306_ (.A1(_18480_),
    .A2(_02509_),
    .B1(_18478_),
    .C1(_18483_),
    .X(_03971_));
 sky130_fd_sc_hd__or2_2 _21307_ (.A(_18481_),
    .B(\reg_next_pc[11] ),
    .X(_18484_));
 sky130_fd_sc_hd__o211a_2 _21308_ (.A1(_18480_),
    .A2(_02508_),
    .B1(_18478_),
    .C1(_18484_),
    .X(_03970_));
 sky130_fd_sc_hd__or2_2 _21309_ (.A(_18481_),
    .B(\reg_next_pc[10] ),
    .X(_18485_));
 sky130_fd_sc_hd__o211a_2 _21310_ (.A1(_18480_),
    .A2(_02507_),
    .B1(_18478_),
    .C1(_18485_),
    .X(_03969_));
 sky130_fd_sc_hd__or2_2 _21311_ (.A(_18481_),
    .B(\reg_next_pc[9] ),
    .X(_18486_));
 sky130_fd_sc_hd__o211a_2 _21312_ (.A1(_18480_),
    .A2(_02537_),
    .B1(_18478_),
    .C1(_18486_),
    .X(_03968_));
 sky130_fd_sc_hd__buf_1 _21313_ (.A(_18339_),
    .X(_18487_));
 sky130_fd_sc_hd__or2_2 _21314_ (.A(_18481_),
    .B(\reg_next_pc[8] ),
    .X(_18488_));
 sky130_fd_sc_hd__o211a_2 _21315_ (.A1(_18480_),
    .A2(_02536_),
    .B1(_18487_),
    .C1(_18488_),
    .X(_03967_));
 sky130_fd_sc_hd__buf_1 _21316_ (.A(_18241_),
    .X(_18489_));
 sky130_fd_sc_hd__buf_1 _21317_ (.A(_18451_),
    .X(_18490_));
 sky130_fd_sc_hd__or2_2 _21318_ (.A(_18490_),
    .B(\reg_next_pc[7] ),
    .X(_18491_));
 sky130_fd_sc_hd__o211a_2 _21319_ (.A1(_18489_),
    .A2(_02535_),
    .B1(_18487_),
    .C1(_18491_),
    .X(_03966_));
 sky130_fd_sc_hd__or2_2 _21320_ (.A(_18490_),
    .B(\reg_next_pc[6] ),
    .X(_18492_));
 sky130_fd_sc_hd__o211a_2 _21321_ (.A1(_18489_),
    .A2(_02534_),
    .B1(_18487_),
    .C1(_18492_),
    .X(_03965_));
 sky130_fd_sc_hd__or2_2 _21322_ (.A(_18490_),
    .B(\reg_next_pc[5] ),
    .X(_18493_));
 sky130_fd_sc_hd__o211a_2 _21323_ (.A1(_18489_),
    .A2(_02533_),
    .B1(_18487_),
    .C1(_18493_),
    .X(_03964_));
 sky130_fd_sc_hd__buf_1 _21324_ (.A(_18241_),
    .X(_18494_));
 sky130_fd_sc_hd__inv_2 _21325_ (.A(\reg_next_pc[4] ),
    .Y(_01471_));
 sky130_fd_sc_hd__nand2_2 _21326_ (.A(_18494_),
    .B(_01471_),
    .Y(_18495_));
 sky130_fd_sc_hd__o211a_2 _21327_ (.A1(_18489_),
    .A2(_02532_),
    .B1(_18487_),
    .C1(_18495_),
    .X(_03963_));
 sky130_fd_sc_hd__or2_2 _21328_ (.A(_18490_),
    .B(\reg_next_pc[3] ),
    .X(_18496_));
 sky130_fd_sc_hd__o211a_2 _21329_ (.A1(_18489_),
    .A2(_02531_),
    .B1(_18487_),
    .C1(_18496_),
    .X(_03962_));
 sky130_fd_sc_hd__buf_1 _21330_ (.A(_18026_),
    .X(_18497_));
 sky130_fd_sc_hd__buf_1 _21331_ (.A(_18497_),
    .X(_18498_));
 sky130_fd_sc_hd__or2_2 _21332_ (.A(_18490_),
    .B(\reg_next_pc[2] ),
    .X(_18499_));
 sky130_fd_sc_hd__o211a_2 _21333_ (.A1(_18489_),
    .A2(_02528_),
    .B1(_18498_),
    .C1(_18499_),
    .X(_03961_));
 sky130_fd_sc_hd__or2_2 _21334_ (.A(_18490_),
    .B(\reg_next_pc[1] ),
    .X(_18500_));
 sky130_fd_sc_hd__o211a_2 _21335_ (.A1(_18450_),
    .A2(_02517_),
    .B1(_18498_),
    .C1(_18500_),
    .X(_03960_));
 sky130_fd_sc_hd__buf_1 _21336_ (.A(_18452_),
    .X(_18501_));
 sky130_fd_sc_hd__inv_2 _21337_ (.A(_02581_),
    .Y(_18502_));
 sky130_fd_sc_hd__buf_1 _21338_ (.A(_18462_),
    .X(_18503_));
 sky130_fd_sc_hd__nand2_2 _21339_ (.A(_18502_),
    .B(_18503_),
    .Y(_18504_));
 sky130_fd_sc_hd__o211a_2 _21340_ (.A1(_18501_),
    .A2(\reg_pc[31] ),
    .B1(_18498_),
    .C1(_18504_),
    .X(_03959_));
 sky130_fd_sc_hd__inv_2 _21341_ (.A(\reg_pc[30] ),
    .Y(_18505_));
 sky130_fd_sc_hd__nand2_2 _21342_ (.A(_18494_),
    .B(_18505_),
    .Y(_18506_));
 sky130_fd_sc_hd__o211a_2 _21343_ (.A1(_18450_),
    .A2(_02580_),
    .B1(_18498_),
    .C1(_18506_),
    .X(_03958_));
 sky130_fd_sc_hd__inv_2 _21344_ (.A(_02579_),
    .Y(_18507_));
 sky130_fd_sc_hd__buf_1 _21345_ (.A(_18462_),
    .X(_18508_));
 sky130_fd_sc_hd__nand2_2 _21346_ (.A(_18507_),
    .B(_18508_),
    .Y(_18509_));
 sky130_fd_sc_hd__o211a_2 _21347_ (.A1(_18501_),
    .A2(\reg_pc[29] ),
    .B1(_18498_),
    .C1(_18509_),
    .X(_03957_));
 sky130_fd_sc_hd__inv_2 _21348_ (.A(_02578_),
    .Y(_18510_));
 sky130_fd_sc_hd__nand2_2 _21349_ (.A(_18510_),
    .B(_18508_),
    .Y(_18511_));
 sky130_fd_sc_hd__o211a_2 _21350_ (.A1(_18501_),
    .A2(\reg_pc[28] ),
    .B1(_18498_),
    .C1(_18511_),
    .X(_03956_));
 sky130_fd_sc_hd__buf_1 _21351_ (.A(_18497_),
    .X(_18512_));
 sky130_fd_sc_hd__inv_2 _21352_ (.A(_02577_),
    .Y(_18513_));
 sky130_fd_sc_hd__nand2_2 _21353_ (.A(_18513_),
    .B(_18508_),
    .Y(_18514_));
 sky130_fd_sc_hd__o211a_2 _21354_ (.A1(_18501_),
    .A2(\reg_pc[27] ),
    .B1(_18512_),
    .C1(_18514_),
    .X(_03955_));
 sky130_fd_sc_hd__inv_2 _21355_ (.A(_02576_),
    .Y(_18515_));
 sky130_fd_sc_hd__nand2_2 _21356_ (.A(_18515_),
    .B(_18508_),
    .Y(_18516_));
 sky130_fd_sc_hd__o211a_2 _21357_ (.A1(_18501_),
    .A2(\reg_pc[26] ),
    .B1(_18512_),
    .C1(_18516_),
    .X(_03954_));
 sky130_fd_sc_hd__buf_1 _21358_ (.A(_18452_),
    .X(_18517_));
 sky130_fd_sc_hd__inv_2 _21359_ (.A(_02575_),
    .Y(_18518_));
 sky130_fd_sc_hd__nand2_2 _21360_ (.A(_18518_),
    .B(_18508_),
    .Y(_18519_));
 sky130_fd_sc_hd__o211a_2 _21361_ (.A1(_18517_),
    .A2(\reg_pc[25] ),
    .B1(_18512_),
    .C1(_18519_),
    .X(_03953_));
 sky130_fd_sc_hd__inv_2 _21362_ (.A(_02574_),
    .Y(_18520_));
 sky130_fd_sc_hd__nand2_2 _21363_ (.A(_18520_),
    .B(_18508_),
    .Y(_18521_));
 sky130_fd_sc_hd__o211a_2 _21364_ (.A1(_18517_),
    .A2(\reg_pc[24] ),
    .B1(_18512_),
    .C1(_18521_),
    .X(_03952_));
 sky130_fd_sc_hd__inv_2 _21365_ (.A(_02573_),
    .Y(_18522_));
 sky130_fd_sc_hd__buf_1 _21366_ (.A(_18462_),
    .X(_18523_));
 sky130_fd_sc_hd__nand2_2 _21367_ (.A(_18522_),
    .B(_18523_),
    .Y(_18524_));
 sky130_fd_sc_hd__o211a_2 _21368_ (.A1(_18517_),
    .A2(\reg_pc[23] ),
    .B1(_18512_),
    .C1(_18524_),
    .X(_03951_));
 sky130_fd_sc_hd__inv_2 _21369_ (.A(_02572_),
    .Y(_18525_));
 sky130_fd_sc_hd__nand2_2 _21370_ (.A(_18525_),
    .B(_18523_),
    .Y(_18526_));
 sky130_fd_sc_hd__o211a_2 _21371_ (.A1(_18517_),
    .A2(\reg_pc[22] ),
    .B1(_18512_),
    .C1(_18526_),
    .X(_03950_));
 sky130_fd_sc_hd__buf_1 _21372_ (.A(_18497_),
    .X(_18527_));
 sky130_fd_sc_hd__inv_2 _21373_ (.A(_02570_),
    .Y(_18528_));
 sky130_fd_sc_hd__nand2_2 _21374_ (.A(_18528_),
    .B(_18523_),
    .Y(_18529_));
 sky130_fd_sc_hd__o211a_2 _21375_ (.A1(_18517_),
    .A2(\reg_pc[21] ),
    .B1(_18527_),
    .C1(_18529_),
    .X(_03949_));
 sky130_fd_sc_hd__inv_2 _21376_ (.A(_02569_),
    .Y(_18530_));
 sky130_fd_sc_hd__nand2_2 _21377_ (.A(_18530_),
    .B(_18523_),
    .Y(_18531_));
 sky130_fd_sc_hd__o211a_2 _21378_ (.A1(_18517_),
    .A2(\reg_pc[20] ),
    .B1(_18527_),
    .C1(_18531_),
    .X(_03948_));
 sky130_fd_sc_hd__buf_1 _21379_ (.A(_18452_),
    .X(_18532_));
 sky130_fd_sc_hd__inv_2 _21380_ (.A(_02568_),
    .Y(_18533_));
 sky130_fd_sc_hd__nand2_2 _21381_ (.A(_18533_),
    .B(_18523_),
    .Y(_18534_));
 sky130_fd_sc_hd__o211a_2 _21382_ (.A1(_18532_),
    .A2(\reg_pc[19] ),
    .B1(_18527_),
    .C1(_18534_),
    .X(_03947_));
 sky130_fd_sc_hd__inv_2 _21383_ (.A(_02567_),
    .Y(_18535_));
 sky130_fd_sc_hd__nand2_2 _21384_ (.A(_18535_),
    .B(_18523_),
    .Y(_18536_));
 sky130_fd_sc_hd__o211a_2 _21385_ (.A1(_18532_),
    .A2(\reg_pc[18] ),
    .B1(_18527_),
    .C1(_18536_),
    .X(_03946_));
 sky130_fd_sc_hd__inv_2 _21386_ (.A(_02566_),
    .Y(_18537_));
 sky130_fd_sc_hd__buf_1 _21387_ (.A(_18462_),
    .X(_18538_));
 sky130_fd_sc_hd__nand2_2 _21388_ (.A(_18537_),
    .B(_18538_),
    .Y(_18539_));
 sky130_fd_sc_hd__o211a_2 _21389_ (.A1(_18532_),
    .A2(\reg_pc[17] ),
    .B1(_18527_),
    .C1(_18539_),
    .X(_03945_));
 sky130_fd_sc_hd__inv_2 _21390_ (.A(_02565_),
    .Y(_18540_));
 sky130_fd_sc_hd__nand2_2 _21391_ (.A(_18540_),
    .B(_18538_),
    .Y(_18541_));
 sky130_fd_sc_hd__o211a_2 _21392_ (.A1(_18532_),
    .A2(\reg_pc[16] ),
    .B1(_18527_),
    .C1(_18541_),
    .X(_03944_));
 sky130_fd_sc_hd__buf_1 _21393_ (.A(_18497_),
    .X(_18542_));
 sky130_fd_sc_hd__inv_2 _21394_ (.A(_02564_),
    .Y(_18543_));
 sky130_fd_sc_hd__nand2_2 _21395_ (.A(_18543_),
    .B(_18538_),
    .Y(_18544_));
 sky130_fd_sc_hd__o211a_2 _21396_ (.A1(_18532_),
    .A2(\reg_pc[15] ),
    .B1(_18542_),
    .C1(_18544_),
    .X(_03943_));
 sky130_fd_sc_hd__inv_2 _21397_ (.A(_02563_),
    .Y(_18545_));
 sky130_fd_sc_hd__nand2_2 _21398_ (.A(_18545_),
    .B(_18538_),
    .Y(_18546_));
 sky130_fd_sc_hd__o211a_2 _21399_ (.A1(_18532_),
    .A2(\reg_pc[14] ),
    .B1(_18542_),
    .C1(_18546_),
    .X(_03942_));
 sky130_fd_sc_hd__buf_1 _21400_ (.A(_18452_),
    .X(_18547_));
 sky130_fd_sc_hd__inv_2 _21401_ (.A(_02562_),
    .Y(_18548_));
 sky130_fd_sc_hd__nand2_2 _21402_ (.A(_18548_),
    .B(_18538_),
    .Y(_18549_));
 sky130_fd_sc_hd__o211a_2 _21403_ (.A1(_18547_),
    .A2(\reg_pc[13] ),
    .B1(_18542_),
    .C1(_18549_),
    .X(_03941_));
 sky130_fd_sc_hd__inv_2 _21404_ (.A(_02561_),
    .Y(_18550_));
 sky130_fd_sc_hd__nand2_2 _21405_ (.A(_18550_),
    .B(_18538_),
    .Y(_18551_));
 sky130_fd_sc_hd__o211a_2 _21406_ (.A1(_18547_),
    .A2(\reg_pc[12] ),
    .B1(_18542_),
    .C1(_18551_),
    .X(_03940_));
 sky130_fd_sc_hd__inv_2 _21407_ (.A(\reg_pc[11] ),
    .Y(_18552_));
 sky130_fd_sc_hd__nand2_2 _21408_ (.A(_18494_),
    .B(_18552_),
    .Y(_18553_));
 sky130_fd_sc_hd__o211a_2 _21409_ (.A1(_18450_),
    .A2(_02589_),
    .B1(_18542_),
    .C1(_18553_),
    .X(_03939_));
 sky130_fd_sc_hd__inv_2 _21410_ (.A(_02588_),
    .Y(_18554_));
 sky130_fd_sc_hd__buf_1 _21411_ (.A(_18462_),
    .X(_18555_));
 sky130_fd_sc_hd__nand2_2 _21412_ (.A(_18554_),
    .B(_18555_),
    .Y(_18556_));
 sky130_fd_sc_hd__o211a_2 _21413_ (.A1(_18547_),
    .A2(\reg_pc[10] ),
    .B1(_18542_),
    .C1(_18556_),
    .X(_03938_));
 sky130_fd_sc_hd__buf_1 _21414_ (.A(_18497_),
    .X(_18557_));
 sky130_fd_sc_hd__inv_2 _21415_ (.A(_02587_),
    .Y(_18558_));
 sky130_fd_sc_hd__nand2_2 _21416_ (.A(_18558_),
    .B(_18555_),
    .Y(_18559_));
 sky130_fd_sc_hd__o211a_2 _21417_ (.A1(_18547_),
    .A2(\reg_pc[9] ),
    .B1(_18557_),
    .C1(_18559_),
    .X(_03937_));
 sky130_fd_sc_hd__inv_2 _21418_ (.A(_02586_),
    .Y(_18560_));
 sky130_fd_sc_hd__nand2_2 _21419_ (.A(_18560_),
    .B(_18555_),
    .Y(_18561_));
 sky130_fd_sc_hd__o211a_2 _21420_ (.A1(_18547_),
    .A2(\reg_pc[8] ),
    .B1(_18557_),
    .C1(_18561_),
    .X(_03936_));
 sky130_fd_sc_hd__inv_2 _21421_ (.A(_02585_),
    .Y(_18562_));
 sky130_fd_sc_hd__nand2_2 _21422_ (.A(_18562_),
    .B(_18555_),
    .Y(_18563_));
 sky130_fd_sc_hd__o211a_2 _21423_ (.A1(_18547_),
    .A2(\reg_pc[7] ),
    .B1(_18557_),
    .C1(_18563_),
    .X(_03935_));
 sky130_fd_sc_hd__inv_2 _21424_ (.A(\reg_pc[6] ),
    .Y(_18564_));
 sky130_fd_sc_hd__nand2_2 _21425_ (.A(_18494_),
    .B(_18564_),
    .Y(_18565_));
 sky130_fd_sc_hd__o211a_2 _21426_ (.A1(_18450_),
    .A2(_02584_),
    .B1(_18557_),
    .C1(_18565_),
    .X(_03934_));
 sky130_fd_sc_hd__inv_2 _21427_ (.A(_02583_),
    .Y(_18566_));
 sky130_fd_sc_hd__nand2_2 _21428_ (.A(_18566_),
    .B(_18555_),
    .Y(_18567_));
 sky130_fd_sc_hd__o211a_2 _21429_ (.A1(_18503_),
    .A2(\reg_pc[5] ),
    .B1(_18557_),
    .C1(_18567_),
    .X(_03933_));
 sky130_fd_sc_hd__nand2_2 _21430_ (.A(_18503_),
    .B(_01475_),
    .Y(_18568_));
 sky130_fd_sc_hd__o211a_2 _21431_ (.A1(_18503_),
    .A2(\reg_pc[4] ),
    .B1(_18557_),
    .C1(_18568_),
    .X(_03932_));
 sky130_fd_sc_hd__inv_2 _21432_ (.A(_01475_),
    .Y(_02582_));
 sky130_fd_sc_hd__buf_1 _21433_ (.A(_18497_),
    .X(_18569_));
 sky130_fd_sc_hd__inv_2 _21434_ (.A(_02571_),
    .Y(_18570_));
 sky130_fd_sc_hd__nand2_2 _21435_ (.A(_18570_),
    .B(_18555_),
    .Y(_18571_));
 sky130_fd_sc_hd__o211a_2 _21436_ (.A1(_18503_),
    .A2(\reg_pc[3] ),
    .B1(_18569_),
    .C1(_18571_),
    .X(_03931_));
 sky130_fd_sc_hd__inv_2 _21437_ (.A(_02560_),
    .Y(_01561_));
 sky130_fd_sc_hd__nand2_2 _21438_ (.A(_01561_),
    .B(_18454_),
    .Y(_18572_));
 sky130_fd_sc_hd__o211a_2 _21439_ (.A1(_18503_),
    .A2(\reg_pc[2] ),
    .B1(_18569_),
    .C1(_18572_),
    .X(_03930_));
 sky130_fd_sc_hd__inv_2 _21440_ (.A(\reg_pc[1] ),
    .Y(_18573_));
 sky130_fd_sc_hd__nand2_2 _21441_ (.A(_18494_),
    .B(_18573_),
    .Y(_18574_));
 sky130_fd_sc_hd__o211a_2 _21442_ (.A1(_18450_),
    .A2(_02590_),
    .B1(_18569_),
    .C1(_18574_),
    .X(_03929_));
 sky130_fd_sc_hd__inv_2 _21443_ (.A(\count_instr[61] ),
    .Y(_18575_));
 sky130_fd_sc_hd__and3_2 _21444_ (.A(\count_instr[58] ),
    .B(\count_instr[57] ),
    .C(\count_instr[56] ),
    .X(_18576_));
 sky130_fd_sc_hd__inv_2 _21445_ (.A(_18576_),
    .Y(_18577_));
 sky130_fd_sc_hd__inv_2 _21446_ (.A(\count_instr[62] ),
    .Y(_18578_));
 sky130_fd_sc_hd__inv_2 _21447_ (.A(\count_instr[60] ),
    .Y(_18579_));
 sky130_fd_sc_hd__inv_2 _21448_ (.A(\count_instr[59] ),
    .Y(_18580_));
 sky130_fd_sc_hd__nor2_2 _21449_ (.A(_18579_),
    .B(_18580_),
    .Y(_18581_));
 sky130_fd_sc_hd__inv_2 _21450_ (.A(_18581_),
    .Y(_18582_));
 sky130_fd_sc_hd__or3b_2 _21451_ (.A(_18578_),
    .B(_18582_),
    .C_N(\count_instr[63] ),
    .X(_18583_));
 sky130_fd_sc_hd__inv_2 _21452_ (.A(\count_instr[43] ),
    .Y(_18584_));
 sky130_fd_sc_hd__inv_2 _21453_ (.A(\count_instr[49] ),
    .Y(_18585_));
 sky130_fd_sc_hd__inv_2 _21454_ (.A(\count_instr[48] ),
    .Y(_18586_));
 sky130_fd_sc_hd__and3_2 _21455_ (.A(\count_instr[47] ),
    .B(\count_instr[46] ),
    .C(\count_instr[45] ),
    .X(_18587_));
 sky130_fd_sc_hd__nand2_2 _21456_ (.A(_18587_),
    .B(\count_instr[44] ),
    .Y(_18588_));
 sky130_fd_sc_hd__or3_2 _21457_ (.A(_18585_),
    .B(_18586_),
    .C(_18588_),
    .X(_18589_));
 sky130_fd_sc_hd__nand2_2 _21458_ (.A(\count_instr[36] ),
    .B(\count_instr[35] ),
    .Y(_18590_));
 sky130_fd_sc_hd__inv_2 _21459_ (.A(\count_instr[26] ),
    .Y(_18591_));
 sky130_fd_sc_hd__inv_2 _21460_ (.A(\count_instr[25] ),
    .Y(_18592_));
 sky130_fd_sc_hd__nand2_2 _21461_ (.A(\count_instr[15] ),
    .B(\count_instr[14] ),
    .Y(_18593_));
 sky130_fd_sc_hd__nand2_2 _21462_ (.A(\count_instr[4] ),
    .B(\count_instr[3] ),
    .Y(_18594_));
 sky130_fd_sc_hd__inv_2 _21463_ (.A(\count_instr[12] ),
    .Y(_18595_));
 sky130_fd_sc_hd__inv_2 _21464_ (.A(\count_instr[11] ),
    .Y(_18596_));
 sky130_fd_sc_hd__inv_2 _21465_ (.A(\count_instr[7] ),
    .Y(_18597_));
 sky130_fd_sc_hd__inv_2 _21466_ (.A(\count_instr[6] ),
    .Y(_18598_));
 sky130_fd_sc_hd__or4_2 _21467_ (.A(_18595_),
    .B(_18596_),
    .C(_18597_),
    .D(_18598_),
    .X(_18599_));
 sky130_fd_sc_hd__inv_2 _21468_ (.A(\count_instr[10] ),
    .Y(_18600_));
 sky130_fd_sc_hd__inv_2 _21469_ (.A(\count_instr[9] ),
    .Y(_18601_));
 sky130_fd_sc_hd__inv_2 _21470_ (.A(\count_instr[8] ),
    .Y(_18602_));
 sky130_fd_sc_hd__inv_2 _21471_ (.A(\count_instr[5] ),
    .Y(_18603_));
 sky130_fd_sc_hd__inv_2 _21472_ (.A(\count_instr[2] ),
    .Y(_18604_));
 sky130_fd_sc_hd__inv_2 _21473_ (.A(\count_instr[1] ),
    .Y(_18605_));
 sky130_fd_sc_hd__inv_2 _21474_ (.A(\count_instr[0] ),
    .Y(_18606_));
 sky130_fd_sc_hd__or4_2 _21475_ (.A(_18603_),
    .B(_18604_),
    .C(_18605_),
    .D(_18606_),
    .X(_18607_));
 sky130_fd_sc_hd__or4_2 _21476_ (.A(_18600_),
    .B(_18601_),
    .C(_18602_),
    .D(_18607_),
    .X(_18608_));
 sky130_fd_sc_hd__nor3_2 _21477_ (.A(_18594_),
    .B(_18599_),
    .C(_18608_),
    .Y(_18609_));
 sky130_fd_sc_hd__inv_2 _21478_ (.A(_18609_),
    .Y(_18610_));
 sky130_fd_sc_hd__or3b_2 _21479_ (.A(_18610_),
    .B(_18152_),
    .C_N(\count_instr[13] ),
    .X(_18611_));
 sky130_fd_sc_hd__nor2_2 _21480_ (.A(_18593_),
    .B(_18611_),
    .Y(_18612_));
 sky130_fd_sc_hd__and4_2 _21481_ (.A(_18612_),
    .B(\count_instr[18] ),
    .C(\count_instr[17] ),
    .D(\count_instr[16] ),
    .X(_18613_));
 sky130_fd_sc_hd__inv_2 _21482_ (.A(\count_instr[20] ),
    .Y(_18614_));
 sky130_fd_sc_hd__inv_2 _21483_ (.A(\count_instr[19] ),
    .Y(_18615_));
 sky130_fd_sc_hd__nor2_2 _21484_ (.A(_18614_),
    .B(_18615_),
    .Y(_18616_));
 sky130_fd_sc_hd__and4_2 _21485_ (.A(\count_instr[24] ),
    .B(\count_instr[23] ),
    .C(\count_instr[22] ),
    .D(\count_instr[21] ),
    .X(_18617_));
 sky130_fd_sc_hd__nand3_2 _21486_ (.A(_18613_),
    .B(_18616_),
    .C(_18617_),
    .Y(_18618_));
 sky130_fd_sc_hd__nor3_2 _21487_ (.A(_18591_),
    .B(_18592_),
    .C(_18618_),
    .Y(_18619_));
 sky130_fd_sc_hd__inv_2 _21488_ (.A(\count_instr[27] ),
    .Y(_18620_));
 sky130_fd_sc_hd__inv_2 _21489_ (.A(\count_instr[31] ),
    .Y(_18621_));
 sky130_fd_sc_hd__inv_2 _21490_ (.A(\count_instr[30] ),
    .Y(_18622_));
 sky130_fd_sc_hd__inv_2 _21491_ (.A(\count_instr[29] ),
    .Y(_18623_));
 sky130_fd_sc_hd__inv_2 _21492_ (.A(\count_instr[28] ),
    .Y(_18624_));
 sky130_fd_sc_hd__or4_2 _21493_ (.A(_18621_),
    .B(_18622_),
    .C(_18623_),
    .D(_18624_),
    .X(_18625_));
 sky130_fd_sc_hd__nor2_2 _21494_ (.A(_18620_),
    .B(_18625_),
    .Y(_18626_));
 sky130_fd_sc_hd__and3_2 _21495_ (.A(\count_instr[34] ),
    .B(\count_instr[33] ),
    .C(\count_instr[32] ),
    .X(_18627_));
 sky130_fd_sc_hd__nand3_2 _21496_ (.A(_18619_),
    .B(_18626_),
    .C(_18627_),
    .Y(_18628_));
 sky130_fd_sc_hd__nor2_2 _21497_ (.A(_18590_),
    .B(_18628_),
    .Y(_18629_));
 sky130_fd_sc_hd__and3_2 _21498_ (.A(\count_instr[39] ),
    .B(\count_instr[38] ),
    .C(\count_instr[37] ),
    .X(_18630_));
 sky130_fd_sc_hd__and3_2 _21499_ (.A(\count_instr[42] ),
    .B(\count_instr[41] ),
    .C(\count_instr[40] ),
    .X(_18631_));
 sky130_fd_sc_hd__nand3_2 _21500_ (.A(_18629_),
    .B(_18630_),
    .C(_18631_),
    .Y(_18632_));
 sky130_fd_sc_hd__nor3_2 _21501_ (.A(_18584_),
    .B(_18589_),
    .C(_18632_),
    .Y(_18633_));
 sky130_fd_sc_hd__and4_2 _21502_ (.A(_18633_),
    .B(\count_instr[52] ),
    .C(\count_instr[51] ),
    .D(\count_instr[50] ),
    .X(_18634_));
 sky130_fd_sc_hd__and3_2 _21503_ (.A(\count_instr[55] ),
    .B(\count_instr[54] ),
    .C(\count_instr[53] ),
    .X(_18635_));
 sky130_fd_sc_hd__nand2_2 _21504_ (.A(_18634_),
    .B(_18635_),
    .Y(_18636_));
 sky130_fd_sc_hd__buf_1 _21505_ (.A(_18025_),
    .X(_18637_));
 sky130_fd_sc_hd__buf_1 _21506_ (.A(_18637_),
    .X(_18638_));
 sky130_fd_sc_hd__o41ai_2 _21507_ (.A1(_18575_),
    .A2(_18577_),
    .A3(_18583_),
    .A4(_18636_),
    .B1(_18638_),
    .Y(_18639_));
 sky130_fd_sc_hd__and4_2 _21508_ (.A(_18634_),
    .B(\count_instr[59] ),
    .C(_18635_),
    .D(_18576_),
    .X(_18640_));
 sky130_fd_sc_hd__buf_1 _21509_ (.A(_18640_),
    .X(_18641_));
 sky130_fd_sc_hd__buf_1 _21510_ (.A(\count_instr[60] ),
    .X(_18642_));
 sky130_fd_sc_hd__nor2_2 _21511_ (.A(_18578_),
    .B(_18575_),
    .Y(_18643_));
 sky130_fd_sc_hd__a31oi_2 _21512_ (.A1(_18641_),
    .A2(_18642_),
    .A3(_18643_),
    .B1(\count_instr[63] ),
    .Y(_18644_));
 sky130_fd_sc_hd__nor2_2 _21513_ (.A(_18639_),
    .B(_18644_),
    .Y(_03928_));
 sky130_fd_sc_hd__nand3_2 _21514_ (.A(_18640_),
    .B(\count_instr[61] ),
    .C(_18642_),
    .Y(_18645_));
 sky130_fd_sc_hd__and3_2 _21515_ (.A(\count_instr[62] ),
    .B(\count_instr[61] ),
    .C(_18642_),
    .X(_18646_));
 sky130_fd_sc_hd__a21o_2 _21516_ (.A1(_18641_),
    .A2(_18646_),
    .B1(_18238_),
    .X(_18647_));
 sky130_fd_sc_hd__a21oi_2 _21517_ (.A1(_18645_),
    .A2(_18578_),
    .B1(_18647_),
    .Y(_03927_));
 sky130_fd_sc_hd__nand2_2 _21518_ (.A(_18641_),
    .B(_18642_),
    .Y(_18648_));
 sky130_fd_sc_hd__nand2_2 _21519_ (.A(_18645_),
    .B(_18638_),
    .Y(_18649_));
 sky130_fd_sc_hd__a21oi_2 _21520_ (.A1(_18575_),
    .A2(_18648_),
    .B1(_18649_),
    .Y(_03926_));
 sky130_fd_sc_hd__a21oi_2 _21521_ (.A1(_18641_),
    .A2(_18642_),
    .B1(_18349_),
    .Y(_18650_));
 sky130_fd_sc_hd__o21a_2 _21522_ (.A1(_18642_),
    .A2(_18641_),
    .B1(_18650_),
    .X(_03925_));
 sky130_fd_sc_hd__nor2_2 _21523_ (.A(_18577_),
    .B(_18636_),
    .Y(_18651_));
 sky130_fd_sc_hd__nor2_2 _21524_ (.A(_18331_),
    .B(_18641_),
    .Y(_18652_));
 sky130_fd_sc_hd__o21a_2 _21525_ (.A1(\count_instr[59] ),
    .A2(_18651_),
    .B1(_18652_),
    .X(_03924_));
 sky130_fd_sc_hd__inv_2 _21526_ (.A(\count_instr[57] ),
    .Y(_18653_));
 sky130_fd_sc_hd__inv_2 _21527_ (.A(\count_instr[56] ),
    .Y(_18654_));
 sky130_fd_sc_hd__nor2_2 _21528_ (.A(_18653_),
    .B(_18654_),
    .Y(_18655_));
 sky130_fd_sc_hd__a31o_2 _21529_ (.A1(_18634_),
    .A2(_18635_),
    .A3(_18655_),
    .B1(\count_instr[58] ),
    .X(_18656_));
 sky130_fd_sc_hd__o211a_2 _21530_ (.A1(_18636_),
    .A2(_18577_),
    .B1(_18569_),
    .C1(_18656_),
    .X(_03923_));
 sky130_fd_sc_hd__inv_2 _21531_ (.A(_18636_),
    .Y(_18657_));
 sky130_fd_sc_hd__nand2_2 _21532_ (.A(_18657_),
    .B(\count_instr[56] ),
    .Y(_18658_));
 sky130_fd_sc_hd__a31o_2 _21533_ (.A1(_18634_),
    .A2(_18635_),
    .A3(_18655_),
    .B1(_18238_),
    .X(_18659_));
 sky130_fd_sc_hd__a21oi_2 _21534_ (.A1(_18658_),
    .A2(_18653_),
    .B1(_18659_),
    .Y(_03922_));
 sky130_fd_sc_hd__buf_1 _21535_ (.A(_18027_),
    .X(_18660_));
 sky130_fd_sc_hd__nand2_2 _21536_ (.A(_18636_),
    .B(_18654_),
    .Y(_18661_));
 sky130_fd_sc_hd__and3_2 _21537_ (.A(_18658_),
    .B(_18660_),
    .C(_18661_),
    .X(_03921_));
 sky130_fd_sc_hd__inv_2 _21538_ (.A(\count_instr[54] ),
    .Y(_18662_));
 sky130_fd_sc_hd__nand2_2 _21539_ (.A(_18634_),
    .B(\count_instr[53] ),
    .Y(_18663_));
 sky130_fd_sc_hd__nor2_2 _21540_ (.A(_18662_),
    .B(_18663_),
    .Y(_18664_));
 sky130_fd_sc_hd__nor2_2 _21541_ (.A(_18331_),
    .B(_18657_),
    .Y(_18665_));
 sky130_fd_sc_hd__o21a_2 _21542_ (.A1(\count_instr[55] ),
    .A2(_18664_),
    .B1(_18665_),
    .X(_03920_));
 sky130_fd_sc_hd__buf_1 _21543_ (.A(_18637_),
    .X(_18666_));
 sky130_fd_sc_hd__nand2_2 _21544_ (.A(_18663_),
    .B(_18662_),
    .Y(_18667_));
 sky130_fd_sc_hd__and3b_2 _21545_ (.A_N(_18664_),
    .B(_18666_),
    .C(_18667_),
    .X(_03919_));
 sky130_fd_sc_hd__inv_2 _21546_ (.A(_18634_),
    .Y(_18668_));
 sky130_fd_sc_hd__inv_2 _21547_ (.A(\count_instr[53] ),
    .Y(_18669_));
 sky130_fd_sc_hd__nand2_2 _21548_ (.A(_18668_),
    .B(_18669_),
    .Y(_18670_));
 sky130_fd_sc_hd__buf_1 _21549_ (.A(_18027_),
    .X(_18671_));
 sky130_fd_sc_hd__and3_2 _21550_ (.A(_18670_),
    .B(_18671_),
    .C(_18663_),
    .X(_03918_));
 sky130_fd_sc_hd__inv_2 _21551_ (.A(\count_instr[51] ),
    .Y(_18672_));
 sky130_fd_sc_hd__nand2_2 _21552_ (.A(_18633_),
    .B(\count_instr[50] ),
    .Y(_18673_));
 sky130_fd_sc_hd__nor2_2 _21553_ (.A(_18672_),
    .B(_18673_),
    .Y(_18674_));
 sky130_fd_sc_hd__o211a_2 _21554_ (.A1(\count_instr[52] ),
    .A2(_18674_),
    .B1(_18569_),
    .C1(_18668_),
    .X(_03917_));
 sky130_fd_sc_hd__or2_2 _21555_ (.A(_18189_),
    .B(_18674_),
    .X(_18675_));
 sky130_fd_sc_hd__a21oi_2 _21556_ (.A1(_18672_),
    .A2(_18673_),
    .B1(_18675_),
    .Y(_03916_));
 sky130_fd_sc_hd__or2_2 _21557_ (.A(\count_instr[50] ),
    .B(_18633_),
    .X(_18676_));
 sky130_fd_sc_hd__and3_2 _21558_ (.A(_18676_),
    .B(_18671_),
    .C(_18673_),
    .X(_03915_));
 sky130_fd_sc_hd__or3_2 _21559_ (.A(_18584_),
    .B(_18588_),
    .C(_18632_),
    .X(_18677_));
 sky130_fd_sc_hd__or2_2 _21560_ (.A(_18586_),
    .B(_18677_),
    .X(_18678_));
 sky130_fd_sc_hd__or2_2 _21561_ (.A(_18189_),
    .B(_18633_),
    .X(_18679_));
 sky130_fd_sc_hd__a21oi_2 _21562_ (.A1(_18678_),
    .A2(_18585_),
    .B1(_18679_),
    .Y(_03914_));
 sky130_fd_sc_hd__nand2_2 _21563_ (.A(_18677_),
    .B(_18586_),
    .Y(_18680_));
 sky130_fd_sc_hd__and3_2 _21564_ (.A(_18678_),
    .B(_18671_),
    .C(_18680_),
    .X(_03913_));
 sky130_fd_sc_hd__inv_2 _21565_ (.A(\count_instr[45] ),
    .Y(_18681_));
 sky130_fd_sc_hd__nor2_2 _21566_ (.A(_18584_),
    .B(_18632_),
    .Y(_18682_));
 sky130_fd_sc_hd__nand2_2 _21567_ (.A(_18682_),
    .B(\count_instr[44] ),
    .Y(_18683_));
 sky130_fd_sc_hd__nor2_2 _21568_ (.A(_18681_),
    .B(_18683_),
    .Y(_18684_));
 sky130_fd_sc_hd__a21o_2 _21569_ (.A1(_18684_),
    .A2(\count_instr[46] ),
    .B1(\count_instr[47] ),
    .X(_18685_));
 sky130_fd_sc_hd__and3_2 _21570_ (.A(_18685_),
    .B(_18671_),
    .C(_18677_),
    .X(_03912_));
 sky130_fd_sc_hd__o21ai_2 _21571_ (.A1(\count_instr[46] ),
    .A2(_18684_),
    .B1(_18666_),
    .Y(_18686_));
 sky130_fd_sc_hd__a21oi_2 _21572_ (.A1(\count_instr[46] ),
    .A2(_18684_),
    .B1(_18686_),
    .Y(_03911_));
 sky130_fd_sc_hd__or2_2 _21573_ (.A(_18189_),
    .B(_18684_),
    .X(_18687_));
 sky130_fd_sc_hd__a21oi_2 _21574_ (.A1(_18681_),
    .A2(_18683_),
    .B1(_18687_),
    .Y(_03910_));
 sky130_fd_sc_hd__inv_2 _21575_ (.A(_18682_),
    .Y(_18688_));
 sky130_fd_sc_hd__inv_2 _21576_ (.A(\count_instr[44] ),
    .Y(_18689_));
 sky130_fd_sc_hd__nand2_2 _21577_ (.A(_18688_),
    .B(_18689_),
    .Y(_18690_));
 sky130_fd_sc_hd__and3_2 _21578_ (.A(_18690_),
    .B(_18671_),
    .C(_18683_),
    .X(_03909_));
 sky130_fd_sc_hd__nand2_2 _21579_ (.A(_18632_),
    .B(_18584_),
    .Y(_18691_));
 sky130_fd_sc_hd__and3_2 _21580_ (.A(_18688_),
    .B(_18671_),
    .C(_18691_),
    .X(_03908_));
 sky130_fd_sc_hd__buf_1 _21581_ (.A(\count_instr[37] ),
    .X(_18692_));
 sky130_fd_sc_hd__and4_2 _21582_ (.A(\count_instr[40] ),
    .B(\count_instr[39] ),
    .C(\count_instr[38] ),
    .D(_18692_),
    .X(_18693_));
 sky130_fd_sc_hd__a31o_2 _21583_ (.A1(_18629_),
    .A2(\count_instr[41] ),
    .A3(_18693_),
    .B1(\count_instr[42] ),
    .X(_18694_));
 sky130_fd_sc_hd__buf_1 _21584_ (.A(_18027_),
    .X(_18695_));
 sky130_fd_sc_hd__and3_2 _21585_ (.A(_18694_),
    .B(_18695_),
    .C(_18632_),
    .X(_03907_));
 sky130_fd_sc_hd__inv_2 _21586_ (.A(\count_instr[41] ),
    .Y(_18696_));
 sky130_fd_sc_hd__inv_2 _21587_ (.A(\count_instr[40] ),
    .Y(_18697_));
 sky130_fd_sc_hd__buf_1 _21588_ (.A(_18629_),
    .X(_18698_));
 sky130_fd_sc_hd__nand2_2 _21589_ (.A(_18698_),
    .B(_18630_),
    .Y(_18699_));
 sky130_fd_sc_hd__a21o_2 _21590_ (.A1(_18629_),
    .A2(_18693_),
    .B1(\count_instr[41] ),
    .X(_18700_));
 sky130_fd_sc_hd__o311a_2 _21591_ (.A1(_18696_),
    .A2(_18697_),
    .A3(_18699_),
    .B1(_18407_),
    .C1(_18700_),
    .X(_03906_));
 sky130_fd_sc_hd__a221oi_2 _21592_ (.A1(_18698_),
    .A2(_18693_),
    .B1(_18699_),
    .B2(_18697_),
    .C1(_18190_),
    .Y(_03905_));
 sky130_fd_sc_hd__and3_2 _21593_ (.A(_18629_),
    .B(\count_instr[38] ),
    .C(_18692_),
    .X(_18701_));
 sky130_fd_sc_hd__or2_2 _21594_ (.A(\count_instr[39] ),
    .B(_18701_),
    .X(_18702_));
 sky130_fd_sc_hd__and3_2 _21595_ (.A(_18702_),
    .B(_18695_),
    .C(_18699_),
    .X(_03904_));
 sky130_fd_sc_hd__a21oi_2 _21596_ (.A1(_18698_),
    .A2(_18692_),
    .B1(\count_instr[38] ),
    .Y(_18703_));
 sky130_fd_sc_hd__nor3_2 _21597_ (.A(_18190_),
    .B(_18703_),
    .C(_18701_),
    .Y(_03903_));
 sky130_fd_sc_hd__o21ai_2 _21598_ (.A1(_18692_),
    .A2(_18698_),
    .B1(_18638_),
    .Y(_18704_));
 sky130_fd_sc_hd__a21oi_2 _21599_ (.A1(_18692_),
    .A2(_18698_),
    .B1(_18704_),
    .Y(_03902_));
 sky130_fd_sc_hd__inv_2 _21600_ (.A(\count_instr[33] ),
    .Y(_18705_));
 sky130_fd_sc_hd__nand2_2 _21601_ (.A(_18619_),
    .B(\count_instr[27] ),
    .Y(_18706_));
 sky130_fd_sc_hd__nor2_2 _21602_ (.A(_18625_),
    .B(_18706_),
    .Y(_18707_));
 sky130_fd_sc_hd__nand2_2 _21603_ (.A(_18707_),
    .B(\count_instr[32] ),
    .Y(_18708_));
 sky130_fd_sc_hd__nor2_2 _21604_ (.A(_18705_),
    .B(_18708_),
    .Y(_18709_));
 sky130_fd_sc_hd__and3_2 _21605_ (.A(_18709_),
    .B(\count_instr[35] ),
    .C(\count_instr[34] ),
    .X(_18710_));
 sky130_fd_sc_hd__nor2_2 _21606_ (.A(_18331_),
    .B(_18698_),
    .Y(_18711_));
 sky130_fd_sc_hd__o21a_2 _21607_ (.A1(\count_instr[36] ),
    .A2(_18710_),
    .B1(_18711_),
    .X(_03901_));
 sky130_fd_sc_hd__inv_2 _21608_ (.A(_18628_),
    .Y(_18712_));
 sky130_fd_sc_hd__o21ai_2 _21609_ (.A1(\count_instr[35] ),
    .A2(_18712_),
    .B1(_18666_),
    .Y(_18713_));
 sky130_fd_sc_hd__nor2_2 _21610_ (.A(_18713_),
    .B(_18710_),
    .Y(_03900_));
 sky130_fd_sc_hd__inv_2 _21611_ (.A(_18709_),
    .Y(_18714_));
 sky130_fd_sc_hd__inv_2 _21612_ (.A(\count_instr[34] ),
    .Y(_18715_));
 sky130_fd_sc_hd__nand2_2 _21613_ (.A(_18714_),
    .B(_18715_),
    .Y(_18716_));
 sky130_fd_sc_hd__and3_2 _21614_ (.A(_18716_),
    .B(_18695_),
    .C(_18628_),
    .X(_03899_));
 sky130_fd_sc_hd__nand2_2 _21615_ (.A(_18708_),
    .B(_18705_),
    .Y(_18717_));
 sky130_fd_sc_hd__and3_2 _21616_ (.A(_18714_),
    .B(_18695_),
    .C(_18717_),
    .X(_03898_));
 sky130_fd_sc_hd__or2_2 _21617_ (.A(\count_instr[32] ),
    .B(_18707_),
    .X(_18718_));
 sky130_fd_sc_hd__and3_2 _21618_ (.A(_18718_),
    .B(_18695_),
    .C(_18708_),
    .X(_03897_));
 sky130_fd_sc_hd__or2_2 _21619_ (.A(_18624_),
    .B(_18706_),
    .X(_18719_));
 sky130_fd_sc_hd__or3_2 _21620_ (.A(_18622_),
    .B(_18623_),
    .C(_18719_),
    .X(_18720_));
 sky130_fd_sc_hd__buf_1 _21621_ (.A(_18051_),
    .X(_18721_));
 sky130_fd_sc_hd__or2_2 _21622_ (.A(_18721_),
    .B(_18707_),
    .X(_18722_));
 sky130_fd_sc_hd__a21oi_2 _21623_ (.A1(_18720_),
    .A2(_18621_),
    .B1(_18722_),
    .Y(_03896_));
 sky130_fd_sc_hd__nor2_2 _21624_ (.A(_18623_),
    .B(_18719_),
    .Y(_18723_));
 sky130_fd_sc_hd__o211a_2 _21625_ (.A1(\count_instr[30] ),
    .A2(_18723_),
    .B1(_18569_),
    .C1(_18720_),
    .X(_03895_));
 sky130_fd_sc_hd__or2_2 _21626_ (.A(_18721_),
    .B(_18723_),
    .X(_18724_));
 sky130_fd_sc_hd__a21oi_2 _21627_ (.A1(_18623_),
    .A2(_18719_),
    .B1(_18724_),
    .Y(_03894_));
 sky130_fd_sc_hd__nand2_2 _21628_ (.A(_18706_),
    .B(_18624_),
    .Y(_18725_));
 sky130_fd_sc_hd__and3_2 _21629_ (.A(_18719_),
    .B(_18695_),
    .C(_18725_),
    .X(_03893_));
 sky130_fd_sc_hd__inv_2 _21630_ (.A(_18619_),
    .Y(_18726_));
 sky130_fd_sc_hd__nand2_2 _21631_ (.A(_18726_),
    .B(_18620_),
    .Y(_18727_));
 sky130_fd_sc_hd__buf_1 _21632_ (.A(_18027_),
    .X(_18728_));
 sky130_fd_sc_hd__and3_2 _21633_ (.A(_18727_),
    .B(_18728_),
    .C(_18706_),
    .X(_03892_));
 sky130_fd_sc_hd__nor2_2 _21634_ (.A(_18592_),
    .B(_18618_),
    .Y(_18729_));
 sky130_fd_sc_hd__or2_2 _21635_ (.A(\count_instr[26] ),
    .B(_18729_),
    .X(_18730_));
 sky130_fd_sc_hd__and3_2 _21636_ (.A(_18730_),
    .B(_18728_),
    .C(_18726_),
    .X(_03891_));
 sky130_fd_sc_hd__or2_2 _21637_ (.A(_18721_),
    .B(_18729_),
    .X(_18731_));
 sky130_fd_sc_hd__a21oi_2 _21638_ (.A1(_18592_),
    .A2(_18618_),
    .B1(_18731_),
    .Y(_03890_));
 sky130_fd_sc_hd__inv_2 _21639_ (.A(\count_instr[23] ),
    .Y(_18732_));
 sky130_fd_sc_hd__inv_2 _21640_ (.A(\count_instr[22] ),
    .Y(_18733_));
 sky130_fd_sc_hd__nand2_2 _21641_ (.A(_18613_),
    .B(\count_instr[19] ),
    .Y(_18734_));
 sky130_fd_sc_hd__nor2_2 _21642_ (.A(_18614_),
    .B(_18734_),
    .Y(_18735_));
 sky130_fd_sc_hd__nand2_2 _21643_ (.A(_18735_),
    .B(\count_instr[21] ),
    .Y(_18736_));
 sky130_fd_sc_hd__or3_2 _21644_ (.A(_18732_),
    .B(_18733_),
    .C(_18736_),
    .X(_18737_));
 sky130_fd_sc_hd__inv_2 _21645_ (.A(\count_instr[24] ),
    .Y(_18738_));
 sky130_fd_sc_hd__nand2_2 _21646_ (.A(_18737_),
    .B(_18738_),
    .Y(_18739_));
 sky130_fd_sc_hd__and3_2 _21647_ (.A(_18739_),
    .B(_18728_),
    .C(_18618_),
    .X(_03889_));
 sky130_fd_sc_hd__nor2_2 _21648_ (.A(_18733_),
    .B(_18736_),
    .Y(_18740_));
 sky130_fd_sc_hd__buf_1 _21649_ (.A(_18026_),
    .X(_18741_));
 sky130_fd_sc_hd__buf_1 _21650_ (.A(_18741_),
    .X(_18742_));
 sky130_fd_sc_hd__o211a_2 _21651_ (.A1(\count_instr[23] ),
    .A2(_18740_),
    .B1(_18742_),
    .C1(_18737_),
    .X(_03888_));
 sky130_fd_sc_hd__or2_2 _21652_ (.A(_18721_),
    .B(_18740_),
    .X(_18743_));
 sky130_fd_sc_hd__a21oi_2 _21653_ (.A1(_18733_),
    .A2(_18736_),
    .B1(_18743_),
    .Y(_03887_));
 sky130_fd_sc_hd__or2_2 _21654_ (.A(\count_instr[21] ),
    .B(_18735_),
    .X(_18744_));
 sky130_fd_sc_hd__and3_2 _21655_ (.A(_18744_),
    .B(_18728_),
    .C(_18736_),
    .X(_03886_));
 sky130_fd_sc_hd__or2_2 _21656_ (.A(_18721_),
    .B(_18735_),
    .X(_18745_));
 sky130_fd_sc_hd__a21oi_2 _21657_ (.A1(_18614_),
    .A2(_18734_),
    .B1(_18745_),
    .Y(_03885_));
 sky130_fd_sc_hd__inv_2 _21658_ (.A(_18613_),
    .Y(_18746_));
 sky130_fd_sc_hd__nand2_2 _21659_ (.A(_18746_),
    .B(_18615_),
    .Y(_18747_));
 sky130_fd_sc_hd__and3_2 _21660_ (.A(_18747_),
    .B(_18728_),
    .C(_18734_),
    .X(_03884_));
 sky130_fd_sc_hd__inv_2 _21661_ (.A(\count_instr[17] ),
    .Y(_18748_));
 sky130_fd_sc_hd__nand2_2 _21662_ (.A(_18612_),
    .B(\count_instr[16] ),
    .Y(_18749_));
 sky130_fd_sc_hd__nor2_2 _21663_ (.A(_18748_),
    .B(_18749_),
    .Y(_18750_));
 sky130_fd_sc_hd__inv_2 _21664_ (.A(_18750_),
    .Y(_18751_));
 sky130_fd_sc_hd__inv_2 _21665_ (.A(\count_instr[18] ),
    .Y(_18752_));
 sky130_fd_sc_hd__nand2_2 _21666_ (.A(_18751_),
    .B(_18752_),
    .Y(_18753_));
 sky130_fd_sc_hd__and3_2 _21667_ (.A(_18753_),
    .B(_18728_),
    .C(_18746_),
    .X(_03883_));
 sky130_fd_sc_hd__buf_1 _21668_ (.A(_18027_),
    .X(_18754_));
 sky130_fd_sc_hd__nand2_2 _21669_ (.A(_18749_),
    .B(_18748_),
    .Y(_18755_));
 sky130_fd_sc_hd__and3_2 _21670_ (.A(_18751_),
    .B(_18754_),
    .C(_18755_),
    .X(_03882_));
 sky130_fd_sc_hd__inv_2 _21671_ (.A(_18612_),
    .Y(_18756_));
 sky130_fd_sc_hd__inv_2 _21672_ (.A(\count_instr[16] ),
    .Y(_18757_));
 sky130_fd_sc_hd__nand2_2 _21673_ (.A(_18756_),
    .B(_18757_),
    .Y(_18758_));
 sky130_fd_sc_hd__and3_2 _21674_ (.A(_18758_),
    .B(_18754_),
    .C(_18749_),
    .X(_03881_));
 sky130_fd_sc_hd__inv_2 _21675_ (.A(\count_instr[14] ),
    .Y(_18759_));
 sky130_fd_sc_hd__or2_2 _21676_ (.A(_18759_),
    .B(_18611_),
    .X(_18760_));
 sky130_fd_sc_hd__or2b_2 _21677_ (.A(\count_instr[15] ),
    .B_N(_18760_),
    .X(_18761_));
 sky130_fd_sc_hd__and3_2 _21678_ (.A(_18761_),
    .B(_18754_),
    .C(_18756_),
    .X(_03880_));
 sky130_fd_sc_hd__nand2_2 _21679_ (.A(_18611_),
    .B(_18759_),
    .Y(_18762_));
 sky130_fd_sc_hd__and3_2 _21680_ (.A(_18760_),
    .B(_18754_),
    .C(_18762_),
    .X(_03879_));
 sky130_fd_sc_hd__nor2_2 _21681_ (.A(_18610_),
    .B(_18152_),
    .Y(_18763_));
 sky130_fd_sc_hd__o211a_2 _21682_ (.A1(\count_instr[13] ),
    .A2(_18763_),
    .B1(_18742_),
    .C1(_18611_),
    .X(_03878_));
 sky130_fd_sc_hd__nand2_2 _21683_ (.A(_18153_),
    .B(\count_instr[0] ),
    .Y(_18764_));
 sky130_fd_sc_hd__or2_2 _21684_ (.A(_18605_),
    .B(_18764_),
    .X(_18765_));
 sky130_fd_sc_hd__or2_2 _21685_ (.A(_18604_),
    .B(_18765_),
    .X(_18766_));
 sky130_fd_sc_hd__or2_2 _21686_ (.A(_18594_),
    .B(_18766_),
    .X(_18767_));
 sky130_fd_sc_hd__nor2_2 _21687_ (.A(_18603_),
    .B(_18767_),
    .Y(_18768_));
 sky130_fd_sc_hd__nand2_2 _21688_ (.A(_18768_),
    .B(\count_instr[6] ),
    .Y(_18769_));
 sky130_fd_sc_hd__nor2_2 _21689_ (.A(_18597_),
    .B(_18769_),
    .Y(_18770_));
 sky130_fd_sc_hd__nand2_2 _21690_ (.A(_18770_),
    .B(\count_instr[8] ),
    .Y(_18771_));
 sky130_fd_sc_hd__nor2_2 _21691_ (.A(_18601_),
    .B(_18771_),
    .Y(_18772_));
 sky130_fd_sc_hd__nand2_2 _21692_ (.A(_18772_),
    .B(\count_instr[10] ),
    .Y(_18773_));
 sky130_fd_sc_hd__or2_2 _21693_ (.A(_18596_),
    .B(_18773_),
    .X(_18774_));
 sky130_fd_sc_hd__a211oi_2 _21694_ (.A1(_18774_),
    .A2(_18595_),
    .B1(_18190_),
    .C1(_18763_),
    .Y(_03877_));
 sky130_fd_sc_hd__nand2_2 _21695_ (.A(_18773_),
    .B(_18596_),
    .Y(_18775_));
 sky130_fd_sc_hd__and3_2 _21696_ (.A(_18774_),
    .B(_18754_),
    .C(_18775_),
    .X(_03876_));
 sky130_fd_sc_hd__inv_2 _21697_ (.A(_18772_),
    .Y(_18776_));
 sky130_fd_sc_hd__nand2_2 _21698_ (.A(_18776_),
    .B(_18600_),
    .Y(_18777_));
 sky130_fd_sc_hd__and3_2 _21699_ (.A(_18777_),
    .B(_18754_),
    .C(_18773_),
    .X(_03875_));
 sky130_fd_sc_hd__buf_1 _21700_ (.A(_18025_),
    .X(_18778_));
 sky130_fd_sc_hd__buf_1 _21701_ (.A(_18778_),
    .X(_18779_));
 sky130_fd_sc_hd__nand2_2 _21702_ (.A(_18771_),
    .B(_18601_),
    .Y(_18780_));
 sky130_fd_sc_hd__and3_2 _21703_ (.A(_18776_),
    .B(_18779_),
    .C(_18780_),
    .X(_03874_));
 sky130_fd_sc_hd__inv_2 _21704_ (.A(_18770_),
    .Y(_18781_));
 sky130_fd_sc_hd__nand2_2 _21705_ (.A(_18781_),
    .B(_18602_),
    .Y(_18782_));
 sky130_fd_sc_hd__and3_2 _21706_ (.A(_18782_),
    .B(_18779_),
    .C(_18771_),
    .X(_03873_));
 sky130_fd_sc_hd__nand2_2 _21707_ (.A(_18769_),
    .B(_18597_),
    .Y(_18783_));
 sky130_fd_sc_hd__and3_2 _21708_ (.A(_18781_),
    .B(_18779_),
    .C(_18783_),
    .X(_03872_));
 sky130_fd_sc_hd__inv_2 _21709_ (.A(_18768_),
    .Y(_18784_));
 sky130_fd_sc_hd__nand2_2 _21710_ (.A(_18784_),
    .B(_18598_),
    .Y(_18785_));
 sky130_fd_sc_hd__and3_2 _21711_ (.A(_18785_),
    .B(_18779_),
    .C(_18769_),
    .X(_03871_));
 sky130_fd_sc_hd__nand2_2 _21712_ (.A(_18767_),
    .B(_18603_),
    .Y(_18786_));
 sky130_fd_sc_hd__and3_2 _21713_ (.A(_18784_),
    .B(_18779_),
    .C(_18786_),
    .X(_03870_));
 sky130_fd_sc_hd__inv_2 _21714_ (.A(\count_instr[3] ),
    .Y(_18787_));
 sky130_fd_sc_hd__or2_2 _21715_ (.A(_18787_),
    .B(_18766_),
    .X(_18788_));
 sky130_fd_sc_hd__inv_2 _21716_ (.A(\count_instr[4] ),
    .Y(_18789_));
 sky130_fd_sc_hd__nand2_2 _21717_ (.A(_18788_),
    .B(_18789_),
    .Y(_18790_));
 sky130_fd_sc_hd__and3_2 _21718_ (.A(_18790_),
    .B(_18779_),
    .C(_18767_),
    .X(_03869_));
 sky130_fd_sc_hd__buf_1 _21719_ (.A(_18778_),
    .X(_18791_));
 sky130_fd_sc_hd__nand2_2 _21720_ (.A(_18766_),
    .B(_18787_),
    .Y(_18792_));
 sky130_fd_sc_hd__and3_2 _21721_ (.A(_18788_),
    .B(_18791_),
    .C(_18792_),
    .X(_03868_));
 sky130_fd_sc_hd__nand2_2 _21722_ (.A(_18765_),
    .B(_18604_),
    .Y(_18793_));
 sky130_fd_sc_hd__and3_2 _21723_ (.A(_18766_),
    .B(_18791_),
    .C(_18793_),
    .X(_03867_));
 sky130_fd_sc_hd__nand2_2 _21724_ (.A(_18764_),
    .B(_18605_),
    .Y(_18794_));
 sky130_fd_sc_hd__and3_2 _21725_ (.A(_18765_),
    .B(_18791_),
    .C(_18794_),
    .X(_03866_));
 sky130_fd_sc_hd__nand2_2 _21726_ (.A(_18152_),
    .B(_18606_),
    .Y(_18795_));
 sky130_fd_sc_hd__and3_2 _21727_ (.A(_18764_),
    .B(_18791_),
    .C(_18795_),
    .X(_03865_));
 sky130_fd_sc_hd__and3_2 _21728_ (.A(_18233_),
    .B(_18034_),
    .C(_18258_),
    .X(_18796_));
 sky130_fd_sc_hd__buf_1 _21729_ (.A(_18796_),
    .X(_18797_));
 sky130_fd_sc_hd__buf_1 _21730_ (.A(_18797_),
    .X(_18798_));
 sky130_fd_sc_hd__buf_1 _21731_ (.A(_18193_),
    .X(_18799_));
 sky130_fd_sc_hd__buf_1 _21732_ (.A(_18799_),
    .X(_18800_));
 sky130_fd_sc_hd__inv_2 _21733_ (.A(_18796_),
    .Y(_18801_));
 sky130_fd_sc_hd__buf_1 _21734_ (.A(_18801_),
    .X(_18802_));
 sky130_fd_sc_hd__buf_1 _21735_ (.A(_18802_),
    .X(_18803_));
 sky130_fd_sc_hd__a21o_2 _21736_ (.A1(_18800_),
    .A2(_18130_),
    .B1(_18803_),
    .X(_18804_));
 sky130_fd_sc_hd__o211a_2 _21737_ (.A1(eoi[31]),
    .A2(_18798_),
    .B1(_18742_),
    .C1(_18804_),
    .X(_03864_));
 sky130_fd_sc_hd__a21o_2 _21738_ (.A1(_18800_),
    .A2(_18132_),
    .B1(_18803_),
    .X(_18805_));
 sky130_fd_sc_hd__o211a_2 _21739_ (.A1(eoi[30]),
    .A2(_18798_),
    .B1(_18742_),
    .C1(_18805_),
    .X(_03863_));
 sky130_fd_sc_hd__buf_1 _21740_ (.A(_18194_),
    .X(_18806_));
 sky130_fd_sc_hd__buf_1 _21741_ (.A(_18801_),
    .X(_18807_));
 sky130_fd_sc_hd__a31o_2 _21742_ (.A1(_18126_),
    .A2(_18806_),
    .A3(\irq_pending[29] ),
    .B1(_18807_),
    .X(_18808_));
 sky130_fd_sc_hd__o211a_2 _21743_ (.A1(eoi[29]),
    .A2(_18798_),
    .B1(_18742_),
    .C1(_18808_),
    .X(_03862_));
 sky130_fd_sc_hd__buf_1 _21744_ (.A(_18799_),
    .X(_18809_));
 sky130_fd_sc_hd__a21o_2 _21745_ (.A1(_18809_),
    .A2(_18128_),
    .B1(_18803_),
    .X(_18810_));
 sky130_fd_sc_hd__o211a_2 _21746_ (.A1(eoi[28]),
    .A2(_18798_),
    .B1(_18742_),
    .C1(_18810_),
    .X(_03861_));
 sky130_fd_sc_hd__buf_1 _21747_ (.A(_18741_),
    .X(_18811_));
 sky130_fd_sc_hd__a21o_2 _21748_ (.A1(_18809_),
    .A2(_18097_),
    .B1(_18803_),
    .X(_18812_));
 sky130_fd_sc_hd__o211a_2 _21749_ (.A1(eoi[27]),
    .A2(_18798_),
    .B1(_18811_),
    .C1(_18812_),
    .X(_03860_));
 sky130_fd_sc_hd__a21o_2 _21750_ (.A1(_18809_),
    .A2(_18098_),
    .B1(_18803_),
    .X(_18813_));
 sky130_fd_sc_hd__o211a_2 _21751_ (.A1(eoi[26]),
    .A2(_18798_),
    .B1(_18811_),
    .C1(_18813_),
    .X(_03859_));
 sky130_fd_sc_hd__buf_1 _21752_ (.A(_18797_),
    .X(_18814_));
 sky130_fd_sc_hd__a31o_2 _21753_ (.A1(_18099_),
    .A2(_18806_),
    .A3(\irq_pending[25] ),
    .B1(_18807_),
    .X(_18815_));
 sky130_fd_sc_hd__o211a_2 _21754_ (.A1(eoi[25]),
    .A2(_18814_),
    .B1(_18811_),
    .C1(_18815_),
    .X(_03858_));
 sky130_fd_sc_hd__a31o_2 _21755_ (.A1(_18100_),
    .A2(_18806_),
    .A3(\irq_pending[24] ),
    .B1(_18807_),
    .X(_18816_));
 sky130_fd_sc_hd__o211a_2 _21756_ (.A1(eoi[24]),
    .A2(_18814_),
    .B1(_18811_),
    .C1(_18816_),
    .X(_03857_));
 sky130_fd_sc_hd__a21o_2 _21757_ (.A1(_18809_),
    .A2(_18104_),
    .B1(_18803_),
    .X(_18817_));
 sky130_fd_sc_hd__o211a_2 _21758_ (.A1(eoi[23]),
    .A2(_18814_),
    .B1(_18811_),
    .C1(_18817_),
    .X(_03856_));
 sky130_fd_sc_hd__buf_1 _21759_ (.A(_18802_),
    .X(_18818_));
 sky130_fd_sc_hd__a21o_2 _21760_ (.A1(_18809_),
    .A2(_18106_),
    .B1(_18818_),
    .X(_18819_));
 sky130_fd_sc_hd__o211a_2 _21761_ (.A1(eoi[22]),
    .A2(_18814_),
    .B1(_18811_),
    .C1(_18819_),
    .X(_03855_));
 sky130_fd_sc_hd__buf_1 _21762_ (.A(_18741_),
    .X(_18820_));
 sky130_fd_sc_hd__a31o_2 _21763_ (.A1(_18107_),
    .A2(_18806_),
    .A3(\irq_pending[21] ),
    .B1(_18807_),
    .X(_18821_));
 sky130_fd_sc_hd__o211a_2 _21764_ (.A1(eoi[21]),
    .A2(_18814_),
    .B1(_18820_),
    .C1(_18821_),
    .X(_03854_));
 sky130_fd_sc_hd__buf_1 _21765_ (.A(_18802_),
    .X(_18822_));
 sky130_fd_sc_hd__a31o_2 _21766_ (.A1(_18108_),
    .A2(_18806_),
    .A3(\irq_pending[20] ),
    .B1(_18822_),
    .X(_18823_));
 sky130_fd_sc_hd__o211a_2 _21767_ (.A1(eoi[20]),
    .A2(_18814_),
    .B1(_18820_),
    .C1(_18823_),
    .X(_03853_));
 sky130_fd_sc_hd__buf_1 _21768_ (.A(_18797_),
    .X(_18824_));
 sky130_fd_sc_hd__a21o_2 _21769_ (.A1(_18809_),
    .A2(_18093_),
    .B1(_18818_),
    .X(_18825_));
 sky130_fd_sc_hd__o211a_2 _21770_ (.A1(eoi[19]),
    .A2(_18824_),
    .B1(_18820_),
    .C1(_18825_),
    .X(_03852_));
 sky130_fd_sc_hd__buf_1 _21771_ (.A(_18799_),
    .X(_18826_));
 sky130_fd_sc_hd__a21o_2 _21772_ (.A1(_18826_),
    .A2(_18095_),
    .B1(_18818_),
    .X(_18827_));
 sky130_fd_sc_hd__o211a_2 _21773_ (.A1(eoi[18]),
    .A2(_18824_),
    .B1(_18820_),
    .C1(_18827_),
    .X(_03851_));
 sky130_fd_sc_hd__buf_1 _21774_ (.A(_18194_),
    .X(_18828_));
 sky130_fd_sc_hd__a31o_2 _21775_ (.A1(_18089_),
    .A2(_18828_),
    .A3(\irq_pending[17] ),
    .B1(_18822_),
    .X(_18829_));
 sky130_fd_sc_hd__o211a_2 _21776_ (.A1(eoi[17]),
    .A2(_18824_),
    .B1(_18820_),
    .C1(_18829_),
    .X(_03850_));
 sky130_fd_sc_hd__a21o_2 _21777_ (.A1(_18826_),
    .A2(_18091_),
    .B1(_18818_),
    .X(_18830_));
 sky130_fd_sc_hd__o211a_2 _21778_ (.A1(eoi[16]),
    .A2(_18824_),
    .B1(_18820_),
    .C1(_18830_),
    .X(_03849_));
 sky130_fd_sc_hd__buf_1 _21779_ (.A(_18741_),
    .X(_18831_));
 sky130_fd_sc_hd__a21o_2 _21780_ (.A1(_18826_),
    .A2(_18138_),
    .B1(_18818_),
    .X(_18832_));
 sky130_fd_sc_hd__o211a_2 _21781_ (.A1(eoi[15]),
    .A2(_18824_),
    .B1(_18831_),
    .C1(_18832_),
    .X(_03848_));
 sky130_fd_sc_hd__a21o_2 _21782_ (.A1(_18826_),
    .A2(_18140_),
    .B1(_18818_),
    .X(_18833_));
 sky130_fd_sc_hd__o211a_2 _21783_ (.A1(eoi[14]),
    .A2(_18824_),
    .B1(_18831_),
    .C1(_18833_),
    .X(_03847_));
 sky130_fd_sc_hd__buf_1 _21784_ (.A(_18797_),
    .X(_18834_));
 sky130_fd_sc_hd__a31o_2 _21785_ (.A1(_18134_),
    .A2(_18828_),
    .A3(\irq_pending[13] ),
    .B1(_18822_),
    .X(_18835_));
 sky130_fd_sc_hd__o211a_2 _21786_ (.A1(eoi[13]),
    .A2(_18834_),
    .B1(_18831_),
    .C1(_18835_),
    .X(_03846_));
 sky130_fd_sc_hd__buf_1 _21787_ (.A(_18802_),
    .X(_18836_));
 sky130_fd_sc_hd__a21o_2 _21788_ (.A1(_18826_),
    .A2(_18136_),
    .B1(_18836_),
    .X(_18837_));
 sky130_fd_sc_hd__o211a_2 _21789_ (.A1(eoi[12]),
    .A2(_18834_),
    .B1(_18831_),
    .C1(_18837_),
    .X(_03845_));
 sky130_fd_sc_hd__a21o_2 _21790_ (.A1(_18826_),
    .A2(_18112_),
    .B1(_18836_),
    .X(_18838_));
 sky130_fd_sc_hd__o211a_2 _21791_ (.A1(eoi[11]),
    .A2(_18834_),
    .B1(_18831_),
    .C1(_18838_),
    .X(_03844_));
 sky130_fd_sc_hd__buf_1 _21792_ (.A(_18799_),
    .X(_18839_));
 sky130_fd_sc_hd__a21o_2 _21793_ (.A1(_18839_),
    .A2(_18113_),
    .B1(_18836_),
    .X(_18840_));
 sky130_fd_sc_hd__o211a_2 _21794_ (.A1(eoi[10]),
    .A2(_18834_),
    .B1(_18831_),
    .C1(_18840_),
    .X(_03843_));
 sky130_fd_sc_hd__buf_1 _21795_ (.A(_18741_),
    .X(_18841_));
 sky130_fd_sc_hd__a31o_2 _21796_ (.A1(_18114_),
    .A2(_18828_),
    .A3(\irq_pending[9] ),
    .B1(_18822_),
    .X(_18842_));
 sky130_fd_sc_hd__o211a_2 _21797_ (.A1(eoi[9]),
    .A2(_18834_),
    .B1(_18841_),
    .C1(_18842_),
    .X(_03842_));
 sky130_fd_sc_hd__a31o_2 _21798_ (.A1(_18115_),
    .A2(_18828_),
    .A3(\irq_pending[8] ),
    .B1(_18822_),
    .X(_18843_));
 sky130_fd_sc_hd__o211a_2 _21799_ (.A1(eoi[8]),
    .A2(_18834_),
    .B1(_18841_),
    .C1(_18843_),
    .X(_03841_));
 sky130_fd_sc_hd__buf_1 _21800_ (.A(_18796_),
    .X(_18844_));
 sky130_fd_sc_hd__a21o_2 _21801_ (.A1(_18839_),
    .A2(_18119_),
    .B1(_18836_),
    .X(_18845_));
 sky130_fd_sc_hd__o211a_2 _21802_ (.A1(eoi[7]),
    .A2(_18844_),
    .B1(_18841_),
    .C1(_18845_),
    .X(_03840_));
 sky130_fd_sc_hd__a21o_2 _21803_ (.A1(_18839_),
    .A2(_18121_),
    .B1(_18836_),
    .X(_18846_));
 sky130_fd_sc_hd__o211a_2 _21804_ (.A1(eoi[6]),
    .A2(_18844_),
    .B1(_18841_),
    .C1(_18846_),
    .X(_03839_));
 sky130_fd_sc_hd__a31o_2 _21805_ (.A1(_18122_),
    .A2(_18828_),
    .A3(\irq_pending[5] ),
    .B1(_18822_),
    .X(_18847_));
 sky130_fd_sc_hd__o211a_2 _21806_ (.A1(eoi[5]),
    .A2(_18844_),
    .B1(_18841_),
    .C1(_18847_),
    .X(_03838_));
 sky130_fd_sc_hd__a31o_2 _21807_ (.A1(_18123_),
    .A2(_18828_),
    .A3(\irq_pending[4] ),
    .B1(_18802_),
    .X(_18848_));
 sky130_fd_sc_hd__o211a_2 _21808_ (.A1(eoi[4]),
    .A2(_18844_),
    .B1(_18841_),
    .C1(_18848_),
    .X(_03837_));
 sky130_fd_sc_hd__buf_1 _21809_ (.A(_18741_),
    .X(_18849_));
 sky130_fd_sc_hd__a21o_2 _21810_ (.A1(_18839_),
    .A2(_18087_),
    .B1(_18836_),
    .X(_18850_));
 sky130_fd_sc_hd__o211a_2 _21811_ (.A1(eoi[3]),
    .A2(_18844_),
    .B1(_18849_),
    .C1(_18850_),
    .X(_03836_));
 sky130_fd_sc_hd__buf_1 _21812_ (.A(_18194_),
    .X(_18851_));
 sky130_fd_sc_hd__a31o_2 _21813_ (.A1(_18081_),
    .A2(_18851_),
    .A3(\irq_pending[2] ),
    .B1(_18802_),
    .X(_18852_));
 sky130_fd_sc_hd__o211a_2 _21814_ (.A1(eoi[2]),
    .A2(_18844_),
    .B1(_18849_),
    .C1(_18852_),
    .X(_03835_));
 sky130_fd_sc_hd__a21o_2 _21815_ (.A1(_18839_),
    .A2(_18085_),
    .B1(_18807_),
    .X(_18853_));
 sky130_fd_sc_hd__o211a_2 _21816_ (.A1(eoi[1]),
    .A2(_18797_),
    .B1(_18849_),
    .C1(_18853_),
    .X(_03834_));
 sky130_fd_sc_hd__a21o_2 _21817_ (.A1(_18839_),
    .A2(_18083_),
    .B1(_18807_),
    .X(_18854_));
 sky130_fd_sc_hd__o211a_2 _21818_ (.A1(eoi[0]),
    .A2(_18797_),
    .B1(_18849_),
    .C1(_18854_),
    .X(_03833_));
 sky130_fd_sc_hd__nor2_2 _21819_ (.A(instr_ecall_ebreak),
    .B(pcpi_timeout),
    .Y(_00311_));
 sky130_fd_sc_hd__inv_2 _21820_ (.A(_00311_),
    .Y(_18855_));
 sky130_fd_sc_hd__nor2_2 _21821_ (.A(_18227_),
    .B(_18246_),
    .Y(_18856_));
 sky130_fd_sc_hd__inv_2 _21822_ (.A(_18856_),
    .Y(_18857_));
 sky130_fd_sc_hd__or3_2 _21823_ (.A(\pcpi_mul.active[1] ),
    .B(_18855_),
    .C(_18857_),
    .X(_18858_));
 sky130_fd_sc_hd__nand2_2 _21824_ (.A(_18857_),
    .B(pcpi_valid),
    .Y(_18859_));
 sky130_fd_sc_hd__a21oi_2 _21825_ (.A1(_18858_),
    .A2(_18859_),
    .B1(_18245_),
    .Y(_03832_));
 sky130_fd_sc_hd__a21oi_2 _21826_ (.A1(_18045_),
    .A2(_18009_),
    .B1(_18005_),
    .Y(_18860_));
 sky130_fd_sc_hd__o21ai_2 _21827_ (.A1(_18860_),
    .A2(_18335_),
    .B1(_18047_),
    .Y(_18861_));
 sky130_fd_sc_hd__nand2_2 _21828_ (.A(_18006_),
    .B(mem_valid),
    .Y(_18862_));
 sky130_fd_sc_hd__a21oi_2 _21829_ (.A1(_18861_),
    .A2(_18862_),
    .B1(_18190_),
    .Y(_03831_));
 sky130_fd_sc_hd__or4_2 _21830_ (.A(\irq_pending[25] ),
    .B(\irq_pending[24] ),
    .C(\irq_pending[27] ),
    .D(\irq_pending[26] ),
    .X(_18863_));
 sky130_fd_sc_hd__or4_2 _21831_ (.A(\irq_pending[21] ),
    .B(\irq_pending[20] ),
    .C(\irq_pending[23] ),
    .D(\irq_pending[22] ),
    .X(_18864_));
 sky130_fd_sc_hd__or4_2 _21832_ (.A(\irq_pending[17] ),
    .B(\irq_pending[16] ),
    .C(\irq_pending[19] ),
    .D(\irq_pending[18] ),
    .X(_18865_));
 sky130_fd_sc_hd__or4_2 _21833_ (.A(\irq_pending[29] ),
    .B(\irq_pending[28] ),
    .C(\irq_pending[31] ),
    .D(\irq_pending[30] ),
    .X(_18866_));
 sky130_fd_sc_hd__or4_2 _21834_ (.A(_18863_),
    .B(_18864_),
    .C(_18865_),
    .D(_18866_),
    .X(_18867_));
 sky130_fd_sc_hd__or4_2 _21835_ (.A(\irq_pending[9] ),
    .B(\irq_pending[8] ),
    .C(\irq_pending[11] ),
    .D(\irq_pending[10] ),
    .X(_18868_));
 sky130_fd_sc_hd__or4_2 _21836_ (.A(\irq_pending[5] ),
    .B(\irq_pending[4] ),
    .C(\irq_pending[7] ),
    .D(\irq_pending[6] ),
    .X(_18869_));
 sky130_fd_sc_hd__or4_2 _21837_ (.A(\irq_pending[1] ),
    .B(\irq_pending[0] ),
    .C(\irq_pending[3] ),
    .D(\irq_pending[2] ),
    .X(_18870_));
 sky130_fd_sc_hd__or4_2 _21838_ (.A(\irq_pending[13] ),
    .B(\irq_pending[12] ),
    .C(\irq_pending[15] ),
    .D(\irq_pending[14] ),
    .X(_18871_));
 sky130_fd_sc_hd__or4_2 _21839_ (.A(_18868_),
    .B(_18869_),
    .C(_18870_),
    .D(_18871_),
    .X(_18872_));
 sky130_fd_sc_hd__nor2_2 _21840_ (.A(_18867_),
    .B(_18872_),
    .Y(_02410_));
 sky130_fd_sc_hd__buf_1 _21841_ (.A(_18146_),
    .X(_00308_));
 sky130_fd_sc_hd__nor2_2 _21842_ (.A(_18017_),
    .B(_00308_),
    .Y(_18873_));
 sky130_fd_sc_hd__inv_2 _21843_ (.A(_18873_),
    .Y(_18874_));
 sky130_fd_sc_hd__nor2_2 _21844_ (.A(_18150_),
    .B(_18874_),
    .Y(_18875_));
 sky130_fd_sc_hd__and3_2 _21845_ (.A(_18875_),
    .B(_18501_),
    .C(_02410_),
    .X(_03830_));
 sky130_fd_sc_hd__or4b_2 _21846_ (.A(_18338_),
    .B(instr_sltu),
    .C(instr_slt),
    .D_N(_18211_),
    .X(_18876_));
 sky130_fd_sc_hd__buf_1 _21847_ (.A(_18392_),
    .X(_18877_));
 sky130_fd_sc_hd__and3_2 _21848_ (.A(_18876_),
    .B(_18791_),
    .C(_18877_),
    .X(_03829_));
 sky130_fd_sc_hd__or2_2 _21849_ (.A(_18015_),
    .B(_18014_),
    .X(_18878_));
 sky130_fd_sc_hd__nor3_2 _21850_ (.A(_18017_),
    .B(_00297_),
    .C(_18878_),
    .Y(_03828_));
 sky130_fd_sc_hd__and2_2 _21851_ (.A(_18442_),
    .B(_18407_),
    .X(_03827_));
 sky130_fd_sc_hd__buf_1 _21852_ (.A(_18395_),
    .X(_18879_));
 sky130_fd_sc_hd__and2_2 _21853_ (.A(_18879_),
    .B(_02435_),
    .X(_03826_));
 sky130_fd_sc_hd__and2_2 _21854_ (.A(_18879_),
    .B(_02434_),
    .X(_03825_));
 sky130_fd_sc_hd__and2_2 _21855_ (.A(_18879_),
    .B(_02432_),
    .X(_03824_));
 sky130_fd_sc_hd__and2_2 _21856_ (.A(_18879_),
    .B(_02431_),
    .X(_03823_));
 sky130_fd_sc_hd__and2_2 _21857_ (.A(_18879_),
    .B(_02430_),
    .X(_03822_));
 sky130_fd_sc_hd__buf_1 _21858_ (.A(_18026_),
    .X(_18880_));
 sky130_fd_sc_hd__buf_1 _21859_ (.A(_18880_),
    .X(_18881_));
 sky130_fd_sc_hd__and2_2 _21860_ (.A(_18881_),
    .B(_02429_),
    .X(_03821_));
 sky130_fd_sc_hd__and2_2 _21861_ (.A(_18881_),
    .B(_02428_),
    .X(_03820_));
 sky130_fd_sc_hd__and2_2 _21862_ (.A(_18881_),
    .B(_02427_),
    .X(_03819_));
 sky130_fd_sc_hd__and2_2 _21863_ (.A(_18881_),
    .B(_02426_),
    .X(_03818_));
 sky130_fd_sc_hd__and2_2 _21864_ (.A(_18881_),
    .B(_02425_),
    .X(_03817_));
 sky130_fd_sc_hd__and2_2 _21865_ (.A(_18881_),
    .B(_02424_),
    .X(_03816_));
 sky130_fd_sc_hd__buf_1 _21866_ (.A(_18880_),
    .X(_18882_));
 sky130_fd_sc_hd__and2_2 _21867_ (.A(_18882_),
    .B(_02423_),
    .X(_03815_));
 sky130_fd_sc_hd__and2_2 _21868_ (.A(_18882_),
    .B(_02421_),
    .X(_03814_));
 sky130_fd_sc_hd__and2_2 _21869_ (.A(_18882_),
    .B(_02420_),
    .X(_03813_));
 sky130_fd_sc_hd__and2_2 _21870_ (.A(_18882_),
    .B(_02419_),
    .X(_03812_));
 sky130_fd_sc_hd__and2_2 _21871_ (.A(_18882_),
    .B(_02418_),
    .X(_03811_));
 sky130_fd_sc_hd__and2_2 _21872_ (.A(_18882_),
    .B(_02417_),
    .X(_03810_));
 sky130_fd_sc_hd__buf_1 _21873_ (.A(_18880_),
    .X(_18883_));
 sky130_fd_sc_hd__and2_2 _21874_ (.A(_18883_),
    .B(_02416_),
    .X(_03809_));
 sky130_fd_sc_hd__and2_2 _21875_ (.A(_18883_),
    .B(_02415_),
    .X(_03808_));
 sky130_fd_sc_hd__and2_2 _21876_ (.A(_18883_),
    .B(_02414_),
    .X(_03807_));
 sky130_fd_sc_hd__and2_2 _21877_ (.A(_18883_),
    .B(_02413_),
    .X(_03806_));
 sky130_fd_sc_hd__and2_2 _21878_ (.A(_18883_),
    .B(_02412_),
    .X(_03805_));
 sky130_fd_sc_hd__and2_2 _21879_ (.A(_18883_),
    .B(_02442_),
    .X(_03804_));
 sky130_fd_sc_hd__buf_1 _21880_ (.A(_18880_),
    .X(_18884_));
 sky130_fd_sc_hd__and2_2 _21881_ (.A(_18884_),
    .B(_02441_),
    .X(_03803_));
 sky130_fd_sc_hd__and2_2 _21882_ (.A(_18884_),
    .B(_02440_),
    .X(_03802_));
 sky130_fd_sc_hd__and2_2 _21883_ (.A(_18884_),
    .B(_02439_),
    .X(_03801_));
 sky130_fd_sc_hd__and2_2 _21884_ (.A(_18884_),
    .B(_02438_),
    .X(_03800_));
 sky130_fd_sc_hd__and2_2 _21885_ (.A(_18884_),
    .B(_02437_),
    .X(_03799_));
 sky130_fd_sc_hd__and2_2 _21886_ (.A(_18884_),
    .B(_02436_),
    .X(_03798_));
 sky130_fd_sc_hd__buf_1 _21887_ (.A(_18880_),
    .X(_18885_));
 sky130_fd_sc_hd__and2_2 _21888_ (.A(_18885_),
    .B(_02433_),
    .X(_03797_));
 sky130_fd_sc_hd__and2_2 _21889_ (.A(_18885_),
    .B(_02422_),
    .X(_03796_));
 sky130_fd_sc_hd__and2_2 _21890_ (.A(_18885_),
    .B(_02411_),
    .X(_03795_));
 sky130_fd_sc_hd__nand2_2 _21891_ (.A(\count_cycle[56] ),
    .B(\count_cycle[57] ),
    .Y(_18886_));
 sky130_fd_sc_hd__inv_2 _21892_ (.A(\count_cycle[58] ),
    .Y(_18887_));
 sky130_fd_sc_hd__inv_2 _21893_ (.A(\count_cycle[59] ),
    .Y(_18888_));
 sky130_fd_sc_hd__inv_2 _21894_ (.A(\count_cycle[62] ),
    .Y(_18889_));
 sky130_fd_sc_hd__inv_2 _21895_ (.A(\count_cycle[60] ),
    .Y(_18890_));
 sky130_fd_sc_hd__inv_2 _21896_ (.A(\count_cycle[61] ),
    .Y(_18891_));
 sky130_fd_sc_hd__nor2_2 _21897_ (.A(_18890_),
    .B(_18891_),
    .Y(_18892_));
 sky130_fd_sc_hd__or4b_2 _21898_ (.A(_18887_),
    .B(_18888_),
    .C(_18889_),
    .D_N(_18892_),
    .X(_18893_));
 sky130_fd_sc_hd__and3_2 _21899_ (.A(\count_cycle[41] ),
    .B(\count_cycle[42] ),
    .C(\count_cycle[43] ),
    .X(_18894_));
 sky130_fd_sc_hd__inv_2 _21900_ (.A(_18894_),
    .Y(_18895_));
 sky130_fd_sc_hd__and3_2 _21901_ (.A(\count_cycle[28] ),
    .B(\count_cycle[29] ),
    .C(\count_cycle[30] ),
    .X(_18896_));
 sky130_fd_sc_hd__and3_2 _21902_ (.A(_18896_),
    .B(\count_cycle[27] ),
    .C(\count_cycle[31] ),
    .X(_18897_));
 sky130_fd_sc_hd__inv_2 _21903_ (.A(_18897_),
    .Y(_18898_));
 sky130_fd_sc_hd__inv_2 _21904_ (.A(\count_cycle[21] ),
    .Y(_01965_));
 sky130_fd_sc_hd__inv_2 _21905_ (.A(\count_cycle[22] ),
    .Y(_01974_));
 sky130_fd_sc_hd__inv_2 _21906_ (.A(\count_cycle[23] ),
    .Y(_01983_));
 sky130_fd_sc_hd__inv_2 _21907_ (.A(\count_cycle[24] ),
    .Y(_01992_));
 sky130_fd_sc_hd__or4_2 _21908_ (.A(_01965_),
    .B(_01974_),
    .C(_01983_),
    .D(_01992_),
    .X(_18899_));
 sky130_fd_sc_hd__inv_2 _21909_ (.A(\count_cycle[20] ),
    .Y(_01956_));
 sky130_fd_sc_hd__inv_2 _21910_ (.A(\count_cycle[18] ),
    .Y(_01938_));
 sky130_fd_sc_hd__inv_2 _21911_ (.A(\count_cycle[16] ),
    .Y(_01920_));
 sky130_fd_sc_hd__inv_2 _21912_ (.A(\count_cycle[15] ),
    .Y(_01911_));
 sky130_fd_sc_hd__inv_2 _21913_ (.A(\count_cycle[13] ),
    .Y(_01885_));
 sky130_fd_sc_hd__inv_2 _21914_ (.A(\count_cycle[12] ),
    .Y(_01872_));
 sky130_fd_sc_hd__inv_2 _21915_ (.A(\count_cycle[10] ),
    .Y(_01846_));
 sky130_fd_sc_hd__inv_2 _21916_ (.A(\count_cycle[9] ),
    .Y(_01833_));
 sky130_fd_sc_hd__inv_2 _21917_ (.A(\count_cycle[7] ),
    .Y(_01806_));
 sky130_fd_sc_hd__inv_2 _21918_ (.A(\count_cycle[8] ),
    .Y(_01820_));
 sky130_fd_sc_hd__inv_2 _21919_ (.A(\count_cycle[5] ),
    .Y(_01780_));
 sky130_fd_sc_hd__inv_2 _21920_ (.A(\count_cycle[3] ),
    .Y(_01754_));
 sky130_fd_sc_hd__nand2_2 _21921_ (.A(\count_cycle[0] ),
    .B(\count_cycle[1] ),
    .Y(_18900_));
 sky130_fd_sc_hd__inv_2 _21922_ (.A(\count_cycle[2] ),
    .Y(_01741_));
 sky130_fd_sc_hd__or2_2 _21923_ (.A(_18900_),
    .B(_01741_),
    .X(_18901_));
 sky130_fd_sc_hd__nor2_2 _21924_ (.A(_01754_),
    .B(_18901_),
    .Y(_18902_));
 sky130_fd_sc_hd__nand2_2 _21925_ (.A(_18902_),
    .B(\count_cycle[4] ),
    .Y(_18903_));
 sky130_fd_sc_hd__nor2_2 _21926_ (.A(_01780_),
    .B(_18903_),
    .Y(_18904_));
 sky130_fd_sc_hd__nand2_2 _21927_ (.A(_18904_),
    .B(\count_cycle[6] ),
    .Y(_18905_));
 sky130_fd_sc_hd__or3_2 _21928_ (.A(_01806_),
    .B(_01820_),
    .C(_18905_),
    .X(_18906_));
 sky130_fd_sc_hd__or2_2 _21929_ (.A(_01833_),
    .B(_18906_),
    .X(_18907_));
 sky130_fd_sc_hd__nor2_2 _21930_ (.A(_01846_),
    .B(_18907_),
    .Y(_18908_));
 sky130_fd_sc_hd__nand2_2 _21931_ (.A(_18908_),
    .B(\count_cycle[11] ),
    .Y(_18909_));
 sky130_fd_sc_hd__or2_2 _21932_ (.A(_01872_),
    .B(_18909_),
    .X(_18910_));
 sky130_fd_sc_hd__nor2_2 _21933_ (.A(_01885_),
    .B(_18910_),
    .Y(_18911_));
 sky130_fd_sc_hd__nand2_2 _21934_ (.A(_18911_),
    .B(\count_cycle[14] ),
    .Y(_18912_));
 sky130_fd_sc_hd__or2_2 _21935_ (.A(_01911_),
    .B(_18912_),
    .X(_18913_));
 sky130_fd_sc_hd__nor2_2 _21936_ (.A(_01920_),
    .B(_18913_),
    .Y(_18914_));
 sky130_fd_sc_hd__nand2_2 _21937_ (.A(_18914_),
    .B(\count_cycle[17] ),
    .Y(_18915_));
 sky130_fd_sc_hd__nor2_2 _21938_ (.A(_01938_),
    .B(_18915_),
    .Y(_18916_));
 sky130_fd_sc_hd__nand2_2 _21939_ (.A(_18916_),
    .B(\count_cycle[19] ),
    .Y(_18917_));
 sky130_fd_sc_hd__or2_2 _21940_ (.A(_01956_),
    .B(_18917_),
    .X(_18918_));
 sky130_fd_sc_hd__nor2_2 _21941_ (.A(_18899_),
    .B(_18918_),
    .Y(_18919_));
 sky130_fd_sc_hd__inv_2 _21942_ (.A(\count_cycle[25] ),
    .Y(_02001_));
 sky130_fd_sc_hd__inv_2 _21943_ (.A(\count_cycle[26] ),
    .Y(_02010_));
 sky130_fd_sc_hd__nor2_2 _21944_ (.A(_02001_),
    .B(_02010_),
    .Y(_18920_));
 sky130_fd_sc_hd__nand2_2 _21945_ (.A(_18919_),
    .B(_18920_),
    .Y(_18921_));
 sky130_fd_sc_hd__nor2_2 _21946_ (.A(_18898_),
    .B(_18921_),
    .Y(_18922_));
 sky130_fd_sc_hd__and3_2 _21947_ (.A(_18922_),
    .B(\count_cycle[32] ),
    .C(\count_cycle[33] ),
    .X(_18923_));
 sky130_fd_sc_hd__and3_2 _21948_ (.A(\count_cycle[34] ),
    .B(\count_cycle[35] ),
    .C(\count_cycle[36] ),
    .X(_18924_));
 sky130_fd_sc_hd__and4_2 _21949_ (.A(\count_cycle[37] ),
    .B(\count_cycle[38] ),
    .C(\count_cycle[39] ),
    .D(\count_cycle[40] ),
    .X(_18925_));
 sky130_fd_sc_hd__nand3_2 _21950_ (.A(_18923_),
    .B(_18924_),
    .C(_18925_),
    .Y(_18926_));
 sky130_fd_sc_hd__nor2_2 _21951_ (.A(_18895_),
    .B(_18926_),
    .Y(_18927_));
 sky130_fd_sc_hd__and3_2 _21952_ (.A(\count_cycle[44] ),
    .B(\count_cycle[45] ),
    .C(\count_cycle[46] ),
    .X(_18928_));
 sky130_fd_sc_hd__and4_2 _21953_ (.A(_18928_),
    .B(\count_cycle[47] ),
    .C(\count_cycle[48] ),
    .D(\count_cycle[49] ),
    .X(_18929_));
 sky130_fd_sc_hd__nand2_2 _21954_ (.A(\count_cycle[50] ),
    .B(\count_cycle[51] ),
    .Y(_18930_));
 sky130_fd_sc_hd__inv_2 _21955_ (.A(\count_cycle[52] ),
    .Y(_18931_));
 sky130_fd_sc_hd__nor2_2 _21956_ (.A(_18930_),
    .B(_18931_),
    .Y(_18932_));
 sky130_fd_sc_hd__and4_2 _21957_ (.A(_18927_),
    .B(\count_cycle[53] ),
    .C(_18929_),
    .D(_18932_),
    .X(_18933_));
 sky130_fd_sc_hd__and2_2 _21958_ (.A(\count_cycle[54] ),
    .B(\count_cycle[55] ),
    .X(_18934_));
 sky130_fd_sc_hd__nand2_2 _21959_ (.A(_18933_),
    .B(_18934_),
    .Y(_18935_));
 sky130_fd_sc_hd__inv_2 _21960_ (.A(\count_cycle[63] ),
    .Y(_18936_));
 sky130_fd_sc_hd__o31a_2 _21961_ (.A1(_18886_),
    .A2(_18893_),
    .A3(_18935_),
    .B1(_18936_),
    .X(_18937_));
 sky130_fd_sc_hd__o41ai_2 _21962_ (.A1(_18936_),
    .A2(_18886_),
    .A3(_18893_),
    .A4(_18935_),
    .B1(_18638_),
    .Y(_18938_));
 sky130_fd_sc_hd__nor2_2 _21963_ (.A(_18937_),
    .B(_18938_),
    .Y(_03794_));
 sky130_fd_sc_hd__nand2_2 _21964_ (.A(\count_cycle[57] ),
    .B(\count_cycle[58] ),
    .Y(_18939_));
 sky130_fd_sc_hd__nor2_2 _21965_ (.A(_18939_),
    .B(_18888_),
    .Y(_18940_));
 sky130_fd_sc_hd__inv_2 _21966_ (.A(_18940_),
    .Y(_18941_));
 sky130_fd_sc_hd__and3_2 _21967_ (.A(\count_cycle[54] ),
    .B(\count_cycle[55] ),
    .C(\count_cycle[56] ),
    .X(_18942_));
 sky130_fd_sc_hd__nand2_2 _21968_ (.A(_18933_),
    .B(_18942_),
    .Y(_18943_));
 sky130_fd_sc_hd__nor2_2 _21969_ (.A(_18941_),
    .B(_18943_),
    .Y(_18944_));
 sky130_fd_sc_hd__nand2_2 _21970_ (.A(_18944_),
    .B(_18892_),
    .Y(_18945_));
 sky130_fd_sc_hd__o31ai_2 _21971_ (.A1(_18886_),
    .A2(_18893_),
    .A3(_18935_),
    .B1(_18638_),
    .Y(_18946_));
 sky130_fd_sc_hd__a21oi_2 _21972_ (.A1(_18945_),
    .A2(_18889_),
    .B1(_18946_),
    .Y(_03793_));
 sky130_fd_sc_hd__nand2_2 _21973_ (.A(_18944_),
    .B(\count_cycle[60] ),
    .Y(_18947_));
 sky130_fd_sc_hd__buf_1 _21974_ (.A(_18933_),
    .X(_18948_));
 sky130_fd_sc_hd__a41o_2 _21975_ (.A1(_18948_),
    .A2(_18892_),
    .A3(_18942_),
    .A4(_18940_),
    .B1(_18189_),
    .X(_18949_));
 sky130_fd_sc_hd__a21oi_2 _21976_ (.A1(_18947_),
    .A2(_18891_),
    .B1(_18949_),
    .Y(_03792_));
 sky130_fd_sc_hd__buf_1 _21977_ (.A(_18943_),
    .X(_18950_));
 sky130_fd_sc_hd__o31a_2 _21978_ (.A1(_18890_),
    .A2(_18941_),
    .A3(_18950_),
    .B1(_18880_),
    .X(_18951_));
 sky130_fd_sc_hd__o21a_2 _21979_ (.A1(\count_cycle[60] ),
    .A2(_18944_),
    .B1(_18951_),
    .X(_03791_));
 sky130_fd_sc_hd__o21ai_2 _21980_ (.A1(_18939_),
    .A2(_18950_),
    .B1(_18888_),
    .Y(_18952_));
 sky130_fd_sc_hd__o211a_2 _21981_ (.A1(_18950_),
    .A2(_18941_),
    .B1(_18849_),
    .C1(_18952_),
    .X(_03790_));
 sky130_fd_sc_hd__a31o_2 _21982_ (.A1(_18933_),
    .A2(\count_cycle[57] ),
    .A3(_18942_),
    .B1(\count_cycle[58] ),
    .X(_18953_));
 sky130_fd_sc_hd__o211a_2 _21983_ (.A1(_18950_),
    .A2(_18939_),
    .B1(_18849_),
    .C1(_18953_),
    .X(_03789_));
 sky130_fd_sc_hd__inv_2 _21984_ (.A(\count_cycle[57] ),
    .Y(_18954_));
 sky130_fd_sc_hd__a31o_2 _21985_ (.A1(_18948_),
    .A2(\count_cycle[57] ),
    .A3(_18942_),
    .B1(_18238_),
    .X(_18955_));
 sky130_fd_sc_hd__a21oi_2 _21986_ (.A1(_18954_),
    .A2(_18950_),
    .B1(_18955_),
    .Y(_03788_));
 sky130_fd_sc_hd__a21o_2 _21987_ (.A1(_18948_),
    .A2(_18934_),
    .B1(\count_cycle[56] ),
    .X(_18956_));
 sky130_fd_sc_hd__and3_2 _21988_ (.A(_18956_),
    .B(_18791_),
    .C(_18950_),
    .X(_03787_));
 sky130_fd_sc_hd__a21o_2 _21989_ (.A1(_18933_),
    .A2(\count_cycle[54] ),
    .B1(\count_cycle[55] ),
    .X(_18957_));
 sky130_fd_sc_hd__buf_1 _21990_ (.A(_18778_),
    .X(_18958_));
 sky130_fd_sc_hd__and3_2 _21991_ (.A(_18957_),
    .B(_18958_),
    .C(_18935_),
    .X(_03786_));
 sky130_fd_sc_hd__o21ai_2 _21992_ (.A1(\count_cycle[54] ),
    .A2(_18948_),
    .B1(_18638_),
    .Y(_18959_));
 sky130_fd_sc_hd__a21oi_2 _21993_ (.A1(\count_cycle[54] ),
    .A2(_18948_),
    .B1(_18959_),
    .Y(_03785_));
 sky130_fd_sc_hd__buf_1 _21994_ (.A(_18927_),
    .X(_18960_));
 sky130_fd_sc_hd__nand2_2 _21995_ (.A(_18960_),
    .B(_18929_),
    .Y(_18961_));
 sky130_fd_sc_hd__or2_2 _21996_ (.A(_18930_),
    .B(_18961_),
    .X(_18962_));
 sky130_fd_sc_hd__nor2_2 _21997_ (.A(_18931_),
    .B(_18962_),
    .Y(_18963_));
 sky130_fd_sc_hd__nor2_2 _21998_ (.A(_18331_),
    .B(_18948_),
    .Y(_18964_));
 sky130_fd_sc_hd__o21a_2 _21999_ (.A1(\count_cycle[53] ),
    .A2(_18963_),
    .B1(_18964_),
    .X(_03784_));
 sky130_fd_sc_hd__inv_2 _22000_ (.A(\count_cycle[50] ),
    .Y(_18965_));
 sky130_fd_sc_hd__nand2_2 _22001_ (.A(\count_cycle[51] ),
    .B(\count_cycle[52] ),
    .Y(_18966_));
 sky130_fd_sc_hd__nand2_2 _22002_ (.A(_18962_),
    .B(_18931_),
    .Y(_18967_));
 sky130_fd_sc_hd__o311a_2 _22003_ (.A1(_18965_),
    .A2(_18961_),
    .A3(_18966_),
    .B1(_18407_),
    .C1(_18967_),
    .X(_03783_));
 sky130_fd_sc_hd__a31o_2 _22004_ (.A1(_18960_),
    .A2(\count_cycle[50] ),
    .A3(_18929_),
    .B1(\count_cycle[51] ),
    .X(_18968_));
 sky130_fd_sc_hd__and3_2 _22005_ (.A(_18962_),
    .B(_18958_),
    .C(_18968_),
    .X(_03782_));
 sky130_fd_sc_hd__a31o_2 _22006_ (.A1(_18960_),
    .A2(\count_cycle[50] ),
    .A3(_18929_),
    .B1(_18189_),
    .X(_18969_));
 sky130_fd_sc_hd__a21oi_2 _22007_ (.A1(_18965_),
    .A2(_18961_),
    .B1(_18969_),
    .Y(_03781_));
 sky130_fd_sc_hd__inv_2 _22008_ (.A(\count_cycle[47] ),
    .Y(_18970_));
 sky130_fd_sc_hd__nand2_2 _22009_ (.A(_18960_),
    .B(_18928_),
    .Y(_18971_));
 sky130_fd_sc_hd__nor2_2 _22010_ (.A(_18970_),
    .B(_18971_),
    .Y(_18972_));
 sky130_fd_sc_hd__nand2_2 _22011_ (.A(_18972_),
    .B(\count_cycle[48] ),
    .Y(_18973_));
 sky130_fd_sc_hd__inv_2 _22012_ (.A(\count_cycle[49] ),
    .Y(_18974_));
 sky130_fd_sc_hd__nand2_2 _22013_ (.A(_18973_),
    .B(_18974_),
    .Y(_18975_));
 sky130_fd_sc_hd__and3_2 _22014_ (.A(_18975_),
    .B(_18958_),
    .C(_18961_),
    .X(_03780_));
 sky130_fd_sc_hd__or2_2 _22015_ (.A(\count_cycle[48] ),
    .B(_18972_),
    .X(_18976_));
 sky130_fd_sc_hd__and3_2 _22016_ (.A(_18976_),
    .B(_18958_),
    .C(_18973_),
    .X(_03779_));
 sky130_fd_sc_hd__a21o_2 _22017_ (.A1(_18971_),
    .A2(_18970_),
    .B1(_18349_),
    .X(_18977_));
 sky130_fd_sc_hd__nor2_2 _22018_ (.A(_18972_),
    .B(_18977_),
    .Y(_03778_));
 sky130_fd_sc_hd__inv_2 _22019_ (.A(\count_cycle[45] ),
    .Y(_18978_));
 sky130_fd_sc_hd__nand2_2 _22020_ (.A(_18960_),
    .B(\count_cycle[44] ),
    .Y(_18979_));
 sky130_fd_sc_hd__or2_2 _22021_ (.A(_18978_),
    .B(_18979_),
    .X(_18980_));
 sky130_fd_sc_hd__inv_2 _22022_ (.A(\count_cycle[46] ),
    .Y(_18981_));
 sky130_fd_sc_hd__nand2_2 _22023_ (.A(_18980_),
    .B(_18981_),
    .Y(_18982_));
 sky130_fd_sc_hd__and3_2 _22024_ (.A(_18982_),
    .B(_18971_),
    .C(_18660_),
    .X(_03777_));
 sky130_fd_sc_hd__nand2_2 _22025_ (.A(_18979_),
    .B(_18978_),
    .Y(_18983_));
 sky130_fd_sc_hd__and3_2 _22026_ (.A(_18980_),
    .B(_18958_),
    .C(_18983_),
    .X(_03776_));
 sky130_fd_sc_hd__or2_2 _22027_ (.A(\count_cycle[44] ),
    .B(_18960_),
    .X(_18984_));
 sky130_fd_sc_hd__and3_2 _22028_ (.A(_18984_),
    .B(_18958_),
    .C(_18979_),
    .X(_03775_));
 sky130_fd_sc_hd__inv_2 _22029_ (.A(_18926_),
    .Y(_18985_));
 sky130_fd_sc_hd__buf_1 _22030_ (.A(\count_cycle[41] ),
    .X(_18986_));
 sky130_fd_sc_hd__a31o_2 _22031_ (.A1(_18985_),
    .A2(_18986_),
    .A3(\count_cycle[42] ),
    .B1(\count_cycle[43] ),
    .X(_18987_));
 sky130_fd_sc_hd__o211a_2 _22032_ (.A1(_18926_),
    .A2(_18895_),
    .B1(_18660_),
    .C1(_18987_),
    .X(_03774_));
 sky130_fd_sc_hd__a21oi_2 _22033_ (.A1(_18985_),
    .A2(_18986_),
    .B1(\count_cycle[42] ),
    .Y(_18988_));
 sky130_fd_sc_hd__a31o_2 _22034_ (.A1(_18985_),
    .A2(_18986_),
    .A3(\count_cycle[42] ),
    .B1(_18238_),
    .X(_18989_));
 sky130_fd_sc_hd__nor2_2 _22035_ (.A(_18988_),
    .B(_18989_),
    .Y(_03773_));
 sky130_fd_sc_hd__a21oi_2 _22036_ (.A1(_18985_),
    .A2(_18986_),
    .B1(_18349_),
    .Y(_18990_));
 sky130_fd_sc_hd__o21a_2 _22037_ (.A1(_18986_),
    .A2(_18985_),
    .B1(_18990_),
    .X(_03772_));
 sky130_fd_sc_hd__inv_2 _22038_ (.A(\count_cycle[38] ),
    .Y(_18991_));
 sky130_fd_sc_hd__inv_2 _22039_ (.A(\count_cycle[39] ),
    .Y(_18992_));
 sky130_fd_sc_hd__inv_2 _22040_ (.A(_18924_),
    .Y(_18993_));
 sky130_fd_sc_hd__inv_2 _22041_ (.A(_18923_),
    .Y(_18994_));
 sky130_fd_sc_hd__nor2_2 _22042_ (.A(_18993_),
    .B(_18994_),
    .Y(_18995_));
 sky130_fd_sc_hd__nand2_2 _22043_ (.A(_18995_),
    .B(\count_cycle[37] ),
    .Y(_18996_));
 sky130_fd_sc_hd__or3_2 _22044_ (.A(_18991_),
    .B(_18992_),
    .C(_18996_),
    .X(_18997_));
 sky130_fd_sc_hd__inv_2 _22045_ (.A(\count_cycle[40] ),
    .Y(_18998_));
 sky130_fd_sc_hd__nand2_2 _22046_ (.A(_18997_),
    .B(_18998_),
    .Y(_18999_));
 sky130_fd_sc_hd__buf_1 _22047_ (.A(_18778_),
    .X(_19000_));
 sky130_fd_sc_hd__and3_2 _22048_ (.A(_18999_),
    .B(_19000_),
    .C(_18926_),
    .X(_03771_));
 sky130_fd_sc_hd__or2_2 _22049_ (.A(_18991_),
    .B(_18996_),
    .X(_19001_));
 sky130_fd_sc_hd__nand2_2 _22050_ (.A(_19001_),
    .B(_18992_),
    .Y(_19002_));
 sky130_fd_sc_hd__and3_2 _22051_ (.A(_19002_),
    .B(_18997_),
    .C(_18660_),
    .X(_03770_));
 sky130_fd_sc_hd__nand2_2 _22052_ (.A(_18996_),
    .B(_18991_),
    .Y(_19003_));
 sky130_fd_sc_hd__and3_2 _22053_ (.A(_19001_),
    .B(_19000_),
    .C(_19003_),
    .X(_03769_));
 sky130_fd_sc_hd__or2_2 _22054_ (.A(\count_cycle[37] ),
    .B(_18995_),
    .X(_19004_));
 sky130_fd_sc_hd__and3_2 _22055_ (.A(_19004_),
    .B(_19000_),
    .C(_18996_),
    .X(_03768_));
 sky130_fd_sc_hd__inv_2 _22056_ (.A(\count_cycle[36] ),
    .Y(_19005_));
 sky130_fd_sc_hd__inv_2 _22057_ (.A(\count_cycle[35] ),
    .Y(_19006_));
 sky130_fd_sc_hd__nand2_2 _22058_ (.A(_18923_),
    .B(\count_cycle[34] ),
    .Y(_19007_));
 sky130_fd_sc_hd__or2_2 _22059_ (.A(_19006_),
    .B(_19007_),
    .X(_19008_));
 sky130_fd_sc_hd__or2_2 _22060_ (.A(_18721_),
    .B(_18995_),
    .X(_19009_));
 sky130_fd_sc_hd__a21oi_2 _22061_ (.A1(_19005_),
    .A2(_19008_),
    .B1(_19009_),
    .Y(_03767_));
 sky130_fd_sc_hd__nand2_2 _22062_ (.A(_19007_),
    .B(_19006_),
    .Y(_19010_));
 sky130_fd_sc_hd__and3_2 _22063_ (.A(_19008_),
    .B(_19000_),
    .C(_19010_),
    .X(_03766_));
 sky130_fd_sc_hd__or2_2 _22064_ (.A(\count_cycle[34] ),
    .B(_18923_),
    .X(_19011_));
 sky130_fd_sc_hd__and3_2 _22065_ (.A(_19011_),
    .B(_19000_),
    .C(_19007_),
    .X(_03765_));
 sky130_fd_sc_hd__inv_2 _22066_ (.A(\count_cycle[32] ),
    .Y(_19012_));
 sky130_fd_sc_hd__inv_2 _22067_ (.A(_18922_),
    .Y(_19013_));
 sky130_fd_sc_hd__nor2_2 _22068_ (.A(_19012_),
    .B(_19013_),
    .Y(_19014_));
 sky130_fd_sc_hd__inv_2 _22069_ (.A(_19014_),
    .Y(_19015_));
 sky130_fd_sc_hd__inv_2 _22070_ (.A(\count_cycle[33] ),
    .Y(_19016_));
 sky130_fd_sc_hd__nand2_2 _22071_ (.A(_19015_),
    .B(_19016_),
    .Y(_19017_));
 sky130_fd_sc_hd__and3_2 _22072_ (.A(_19017_),
    .B(_19000_),
    .C(_18994_),
    .X(_03764_));
 sky130_fd_sc_hd__buf_1 _22073_ (.A(_18778_),
    .X(_19018_));
 sky130_fd_sc_hd__nand2_2 _22074_ (.A(_19013_),
    .B(_19012_),
    .Y(_19019_));
 sky130_fd_sc_hd__and3_2 _22075_ (.A(_19015_),
    .B(_19018_),
    .C(_19019_),
    .X(_03763_));
 sky130_fd_sc_hd__inv_2 _22076_ (.A(\count_cycle[30] ),
    .Y(_02046_));
 sky130_fd_sc_hd__inv_2 _22077_ (.A(\count_cycle[29] ),
    .Y(_02037_));
 sky130_fd_sc_hd__inv_2 _22078_ (.A(\count_cycle[28] ),
    .Y(_02028_));
 sky130_fd_sc_hd__inv_2 _22079_ (.A(\count_cycle[27] ),
    .Y(_02019_));
 sky130_fd_sc_hd__or2_2 _22080_ (.A(_02019_),
    .B(_18921_),
    .X(_19020_));
 sky130_fd_sc_hd__or2_2 _22081_ (.A(_02028_),
    .B(_19020_),
    .X(_19021_));
 sky130_fd_sc_hd__or2_2 _22082_ (.A(_02037_),
    .B(_19021_),
    .X(_19022_));
 sky130_fd_sc_hd__nor2_2 _22083_ (.A(_02046_),
    .B(_19022_),
    .Y(_19023_));
 sky130_fd_sc_hd__or2_2 _22084_ (.A(\count_cycle[31] ),
    .B(_19023_),
    .X(_19024_));
 sky130_fd_sc_hd__and3_2 _22085_ (.A(_19024_),
    .B(_19018_),
    .C(_19013_),
    .X(_03762_));
 sky130_fd_sc_hd__a21o_2 _22086_ (.A1(_19022_),
    .A2(_02046_),
    .B1(_18349_),
    .X(_19025_));
 sky130_fd_sc_hd__nor2_2 _22087_ (.A(_19023_),
    .B(_19025_),
    .Y(_03761_));
 sky130_fd_sc_hd__nand2_2 _22088_ (.A(_19021_),
    .B(_02037_),
    .Y(_19026_));
 sky130_fd_sc_hd__and3_2 _22089_ (.A(_19022_),
    .B(_19018_),
    .C(_19026_),
    .X(_03760_));
 sky130_fd_sc_hd__nand2_2 _22090_ (.A(_19020_),
    .B(_02028_),
    .Y(_19027_));
 sky130_fd_sc_hd__and3_2 _22091_ (.A(_19021_),
    .B(_19018_),
    .C(_19027_),
    .X(_03759_));
 sky130_fd_sc_hd__nand2_2 _22092_ (.A(_18921_),
    .B(_02019_),
    .Y(_19028_));
 sky130_fd_sc_hd__and3_2 _22093_ (.A(_19020_),
    .B(_19018_),
    .C(_19028_),
    .X(_03758_));
 sky130_fd_sc_hd__nand2_2 _22094_ (.A(_18919_),
    .B(\count_cycle[25] ),
    .Y(_19029_));
 sky130_fd_sc_hd__nand2_2 _22095_ (.A(_19029_),
    .B(_02010_),
    .Y(_19030_));
 sky130_fd_sc_hd__and3_2 _22096_ (.A(_19030_),
    .B(_19018_),
    .C(_18921_),
    .X(_03757_));
 sky130_fd_sc_hd__or2_2 _22097_ (.A(\count_cycle[25] ),
    .B(_18919_),
    .X(_19031_));
 sky130_fd_sc_hd__buf_1 _22098_ (.A(_18778_),
    .X(_19032_));
 sky130_fd_sc_hd__and3_2 _22099_ (.A(_19031_),
    .B(_19032_),
    .C(_19029_),
    .X(_03756_));
 sky130_fd_sc_hd__or2_2 _22100_ (.A(_01965_),
    .B(_18918_),
    .X(_19033_));
 sky130_fd_sc_hd__nor2_2 _22101_ (.A(_01974_),
    .B(_19033_),
    .Y(_19034_));
 sky130_fd_sc_hd__nand2_2 _22102_ (.A(_19034_),
    .B(\count_cycle[23] ),
    .Y(_19035_));
 sky130_fd_sc_hd__or2_2 _22103_ (.A(_18278_),
    .B(_18919_),
    .X(_19036_));
 sky130_fd_sc_hd__a21oi_2 _22104_ (.A1(_19035_),
    .A2(_01992_),
    .B1(_19036_),
    .Y(_03755_));
 sky130_fd_sc_hd__inv_2 _22105_ (.A(_19034_),
    .Y(_19037_));
 sky130_fd_sc_hd__nand2_2 _22106_ (.A(_19037_),
    .B(_01983_),
    .Y(_19038_));
 sky130_fd_sc_hd__and3_2 _22107_ (.A(_19038_),
    .B(_19032_),
    .C(_19035_),
    .X(_03754_));
 sky130_fd_sc_hd__nand2_2 _22108_ (.A(_19033_),
    .B(_01974_),
    .Y(_19039_));
 sky130_fd_sc_hd__and3_2 _22109_ (.A(_19037_),
    .B(_19032_),
    .C(_19039_),
    .X(_03753_));
 sky130_fd_sc_hd__nand2_2 _22110_ (.A(_18918_),
    .B(_01965_),
    .Y(_19040_));
 sky130_fd_sc_hd__and3_2 _22111_ (.A(_19033_),
    .B(_19032_),
    .C(_19040_),
    .X(_03752_));
 sky130_fd_sc_hd__nand2_2 _22112_ (.A(_18917_),
    .B(_01956_),
    .Y(_19041_));
 sky130_fd_sc_hd__and3_2 _22113_ (.A(_18918_),
    .B(_19032_),
    .C(_19041_),
    .X(_03751_));
 sky130_fd_sc_hd__or2_2 _22114_ (.A(\count_cycle[19] ),
    .B(_18916_),
    .X(_19042_));
 sky130_fd_sc_hd__and3_2 _22115_ (.A(_19042_),
    .B(_19032_),
    .C(_18917_),
    .X(_03750_));
 sky130_fd_sc_hd__or2_2 _22116_ (.A(_18278_),
    .B(_18916_),
    .X(_19043_));
 sky130_fd_sc_hd__a21oi_2 _22117_ (.A1(_01938_),
    .A2(_18915_),
    .B1(_19043_),
    .Y(_03749_));
 sky130_fd_sc_hd__inv_2 _22118_ (.A(_18914_),
    .Y(_19044_));
 sky130_fd_sc_hd__inv_2 _22119_ (.A(\count_cycle[17] ),
    .Y(_01929_));
 sky130_fd_sc_hd__nand2_2 _22120_ (.A(_19044_),
    .B(_01929_),
    .Y(_19045_));
 sky130_fd_sc_hd__buf_1 _22121_ (.A(_18637_),
    .X(_19046_));
 sky130_fd_sc_hd__and3_2 _22122_ (.A(_19045_),
    .B(_19046_),
    .C(_18915_),
    .X(_03748_));
 sky130_fd_sc_hd__nand2_2 _22123_ (.A(_18913_),
    .B(_01920_),
    .Y(_19047_));
 sky130_fd_sc_hd__and3_2 _22124_ (.A(_19044_),
    .B(_19046_),
    .C(_19047_),
    .X(_03747_));
 sky130_fd_sc_hd__nand2_2 _22125_ (.A(_18912_),
    .B(_01911_),
    .Y(_19048_));
 sky130_fd_sc_hd__and3_2 _22126_ (.A(_18913_),
    .B(_19046_),
    .C(_19048_),
    .X(_03746_));
 sky130_fd_sc_hd__or2_2 _22127_ (.A(\count_cycle[14] ),
    .B(_18911_),
    .X(_19049_));
 sky130_fd_sc_hd__and3_2 _22128_ (.A(_19049_),
    .B(_19046_),
    .C(_18912_),
    .X(_03745_));
 sky130_fd_sc_hd__or2_2 _22129_ (.A(_18278_),
    .B(_18911_),
    .X(_19050_));
 sky130_fd_sc_hd__a21oi_2 _22130_ (.A1(_01885_),
    .A2(_18910_),
    .B1(_19050_),
    .Y(_03744_));
 sky130_fd_sc_hd__nand2_2 _22131_ (.A(_18909_),
    .B(_01872_),
    .Y(_19051_));
 sky130_fd_sc_hd__and3_2 _22132_ (.A(_18910_),
    .B(_19046_),
    .C(_19051_),
    .X(_03743_));
 sky130_fd_sc_hd__inv_2 _22133_ (.A(_18908_),
    .Y(_19052_));
 sky130_fd_sc_hd__inv_2 _22134_ (.A(\count_cycle[11] ),
    .Y(_01859_));
 sky130_fd_sc_hd__nand2_2 _22135_ (.A(_19052_),
    .B(_01859_),
    .Y(_19053_));
 sky130_fd_sc_hd__and3_2 _22136_ (.A(_19053_),
    .B(_19046_),
    .C(_18909_),
    .X(_03742_));
 sky130_fd_sc_hd__buf_1 _22137_ (.A(_18637_),
    .X(_19054_));
 sky130_fd_sc_hd__nand2_2 _22138_ (.A(_18907_),
    .B(_01846_),
    .Y(_19055_));
 sky130_fd_sc_hd__and3_2 _22139_ (.A(_19052_),
    .B(_19054_),
    .C(_19055_),
    .X(_03741_));
 sky130_fd_sc_hd__nand2_2 _22140_ (.A(_18906_),
    .B(_01833_),
    .Y(_19056_));
 sky130_fd_sc_hd__and3_2 _22141_ (.A(_18907_),
    .B(_19054_),
    .C(_19056_),
    .X(_03740_));
 sky130_fd_sc_hd__or2_2 _22142_ (.A(_01806_),
    .B(_18905_),
    .X(_19057_));
 sky130_fd_sc_hd__nand2_2 _22143_ (.A(_19057_),
    .B(_01820_),
    .Y(_19058_));
 sky130_fd_sc_hd__and3_2 _22144_ (.A(_19058_),
    .B(_18906_),
    .C(_18660_),
    .X(_03739_));
 sky130_fd_sc_hd__nand2_2 _22145_ (.A(_18905_),
    .B(_01806_),
    .Y(_19059_));
 sky130_fd_sc_hd__and3_2 _22146_ (.A(_19057_),
    .B(_19054_),
    .C(_19059_),
    .X(_03738_));
 sky130_fd_sc_hd__inv_2 _22147_ (.A(_18904_),
    .Y(_19060_));
 sky130_fd_sc_hd__inv_2 _22148_ (.A(\count_cycle[6] ),
    .Y(_01793_));
 sky130_fd_sc_hd__nand2_2 _22149_ (.A(_19060_),
    .B(_01793_),
    .Y(_19061_));
 sky130_fd_sc_hd__and3_2 _22150_ (.A(_19061_),
    .B(_19054_),
    .C(_18905_),
    .X(_03737_));
 sky130_fd_sc_hd__nand2_2 _22151_ (.A(_18903_),
    .B(_01780_),
    .Y(_19062_));
 sky130_fd_sc_hd__and3_2 _22152_ (.A(_19060_),
    .B(_19054_),
    .C(_19062_),
    .X(_03736_));
 sky130_fd_sc_hd__inv_2 _22153_ (.A(_18902_),
    .Y(_19063_));
 sky130_fd_sc_hd__inv_2 _22154_ (.A(\count_cycle[4] ),
    .Y(_01767_));
 sky130_fd_sc_hd__nand2_2 _22155_ (.A(_19063_),
    .B(_01767_),
    .Y(_19064_));
 sky130_fd_sc_hd__and3_2 _22156_ (.A(_19064_),
    .B(_19054_),
    .C(_18903_),
    .X(_03735_));
 sky130_fd_sc_hd__nand2_2 _22157_ (.A(_18901_),
    .B(_01754_),
    .Y(_19065_));
 sky130_fd_sc_hd__and3_2 _22158_ (.A(_19063_),
    .B(_18666_),
    .C(_19065_),
    .X(_03734_));
 sky130_fd_sc_hd__nand2_2 _22159_ (.A(_01741_),
    .B(_18900_),
    .Y(_19066_));
 sky130_fd_sc_hd__and3_2 _22160_ (.A(_18901_),
    .B(_18666_),
    .C(_19066_),
    .X(_03733_));
 sky130_fd_sc_hd__inv_2 _22161_ (.A(\count_cycle[0] ),
    .Y(_02559_));
 sky130_fd_sc_hd__inv_2 _22162_ (.A(\count_cycle[1] ),
    .Y(_01728_));
 sky130_fd_sc_hd__nand2_2 _22163_ (.A(_02559_),
    .B(_01728_),
    .Y(_19067_));
 sky130_fd_sc_hd__and3_2 _22164_ (.A(_19067_),
    .B(_18666_),
    .C(_18900_),
    .X(_03732_));
 sky130_fd_sc_hd__nor2_2 _22165_ (.A(\count_cycle[0] ),
    .B(_18350_),
    .Y(_03731_));
 sky130_fd_sc_hd__nor2_2 _22166_ (.A(_18239_),
    .B(_18445_),
    .Y(_03730_));
 sky130_fd_sc_hd__nor2_2 _22167_ (.A(_18239_),
    .B(_18162_),
    .Y(_03729_));
 sky130_fd_sc_hd__buf_1 _22168_ (.A(\cpuregs_wrdata[31] ),
    .X(_19068_));
 sky130_fd_sc_hd__inv_2 _22169_ (.A(\latched_rd[1] ),
    .Y(_19069_));
 sky130_fd_sc_hd__inv_2 _22170_ (.A(\latched_rd[0] ),
    .Y(_19070_));
 sky130_fd_sc_hd__nand2_2 _22171_ (.A(_19070_),
    .B(_19069_),
    .Y(_19071_));
 sky130_fd_sc_hd__nor2_2 _22172_ (.A(\latched_rd[4] ),
    .B(\latched_rd[2] ),
    .Y(_19072_));
 sky130_fd_sc_hd__inv_2 _22173_ (.A(\latched_rd[3] ),
    .Y(_19073_));
 sky130_fd_sc_hd__nand2_2 _22174_ (.A(_19072_),
    .B(_19073_),
    .Y(_19074_));
 sky130_fd_sc_hd__inv_2 _22175_ (.A(_18145_),
    .Y(_19075_));
 sky130_fd_sc_hd__nor2_2 _22176_ (.A(_18016_),
    .B(_18203_),
    .Y(_19076_));
 sky130_fd_sc_hd__o31a_2 _22177_ (.A1(latched_branch),
    .A2(latched_store),
    .A3(_19075_),
    .B1(_19076_),
    .X(_19077_));
 sky130_fd_sc_hd__o21ai_2 _22178_ (.A1(_19071_),
    .A2(_19074_),
    .B1(_19077_),
    .Y(_19078_));
 sky130_fd_sc_hd__or2_2 _22179_ (.A(_19069_),
    .B(_19078_),
    .X(_19079_));
 sky130_fd_sc_hd__nor2_2 _22180_ (.A(\latched_rd[0] ),
    .B(_19079_),
    .Y(_19080_));
 sky130_fd_sc_hd__inv_2 _22181_ (.A(\latched_rd[4] ),
    .Y(_19081_));
 sky130_fd_sc_hd__and3_2 _22182_ (.A(_19081_),
    .B(_19073_),
    .C(\latched_rd[2] ),
    .X(_19082_));
 sky130_fd_sc_hd__nand2_2 _22183_ (.A(_19080_),
    .B(_19082_),
    .Y(_19083_));
 sky130_fd_sc_hd__buf_1 _22184_ (.A(_19083_),
    .X(_19084_));
 sky130_fd_sc_hd__buf_1 _22185_ (.A(_19084_),
    .X(_19085_));
 sky130_fd_sc_hd__mux2_2 _22186_ (.A0(_19068_),
    .A1(\cpuregs[6][31] ),
    .S(_19085_),
    .X(_03727_));
 sky130_fd_sc_hd__buf_1 _22187_ (.A(\cpuregs_wrdata[30] ),
    .X(_19086_));
 sky130_fd_sc_hd__mux2_2 _22188_ (.A0(_19086_),
    .A1(\cpuregs[6][30] ),
    .S(_19085_),
    .X(_03726_));
 sky130_fd_sc_hd__buf_1 _22189_ (.A(\cpuregs_wrdata[29] ),
    .X(_19087_));
 sky130_fd_sc_hd__mux2_2 _22190_ (.A0(_19087_),
    .A1(\cpuregs[6][29] ),
    .S(_19085_),
    .X(_03725_));
 sky130_fd_sc_hd__buf_1 _22191_ (.A(\cpuregs_wrdata[28] ),
    .X(_19088_));
 sky130_fd_sc_hd__mux2_2 _22192_ (.A0(_19088_),
    .A1(\cpuregs[6][28] ),
    .S(_19085_),
    .X(_03724_));
 sky130_fd_sc_hd__buf_1 _22193_ (.A(\cpuregs_wrdata[27] ),
    .X(_19089_));
 sky130_fd_sc_hd__mux2_2 _22194_ (.A0(_19089_),
    .A1(\cpuregs[6][27] ),
    .S(_19085_),
    .X(_03723_));
 sky130_fd_sc_hd__buf_1 _22195_ (.A(\cpuregs_wrdata[26] ),
    .X(_19090_));
 sky130_fd_sc_hd__mux2_2 _22196_ (.A0(_19090_),
    .A1(\cpuregs[6][26] ),
    .S(_19085_),
    .X(_03722_));
 sky130_fd_sc_hd__buf_1 _22197_ (.A(\cpuregs_wrdata[25] ),
    .X(_19091_));
 sky130_fd_sc_hd__buf_1 _22198_ (.A(_19084_),
    .X(_19092_));
 sky130_fd_sc_hd__mux2_2 _22199_ (.A0(_19091_),
    .A1(\cpuregs[6][25] ),
    .S(_19092_),
    .X(_03721_));
 sky130_fd_sc_hd__buf_1 _22200_ (.A(\cpuregs_wrdata[24] ),
    .X(_19093_));
 sky130_fd_sc_hd__mux2_2 _22201_ (.A0(_19093_),
    .A1(\cpuregs[6][24] ),
    .S(_19092_),
    .X(_03720_));
 sky130_fd_sc_hd__buf_1 _22202_ (.A(\cpuregs_wrdata[23] ),
    .X(_19094_));
 sky130_fd_sc_hd__mux2_2 _22203_ (.A0(_19094_),
    .A1(\cpuregs[6][23] ),
    .S(_19092_),
    .X(_03719_));
 sky130_fd_sc_hd__buf_1 _22204_ (.A(\cpuregs_wrdata[22] ),
    .X(_19095_));
 sky130_fd_sc_hd__mux2_2 _22205_ (.A0(_19095_),
    .A1(\cpuregs[6][22] ),
    .S(_19092_),
    .X(_03718_));
 sky130_fd_sc_hd__buf_1 _22206_ (.A(\cpuregs_wrdata[21] ),
    .X(_19096_));
 sky130_fd_sc_hd__mux2_2 _22207_ (.A0(_19096_),
    .A1(\cpuregs[6][21] ),
    .S(_19092_),
    .X(_03717_));
 sky130_fd_sc_hd__buf_1 _22208_ (.A(\cpuregs_wrdata[20] ),
    .X(_19097_));
 sky130_fd_sc_hd__mux2_2 _22209_ (.A0(_19097_),
    .A1(\cpuregs[6][20] ),
    .S(_19092_),
    .X(_03716_));
 sky130_fd_sc_hd__buf_1 _22210_ (.A(\cpuregs_wrdata[19] ),
    .X(_19098_));
 sky130_fd_sc_hd__buf_1 _22211_ (.A(_19084_),
    .X(_19099_));
 sky130_fd_sc_hd__mux2_2 _22212_ (.A0(_19098_),
    .A1(\cpuregs[6][19] ),
    .S(_19099_),
    .X(_03715_));
 sky130_fd_sc_hd__buf_1 _22213_ (.A(\cpuregs_wrdata[18] ),
    .X(_19100_));
 sky130_fd_sc_hd__mux2_2 _22214_ (.A0(_19100_),
    .A1(\cpuregs[6][18] ),
    .S(_19099_),
    .X(_03714_));
 sky130_fd_sc_hd__buf_1 _22215_ (.A(\cpuregs_wrdata[17] ),
    .X(_19101_));
 sky130_fd_sc_hd__mux2_2 _22216_ (.A0(_19101_),
    .A1(\cpuregs[6][17] ),
    .S(_19099_),
    .X(_03713_));
 sky130_fd_sc_hd__buf_1 _22217_ (.A(\cpuregs_wrdata[16] ),
    .X(_19102_));
 sky130_fd_sc_hd__mux2_2 _22218_ (.A0(_19102_),
    .A1(\cpuregs[6][16] ),
    .S(_19099_),
    .X(_03712_));
 sky130_fd_sc_hd__buf_1 _22219_ (.A(\cpuregs_wrdata[15] ),
    .X(_19103_));
 sky130_fd_sc_hd__mux2_2 _22220_ (.A0(_19103_),
    .A1(\cpuregs[6][15] ),
    .S(_19099_),
    .X(_03711_));
 sky130_fd_sc_hd__buf_1 _22221_ (.A(\cpuregs_wrdata[14] ),
    .X(_19104_));
 sky130_fd_sc_hd__mux2_2 _22222_ (.A0(_19104_),
    .A1(\cpuregs[6][14] ),
    .S(_19099_),
    .X(_03710_));
 sky130_fd_sc_hd__buf_1 _22223_ (.A(\cpuregs_wrdata[13] ),
    .X(_19105_));
 sky130_fd_sc_hd__buf_1 _22224_ (.A(_19084_),
    .X(_19106_));
 sky130_fd_sc_hd__mux2_2 _22225_ (.A0(_19105_),
    .A1(\cpuregs[6][13] ),
    .S(_19106_),
    .X(_03709_));
 sky130_fd_sc_hd__buf_1 _22226_ (.A(\cpuregs_wrdata[12] ),
    .X(_19107_));
 sky130_fd_sc_hd__mux2_2 _22227_ (.A0(_19107_),
    .A1(\cpuregs[6][12] ),
    .S(_19106_),
    .X(_03708_));
 sky130_fd_sc_hd__buf_1 _22228_ (.A(\cpuregs_wrdata[11] ),
    .X(_19108_));
 sky130_fd_sc_hd__mux2_2 _22229_ (.A0(_19108_),
    .A1(\cpuregs[6][11] ),
    .S(_19106_),
    .X(_03707_));
 sky130_fd_sc_hd__buf_1 _22230_ (.A(\cpuregs_wrdata[10] ),
    .X(_19109_));
 sky130_fd_sc_hd__mux2_2 _22231_ (.A0(_19109_),
    .A1(\cpuregs[6][10] ),
    .S(_19106_),
    .X(_03706_));
 sky130_fd_sc_hd__buf_1 _22232_ (.A(\cpuregs_wrdata[9] ),
    .X(_19110_));
 sky130_fd_sc_hd__mux2_2 _22233_ (.A0(_19110_),
    .A1(\cpuregs[6][9] ),
    .S(_19106_),
    .X(_03705_));
 sky130_fd_sc_hd__buf_1 _22234_ (.A(\cpuregs_wrdata[8] ),
    .X(_19111_));
 sky130_fd_sc_hd__mux2_2 _22235_ (.A0(_19111_),
    .A1(\cpuregs[6][8] ),
    .S(_19106_),
    .X(_03704_));
 sky130_fd_sc_hd__buf_1 _22236_ (.A(\cpuregs_wrdata[7] ),
    .X(_19112_));
 sky130_fd_sc_hd__buf_1 _22237_ (.A(_19083_),
    .X(_19113_));
 sky130_fd_sc_hd__mux2_2 _22238_ (.A0(_19112_),
    .A1(\cpuregs[6][7] ),
    .S(_19113_),
    .X(_03703_));
 sky130_fd_sc_hd__buf_1 _22239_ (.A(\cpuregs_wrdata[6] ),
    .X(_19114_));
 sky130_fd_sc_hd__mux2_2 _22240_ (.A0(_19114_),
    .A1(\cpuregs[6][6] ),
    .S(_19113_),
    .X(_03702_));
 sky130_fd_sc_hd__buf_1 _22241_ (.A(\cpuregs_wrdata[5] ),
    .X(_19115_));
 sky130_fd_sc_hd__mux2_2 _22242_ (.A0(_19115_),
    .A1(\cpuregs[6][5] ),
    .S(_19113_),
    .X(_03701_));
 sky130_fd_sc_hd__buf_1 _22243_ (.A(\cpuregs_wrdata[4] ),
    .X(_19116_));
 sky130_fd_sc_hd__mux2_2 _22244_ (.A0(_19116_),
    .A1(\cpuregs[6][4] ),
    .S(_19113_),
    .X(_03700_));
 sky130_fd_sc_hd__buf_1 _22245_ (.A(\cpuregs_wrdata[3] ),
    .X(_19117_));
 sky130_fd_sc_hd__mux2_2 _22246_ (.A0(_19117_),
    .A1(\cpuregs[6][3] ),
    .S(_19113_),
    .X(_03699_));
 sky130_fd_sc_hd__buf_1 _22247_ (.A(\cpuregs_wrdata[2] ),
    .X(_19118_));
 sky130_fd_sc_hd__mux2_2 _22248_ (.A0(_19118_),
    .A1(\cpuregs[6][2] ),
    .S(_19113_),
    .X(_03698_));
 sky130_fd_sc_hd__buf_1 _22249_ (.A(\cpuregs_wrdata[1] ),
    .X(_19119_));
 sky130_fd_sc_hd__mux2_2 _22250_ (.A0(_19119_),
    .A1(\cpuregs[6][1] ),
    .S(_19084_),
    .X(_03697_));
 sky130_fd_sc_hd__buf_1 _22251_ (.A(\cpuregs_wrdata[0] ),
    .X(_19120_));
 sky130_fd_sc_hd__mux2_2 _22252_ (.A0(_19120_),
    .A1(\cpuregs[6][0] ),
    .S(_19084_),
    .X(_03696_));
 sky130_fd_sc_hd__nor3_2 _22253_ (.A(_19070_),
    .B(\latched_rd[1] ),
    .C(_19078_),
    .Y(_19121_));
 sky130_fd_sc_hd__nand2_2 _22254_ (.A(_19072_),
    .B(\latched_rd[3] ),
    .Y(_19122_));
 sky130_fd_sc_hd__inv_2 _22255_ (.A(_19122_),
    .Y(_19123_));
 sky130_fd_sc_hd__nand2_2 _22256_ (.A(_19121_),
    .B(_19123_),
    .Y(_19124_));
 sky130_fd_sc_hd__buf_1 _22257_ (.A(_19124_),
    .X(_19125_));
 sky130_fd_sc_hd__buf_1 _22258_ (.A(_19125_),
    .X(_19126_));
 sky130_fd_sc_hd__mux2_2 _22259_ (.A0(_19068_),
    .A1(\cpuregs[9][31] ),
    .S(_19126_),
    .X(_03695_));
 sky130_fd_sc_hd__mux2_2 _22260_ (.A0(_19086_),
    .A1(\cpuregs[9][30] ),
    .S(_19126_),
    .X(_03694_));
 sky130_fd_sc_hd__mux2_2 _22261_ (.A0(_19087_),
    .A1(\cpuregs[9][29] ),
    .S(_19126_),
    .X(_03693_));
 sky130_fd_sc_hd__mux2_2 _22262_ (.A0(_19088_),
    .A1(\cpuregs[9][28] ),
    .S(_19126_),
    .X(_03692_));
 sky130_fd_sc_hd__mux2_2 _22263_ (.A0(_19089_),
    .A1(\cpuregs[9][27] ),
    .S(_19126_),
    .X(_03691_));
 sky130_fd_sc_hd__mux2_2 _22264_ (.A0(_19090_),
    .A1(\cpuregs[9][26] ),
    .S(_19126_),
    .X(_03690_));
 sky130_fd_sc_hd__buf_1 _22265_ (.A(_19125_),
    .X(_19127_));
 sky130_fd_sc_hd__mux2_2 _22266_ (.A0(_19091_),
    .A1(\cpuregs[9][25] ),
    .S(_19127_),
    .X(_03689_));
 sky130_fd_sc_hd__mux2_2 _22267_ (.A0(_19093_),
    .A1(\cpuregs[9][24] ),
    .S(_19127_),
    .X(_03688_));
 sky130_fd_sc_hd__mux2_2 _22268_ (.A0(_19094_),
    .A1(\cpuregs[9][23] ),
    .S(_19127_),
    .X(_03687_));
 sky130_fd_sc_hd__mux2_2 _22269_ (.A0(_19095_),
    .A1(\cpuregs[9][22] ),
    .S(_19127_),
    .X(_03686_));
 sky130_fd_sc_hd__mux2_2 _22270_ (.A0(_19096_),
    .A1(\cpuregs[9][21] ),
    .S(_19127_),
    .X(_03685_));
 sky130_fd_sc_hd__mux2_2 _22271_ (.A0(_19097_),
    .A1(\cpuregs[9][20] ),
    .S(_19127_),
    .X(_03684_));
 sky130_fd_sc_hd__buf_1 _22272_ (.A(_19125_),
    .X(_19128_));
 sky130_fd_sc_hd__mux2_2 _22273_ (.A0(_19098_),
    .A1(\cpuregs[9][19] ),
    .S(_19128_),
    .X(_03683_));
 sky130_fd_sc_hd__mux2_2 _22274_ (.A0(_19100_),
    .A1(\cpuregs[9][18] ),
    .S(_19128_),
    .X(_03682_));
 sky130_fd_sc_hd__mux2_2 _22275_ (.A0(_19101_),
    .A1(\cpuregs[9][17] ),
    .S(_19128_),
    .X(_03681_));
 sky130_fd_sc_hd__mux2_2 _22276_ (.A0(_19102_),
    .A1(\cpuregs[9][16] ),
    .S(_19128_),
    .X(_03680_));
 sky130_fd_sc_hd__mux2_2 _22277_ (.A0(_19103_),
    .A1(\cpuregs[9][15] ),
    .S(_19128_),
    .X(_03679_));
 sky130_fd_sc_hd__mux2_2 _22278_ (.A0(_19104_),
    .A1(\cpuregs[9][14] ),
    .S(_19128_),
    .X(_03678_));
 sky130_fd_sc_hd__buf_1 _22279_ (.A(_19125_),
    .X(_19129_));
 sky130_fd_sc_hd__mux2_2 _22280_ (.A0(_19105_),
    .A1(\cpuregs[9][13] ),
    .S(_19129_),
    .X(_03677_));
 sky130_fd_sc_hd__mux2_2 _22281_ (.A0(_19107_),
    .A1(\cpuregs[9][12] ),
    .S(_19129_),
    .X(_03676_));
 sky130_fd_sc_hd__mux2_2 _22282_ (.A0(_19108_),
    .A1(\cpuregs[9][11] ),
    .S(_19129_),
    .X(_03675_));
 sky130_fd_sc_hd__mux2_2 _22283_ (.A0(_19109_),
    .A1(\cpuregs[9][10] ),
    .S(_19129_),
    .X(_03674_));
 sky130_fd_sc_hd__mux2_2 _22284_ (.A0(_19110_),
    .A1(\cpuregs[9][9] ),
    .S(_19129_),
    .X(_03673_));
 sky130_fd_sc_hd__mux2_2 _22285_ (.A0(_19111_),
    .A1(\cpuregs[9][8] ),
    .S(_19129_),
    .X(_03672_));
 sky130_fd_sc_hd__buf_1 _22286_ (.A(_19124_),
    .X(_19130_));
 sky130_fd_sc_hd__mux2_2 _22287_ (.A0(_19112_),
    .A1(\cpuregs[9][7] ),
    .S(_19130_),
    .X(_03671_));
 sky130_fd_sc_hd__mux2_2 _22288_ (.A0(_19114_),
    .A1(\cpuregs[9][6] ),
    .S(_19130_),
    .X(_03670_));
 sky130_fd_sc_hd__mux2_2 _22289_ (.A0(_19115_),
    .A1(\cpuregs[9][5] ),
    .S(_19130_),
    .X(_03669_));
 sky130_fd_sc_hd__mux2_2 _22290_ (.A0(_19116_),
    .A1(\cpuregs[9][4] ),
    .S(_19130_),
    .X(_03668_));
 sky130_fd_sc_hd__mux2_2 _22291_ (.A0(_19117_),
    .A1(\cpuregs[9][3] ),
    .S(_19130_),
    .X(_03667_));
 sky130_fd_sc_hd__mux2_2 _22292_ (.A0(_19118_),
    .A1(\cpuregs[9][2] ),
    .S(_19130_),
    .X(_03666_));
 sky130_fd_sc_hd__mux2_2 _22293_ (.A0(_19119_),
    .A1(\cpuregs[9][1] ),
    .S(_19125_),
    .X(_03665_));
 sky130_fd_sc_hd__mux2_2 _22294_ (.A0(_19120_),
    .A1(\cpuregs[9][0] ),
    .S(_19125_),
    .X(_03664_));
 sky130_fd_sc_hd__nor2_2 _22295_ (.A(_18048_),
    .B(_18443_),
    .Y(_19131_));
 sky130_fd_sc_hd__buf_1 _22296_ (.A(_19131_),
    .X(_19132_));
 sky130_fd_sc_hd__buf_1 _22297_ (.A(_19132_),
    .X(_19133_));
 sky130_fd_sc_hd__mux2_2 _22298_ (.A0(pcpi_rs2[31]),
    .A1(_02467_),
    .S(_19133_),
    .X(_03663_));
 sky130_fd_sc_hd__mux2_2 _22299_ (.A0(pcpi_rs2[30]),
    .A1(_02466_),
    .S(_19133_),
    .X(_03662_));
 sky130_fd_sc_hd__buf_1 _22300_ (.A(pcpi_rs2[29]),
    .X(_19134_));
 sky130_fd_sc_hd__mux2_2 _22301_ (.A0(_19134_),
    .A1(_02464_),
    .S(_19133_),
    .X(_03661_));
 sky130_fd_sc_hd__mux2_2 _22302_ (.A0(pcpi_rs2[28]),
    .A1(_02463_),
    .S(_19133_),
    .X(_03660_));
 sky130_fd_sc_hd__buf_1 _22303_ (.A(pcpi_rs2[27]),
    .X(_19135_));
 sky130_fd_sc_hd__mux2_2 _22304_ (.A0(_19135_),
    .A1(_02462_),
    .S(_19133_),
    .X(_03659_));
 sky130_fd_sc_hd__buf_1 _22305_ (.A(_19132_),
    .X(_19136_));
 sky130_fd_sc_hd__mux2_2 _22306_ (.A0(pcpi_rs2[26]),
    .A1(_02461_),
    .S(_19136_),
    .X(_03658_));
 sky130_fd_sc_hd__buf_1 _22307_ (.A(pcpi_rs2[25]),
    .X(_19137_));
 sky130_fd_sc_hd__mux2_2 _22308_ (.A0(_19137_),
    .A1(_02460_),
    .S(_19136_),
    .X(_03657_));
 sky130_fd_sc_hd__mux2_2 _22309_ (.A0(pcpi_rs2[24]),
    .A1(_02459_),
    .S(_19136_),
    .X(_03656_));
 sky130_fd_sc_hd__buf_1 _22310_ (.A(pcpi_rs2[23]),
    .X(_19138_));
 sky130_fd_sc_hd__mux2_2 _22311_ (.A0(_19138_),
    .A1(_02458_),
    .S(_19136_),
    .X(_03655_));
 sky130_fd_sc_hd__mux2_2 _22312_ (.A0(pcpi_rs2[22]),
    .A1(_02457_),
    .S(_19136_),
    .X(_03654_));
 sky130_fd_sc_hd__buf_1 _22313_ (.A(pcpi_rs2[21]),
    .X(_19139_));
 sky130_fd_sc_hd__mux2_2 _22314_ (.A0(_19139_),
    .A1(_02456_),
    .S(_19136_),
    .X(_03653_));
 sky130_fd_sc_hd__buf_1 _22315_ (.A(_19132_),
    .X(_19140_));
 sky130_fd_sc_hd__mux2_2 _22316_ (.A0(pcpi_rs2[20]),
    .A1(_02455_),
    .S(_19140_),
    .X(_03652_));
 sky130_fd_sc_hd__mux2_2 _22317_ (.A0(pcpi_rs2[19]),
    .A1(_02453_),
    .S(_19140_),
    .X(_03651_));
 sky130_fd_sc_hd__buf_1 _22318_ (.A(pcpi_rs2[18]),
    .X(_19141_));
 sky130_fd_sc_hd__mux2_2 _22319_ (.A0(_19141_),
    .A1(_02452_),
    .S(_19140_),
    .X(_03650_));
 sky130_fd_sc_hd__mux2_2 _22320_ (.A0(pcpi_rs2[17]),
    .A1(_02451_),
    .S(_19140_),
    .X(_03649_));
 sky130_fd_sc_hd__mux2_2 _22321_ (.A0(pcpi_rs2[16]),
    .A1(_02450_),
    .S(_19140_),
    .X(_03648_));
 sky130_fd_sc_hd__buf_1 _22322_ (.A(pcpi_rs2[15]),
    .X(_19142_));
 sky130_fd_sc_hd__mux2_2 _22323_ (.A0(_19142_),
    .A1(_02449_),
    .S(_19140_),
    .X(_03647_));
 sky130_fd_sc_hd__buf_1 _22324_ (.A(pcpi_rs2[14]),
    .X(_19143_));
 sky130_fd_sc_hd__buf_1 _22325_ (.A(_19131_),
    .X(_19144_));
 sky130_fd_sc_hd__mux2_2 _22326_ (.A0(_19143_),
    .A1(_02448_),
    .S(_19144_),
    .X(_03646_));
 sky130_fd_sc_hd__buf_1 _22327_ (.A(pcpi_rs2[13]),
    .X(_19145_));
 sky130_fd_sc_hd__mux2_2 _22328_ (.A0(_19145_),
    .A1(_02447_),
    .S(_19144_),
    .X(_03645_));
 sky130_fd_sc_hd__mux2_2 _22329_ (.A0(pcpi_rs2[12]),
    .A1(_02446_),
    .S(_19144_),
    .X(_03644_));
 sky130_fd_sc_hd__buf_1 _22330_ (.A(pcpi_rs2[11]),
    .X(_19146_));
 sky130_fd_sc_hd__mux2_2 _22331_ (.A0(_19146_),
    .A1(_02445_),
    .S(_19144_),
    .X(_03643_));
 sky130_fd_sc_hd__mux2_2 _22332_ (.A0(pcpi_rs2[10]),
    .A1(_02444_),
    .S(_19144_),
    .X(_03642_));
 sky130_fd_sc_hd__buf_1 _22333_ (.A(pcpi_rs2[9]),
    .X(_19147_));
 sky130_fd_sc_hd__mux2_2 _22334_ (.A0(_19147_),
    .A1(_02474_),
    .S(_19144_),
    .X(_03641_));
 sky130_fd_sc_hd__buf_1 _22335_ (.A(_19131_),
    .X(_19148_));
 sky130_fd_sc_hd__mux2_2 _22336_ (.A0(pcpi_rs2[8]),
    .A1(_02473_),
    .S(_19148_),
    .X(_03640_));
 sky130_fd_sc_hd__buf_1 _22337_ (.A(mem_la_wdata[7]),
    .X(_19149_));
 sky130_fd_sc_hd__mux2_2 _22338_ (.A0(_19149_),
    .A1(_02472_),
    .S(_19148_),
    .X(_03639_));
 sky130_fd_sc_hd__buf_1 _22339_ (.A(mem_la_wdata[6]),
    .X(_19150_));
 sky130_fd_sc_hd__mux2_2 _22340_ (.A0(_19150_),
    .A1(_02471_),
    .S(_19148_),
    .X(_03638_));
 sky130_fd_sc_hd__buf_1 _22341_ (.A(mem_la_wdata[5]),
    .X(_19151_));
 sky130_fd_sc_hd__mux2_2 _22342_ (.A0(_19151_),
    .A1(_02470_),
    .S(_19148_),
    .X(_03637_));
 sky130_fd_sc_hd__buf_1 _22343_ (.A(mem_la_wdata[4]),
    .X(_19152_));
 sky130_fd_sc_hd__mux2_2 _22344_ (.A0(_19152_),
    .A1(_02469_),
    .S(_19148_),
    .X(_03636_));
 sky130_fd_sc_hd__buf_1 _22345_ (.A(mem_la_wdata[3]),
    .X(_19153_));
 sky130_fd_sc_hd__mux2_2 _22346_ (.A0(_19153_),
    .A1(_02468_),
    .S(_19148_),
    .X(_03635_));
 sky130_fd_sc_hd__buf_1 _22347_ (.A(mem_la_wdata[2]),
    .X(_19154_));
 sky130_fd_sc_hd__mux2_2 _22348_ (.A0(_19154_),
    .A1(_02465_),
    .S(_19132_),
    .X(_03634_));
 sky130_fd_sc_hd__buf_1 _22349_ (.A(mem_la_wdata[1]),
    .X(_19155_));
 sky130_fd_sc_hd__mux2_2 _22350_ (.A0(_19155_),
    .A1(_02454_),
    .S(_19132_),
    .X(_03633_));
 sky130_fd_sc_hd__buf_1 _22351_ (.A(mem_la_wdata[0]),
    .X(_19156_));
 sky130_fd_sc_hd__mux2_2 _22352_ (.A0(_19156_),
    .A1(_02443_),
    .S(_19132_),
    .X(_03632_));
 sky130_fd_sc_hd__or3b_2 _22353_ (.A(_19071_),
    .B(_19078_),
    .C_N(_19082_),
    .X(_19157_));
 sky130_fd_sc_hd__buf_1 _22354_ (.A(_19157_),
    .X(_19158_));
 sky130_fd_sc_hd__buf_1 _22355_ (.A(_19158_),
    .X(_19159_));
 sky130_fd_sc_hd__mux2_2 _22356_ (.A0(_19068_),
    .A1(\cpuregs[4][31] ),
    .S(_19159_),
    .X(_03631_));
 sky130_fd_sc_hd__mux2_2 _22357_ (.A0(_19086_),
    .A1(\cpuregs[4][30] ),
    .S(_19159_),
    .X(_03630_));
 sky130_fd_sc_hd__mux2_2 _22358_ (.A0(_19087_),
    .A1(\cpuregs[4][29] ),
    .S(_19159_),
    .X(_03629_));
 sky130_fd_sc_hd__mux2_2 _22359_ (.A0(_19088_),
    .A1(\cpuregs[4][28] ),
    .S(_19159_),
    .X(_03628_));
 sky130_fd_sc_hd__mux2_2 _22360_ (.A0(_19089_),
    .A1(\cpuregs[4][27] ),
    .S(_19159_),
    .X(_03627_));
 sky130_fd_sc_hd__mux2_2 _22361_ (.A0(_19090_),
    .A1(\cpuregs[4][26] ),
    .S(_19159_),
    .X(_03626_));
 sky130_fd_sc_hd__buf_1 _22362_ (.A(_19158_),
    .X(_19160_));
 sky130_fd_sc_hd__mux2_2 _22363_ (.A0(_19091_),
    .A1(\cpuregs[4][25] ),
    .S(_19160_),
    .X(_03625_));
 sky130_fd_sc_hd__mux2_2 _22364_ (.A0(_19093_),
    .A1(\cpuregs[4][24] ),
    .S(_19160_),
    .X(_03624_));
 sky130_fd_sc_hd__mux2_2 _22365_ (.A0(_19094_),
    .A1(\cpuregs[4][23] ),
    .S(_19160_),
    .X(_03623_));
 sky130_fd_sc_hd__mux2_2 _22366_ (.A0(_19095_),
    .A1(\cpuregs[4][22] ),
    .S(_19160_),
    .X(_03622_));
 sky130_fd_sc_hd__mux2_2 _22367_ (.A0(_19096_),
    .A1(\cpuregs[4][21] ),
    .S(_19160_),
    .X(_03621_));
 sky130_fd_sc_hd__mux2_2 _22368_ (.A0(_19097_),
    .A1(\cpuregs[4][20] ),
    .S(_19160_),
    .X(_03620_));
 sky130_fd_sc_hd__buf_1 _22369_ (.A(_19158_),
    .X(_19161_));
 sky130_fd_sc_hd__mux2_2 _22370_ (.A0(_19098_),
    .A1(\cpuregs[4][19] ),
    .S(_19161_),
    .X(_03619_));
 sky130_fd_sc_hd__mux2_2 _22371_ (.A0(_19100_),
    .A1(\cpuregs[4][18] ),
    .S(_19161_),
    .X(_03618_));
 sky130_fd_sc_hd__mux2_2 _22372_ (.A0(_19101_),
    .A1(\cpuregs[4][17] ),
    .S(_19161_),
    .X(_03617_));
 sky130_fd_sc_hd__mux2_2 _22373_ (.A0(_19102_),
    .A1(\cpuregs[4][16] ),
    .S(_19161_),
    .X(_03616_));
 sky130_fd_sc_hd__mux2_2 _22374_ (.A0(_19103_),
    .A1(\cpuregs[4][15] ),
    .S(_19161_),
    .X(_03615_));
 sky130_fd_sc_hd__mux2_2 _22375_ (.A0(_19104_),
    .A1(\cpuregs[4][14] ),
    .S(_19161_),
    .X(_03614_));
 sky130_fd_sc_hd__buf_1 _22376_ (.A(_19158_),
    .X(_19162_));
 sky130_fd_sc_hd__mux2_2 _22377_ (.A0(_19105_),
    .A1(\cpuregs[4][13] ),
    .S(_19162_),
    .X(_03613_));
 sky130_fd_sc_hd__mux2_2 _22378_ (.A0(_19107_),
    .A1(\cpuregs[4][12] ),
    .S(_19162_),
    .X(_03612_));
 sky130_fd_sc_hd__mux2_2 _22379_ (.A0(_19108_),
    .A1(\cpuregs[4][11] ),
    .S(_19162_),
    .X(_03611_));
 sky130_fd_sc_hd__mux2_2 _22380_ (.A0(_19109_),
    .A1(\cpuregs[4][10] ),
    .S(_19162_),
    .X(_03610_));
 sky130_fd_sc_hd__mux2_2 _22381_ (.A0(_19110_),
    .A1(\cpuregs[4][9] ),
    .S(_19162_),
    .X(_03609_));
 sky130_fd_sc_hd__mux2_2 _22382_ (.A0(_19111_),
    .A1(\cpuregs[4][8] ),
    .S(_19162_),
    .X(_03608_));
 sky130_fd_sc_hd__buf_1 _22383_ (.A(_19157_),
    .X(_19163_));
 sky130_fd_sc_hd__mux2_2 _22384_ (.A0(_19112_),
    .A1(\cpuregs[4][7] ),
    .S(_19163_),
    .X(_03607_));
 sky130_fd_sc_hd__mux2_2 _22385_ (.A0(_19114_),
    .A1(\cpuregs[4][6] ),
    .S(_19163_),
    .X(_03606_));
 sky130_fd_sc_hd__mux2_2 _22386_ (.A0(_19115_),
    .A1(\cpuregs[4][5] ),
    .S(_19163_),
    .X(_03605_));
 sky130_fd_sc_hd__mux2_2 _22387_ (.A0(_19116_),
    .A1(\cpuregs[4][4] ),
    .S(_19163_),
    .X(_03604_));
 sky130_fd_sc_hd__mux2_2 _22388_ (.A0(_19117_),
    .A1(\cpuregs[4][3] ),
    .S(_19163_),
    .X(_03603_));
 sky130_fd_sc_hd__mux2_2 _22389_ (.A0(_19118_),
    .A1(\cpuregs[4][2] ),
    .S(_19163_),
    .X(_03602_));
 sky130_fd_sc_hd__mux2_2 _22390_ (.A0(_19119_),
    .A1(\cpuregs[4][1] ),
    .S(_19158_),
    .X(_03601_));
 sky130_fd_sc_hd__mux2_2 _22391_ (.A0(_19120_),
    .A1(\cpuregs[4][0] ),
    .S(_19158_),
    .X(_03600_));
 sky130_fd_sc_hd__nor2_2 _22392_ (.A(_19070_),
    .B(_19079_),
    .Y(_19164_));
 sky130_fd_sc_hd__nor3_2 _22393_ (.A(\latched_rd[2] ),
    .B(\latched_rd[3] ),
    .C(_19081_),
    .Y(_19165_));
 sky130_fd_sc_hd__nand2_2 _22394_ (.A(_19164_),
    .B(_19165_),
    .Y(_19166_));
 sky130_fd_sc_hd__buf_1 _22395_ (.A(_19166_),
    .X(_19167_));
 sky130_fd_sc_hd__buf_1 _22396_ (.A(_19167_),
    .X(_19168_));
 sky130_fd_sc_hd__mux2_2 _22397_ (.A0(_19068_),
    .A1(\cpuregs[19][31] ),
    .S(_19168_),
    .X(_03599_));
 sky130_fd_sc_hd__mux2_2 _22398_ (.A0(_19086_),
    .A1(\cpuregs[19][30] ),
    .S(_19168_),
    .X(_03598_));
 sky130_fd_sc_hd__mux2_2 _22399_ (.A0(_19087_),
    .A1(\cpuregs[19][29] ),
    .S(_19168_),
    .X(_03597_));
 sky130_fd_sc_hd__mux2_2 _22400_ (.A0(_19088_),
    .A1(\cpuregs[19][28] ),
    .S(_19168_),
    .X(_03596_));
 sky130_fd_sc_hd__mux2_2 _22401_ (.A0(_19089_),
    .A1(\cpuregs[19][27] ),
    .S(_19168_),
    .X(_03595_));
 sky130_fd_sc_hd__mux2_2 _22402_ (.A0(_19090_),
    .A1(\cpuregs[19][26] ),
    .S(_19168_),
    .X(_03594_));
 sky130_fd_sc_hd__buf_1 _22403_ (.A(_19167_),
    .X(_19169_));
 sky130_fd_sc_hd__mux2_2 _22404_ (.A0(_19091_),
    .A1(\cpuregs[19][25] ),
    .S(_19169_),
    .X(_03593_));
 sky130_fd_sc_hd__mux2_2 _22405_ (.A0(_19093_),
    .A1(\cpuregs[19][24] ),
    .S(_19169_),
    .X(_03592_));
 sky130_fd_sc_hd__mux2_2 _22406_ (.A0(_19094_),
    .A1(\cpuregs[19][23] ),
    .S(_19169_),
    .X(_03591_));
 sky130_fd_sc_hd__mux2_2 _22407_ (.A0(_19095_),
    .A1(\cpuregs[19][22] ),
    .S(_19169_),
    .X(_03590_));
 sky130_fd_sc_hd__mux2_2 _22408_ (.A0(_19096_),
    .A1(\cpuregs[19][21] ),
    .S(_19169_),
    .X(_03589_));
 sky130_fd_sc_hd__mux2_2 _22409_ (.A0(_19097_),
    .A1(\cpuregs[19][20] ),
    .S(_19169_),
    .X(_03588_));
 sky130_fd_sc_hd__buf_1 _22410_ (.A(_19167_),
    .X(_19170_));
 sky130_fd_sc_hd__mux2_2 _22411_ (.A0(_19098_),
    .A1(\cpuregs[19][19] ),
    .S(_19170_),
    .X(_03587_));
 sky130_fd_sc_hd__mux2_2 _22412_ (.A0(_19100_),
    .A1(\cpuregs[19][18] ),
    .S(_19170_),
    .X(_03586_));
 sky130_fd_sc_hd__mux2_2 _22413_ (.A0(_19101_),
    .A1(\cpuregs[19][17] ),
    .S(_19170_),
    .X(_03585_));
 sky130_fd_sc_hd__mux2_2 _22414_ (.A0(_19102_),
    .A1(\cpuregs[19][16] ),
    .S(_19170_),
    .X(_03584_));
 sky130_fd_sc_hd__mux2_2 _22415_ (.A0(_19103_),
    .A1(\cpuregs[19][15] ),
    .S(_19170_),
    .X(_03583_));
 sky130_fd_sc_hd__mux2_2 _22416_ (.A0(_19104_),
    .A1(\cpuregs[19][14] ),
    .S(_19170_),
    .X(_03582_));
 sky130_fd_sc_hd__buf_1 _22417_ (.A(_19167_),
    .X(_19171_));
 sky130_fd_sc_hd__mux2_2 _22418_ (.A0(_19105_),
    .A1(\cpuregs[19][13] ),
    .S(_19171_),
    .X(_03581_));
 sky130_fd_sc_hd__mux2_2 _22419_ (.A0(_19107_),
    .A1(\cpuregs[19][12] ),
    .S(_19171_),
    .X(_03580_));
 sky130_fd_sc_hd__mux2_2 _22420_ (.A0(_19108_),
    .A1(\cpuregs[19][11] ),
    .S(_19171_),
    .X(_03579_));
 sky130_fd_sc_hd__mux2_2 _22421_ (.A0(_19109_),
    .A1(\cpuregs[19][10] ),
    .S(_19171_),
    .X(_03578_));
 sky130_fd_sc_hd__mux2_2 _22422_ (.A0(_19110_),
    .A1(\cpuregs[19][9] ),
    .S(_19171_),
    .X(_03577_));
 sky130_fd_sc_hd__mux2_2 _22423_ (.A0(_19111_),
    .A1(\cpuregs[19][8] ),
    .S(_19171_),
    .X(_03576_));
 sky130_fd_sc_hd__buf_1 _22424_ (.A(_19166_),
    .X(_19172_));
 sky130_fd_sc_hd__mux2_2 _22425_ (.A0(_19112_),
    .A1(\cpuregs[19][7] ),
    .S(_19172_),
    .X(_03575_));
 sky130_fd_sc_hd__mux2_2 _22426_ (.A0(_19114_),
    .A1(\cpuregs[19][6] ),
    .S(_19172_),
    .X(_03574_));
 sky130_fd_sc_hd__mux2_2 _22427_ (.A0(_19115_),
    .A1(\cpuregs[19][5] ),
    .S(_19172_),
    .X(_03573_));
 sky130_fd_sc_hd__mux2_2 _22428_ (.A0(_19116_),
    .A1(\cpuregs[19][4] ),
    .S(_19172_),
    .X(_03572_));
 sky130_fd_sc_hd__mux2_2 _22429_ (.A0(_19117_),
    .A1(\cpuregs[19][3] ),
    .S(_19172_),
    .X(_03571_));
 sky130_fd_sc_hd__mux2_2 _22430_ (.A0(_19118_),
    .A1(\cpuregs[19][2] ),
    .S(_19172_),
    .X(_03570_));
 sky130_fd_sc_hd__mux2_2 _22431_ (.A0(_19119_),
    .A1(\cpuregs[19][1] ),
    .S(_19167_),
    .X(_03569_));
 sky130_fd_sc_hd__mux2_2 _22432_ (.A0(_19120_),
    .A1(\cpuregs[19][0] ),
    .S(_19167_),
    .X(_03568_));
 sky130_fd_sc_hd__and3_2 _22433_ (.A(_00290_),
    .B(_18024_),
    .C(mem_do_wdata),
    .X(_19173_));
 sky130_fd_sc_hd__buf_1 _22434_ (.A(_19173_),
    .X(mem_la_write));
 sky130_fd_sc_hd__nand2_2 _22435_ (.A(mem_la_write),
    .B(_18047_),
    .Y(_19174_));
 sky130_fd_sc_hd__buf_1 _22436_ (.A(_19174_),
    .X(_19175_));
 sky130_fd_sc_hd__buf_1 _22437_ (.A(_19175_),
    .X(_19176_));
 sky130_fd_sc_hd__mux2_2 _22438_ (.A0(mem_la_wdata[31]),
    .A1(mem_wdata[31]),
    .S(_19176_),
    .X(_03567_));
 sky130_fd_sc_hd__mux2_2 _22439_ (.A0(mem_la_wdata[30]),
    .A1(mem_wdata[30]),
    .S(_19176_),
    .X(_03566_));
 sky130_fd_sc_hd__mux2_2 _22440_ (.A0(mem_la_wdata[29]),
    .A1(mem_wdata[29]),
    .S(_19176_),
    .X(_03565_));
 sky130_fd_sc_hd__mux2_2 _22441_ (.A0(mem_la_wdata[28]),
    .A1(mem_wdata[28]),
    .S(_19176_),
    .X(_03564_));
 sky130_fd_sc_hd__mux2_2 _22442_ (.A0(mem_la_wdata[27]),
    .A1(mem_wdata[27]),
    .S(_19176_),
    .X(_03563_));
 sky130_fd_sc_hd__mux2_2 _22443_ (.A0(mem_la_wdata[26]),
    .A1(mem_wdata[26]),
    .S(_19176_),
    .X(_03562_));
 sky130_fd_sc_hd__buf_1 _22444_ (.A(_19175_),
    .X(_19177_));
 sky130_fd_sc_hd__mux2_2 _22445_ (.A0(mem_la_wdata[25]),
    .A1(mem_wdata[25]),
    .S(_19177_),
    .X(_03561_));
 sky130_fd_sc_hd__mux2_2 _22446_ (.A0(mem_la_wdata[24]),
    .A1(mem_wdata[24]),
    .S(_19177_),
    .X(_03560_));
 sky130_fd_sc_hd__mux2_2 _22447_ (.A0(mem_la_wdata[23]),
    .A1(mem_wdata[23]),
    .S(_19177_),
    .X(_03559_));
 sky130_fd_sc_hd__mux2_2 _22448_ (.A0(mem_la_wdata[22]),
    .A1(mem_wdata[22]),
    .S(_19177_),
    .X(_03558_));
 sky130_fd_sc_hd__mux2_2 _22449_ (.A0(mem_la_wdata[21]),
    .A1(mem_wdata[21]),
    .S(_19177_),
    .X(_03557_));
 sky130_fd_sc_hd__mux2_2 _22450_ (.A0(mem_la_wdata[20]),
    .A1(mem_wdata[20]),
    .S(_19177_),
    .X(_03556_));
 sky130_fd_sc_hd__buf_1 _22451_ (.A(_19175_),
    .X(_19178_));
 sky130_fd_sc_hd__mux2_2 _22452_ (.A0(mem_la_wdata[19]),
    .A1(mem_wdata[19]),
    .S(_19178_),
    .X(_03555_));
 sky130_fd_sc_hd__mux2_2 _22453_ (.A0(mem_la_wdata[18]),
    .A1(mem_wdata[18]),
    .S(_19178_),
    .X(_03554_));
 sky130_fd_sc_hd__mux2_2 _22454_ (.A0(mem_la_wdata[17]),
    .A1(mem_wdata[17]),
    .S(_19178_),
    .X(_03553_));
 sky130_fd_sc_hd__mux2_2 _22455_ (.A0(mem_la_wdata[16]),
    .A1(mem_wdata[16]),
    .S(_19178_),
    .X(_03552_));
 sky130_fd_sc_hd__mux2_2 _22456_ (.A0(mem_la_wdata[15]),
    .A1(mem_wdata[15]),
    .S(_19178_),
    .X(_03551_));
 sky130_fd_sc_hd__mux2_2 _22457_ (.A0(mem_la_wdata[14]),
    .A1(mem_wdata[14]),
    .S(_19178_),
    .X(_03550_));
 sky130_fd_sc_hd__buf_1 _22458_ (.A(_19175_),
    .X(_19179_));
 sky130_fd_sc_hd__mux2_2 _22459_ (.A0(mem_la_wdata[13]),
    .A1(mem_wdata[13]),
    .S(_19179_),
    .X(_03549_));
 sky130_fd_sc_hd__mux2_2 _22460_ (.A0(mem_la_wdata[12]),
    .A1(mem_wdata[12]),
    .S(_19179_),
    .X(_03548_));
 sky130_fd_sc_hd__mux2_2 _22461_ (.A0(mem_la_wdata[11]),
    .A1(mem_wdata[11]),
    .S(_19179_),
    .X(_03547_));
 sky130_fd_sc_hd__mux2_2 _22462_ (.A0(mem_la_wdata[10]),
    .A1(mem_wdata[10]),
    .S(_19179_),
    .X(_03546_));
 sky130_fd_sc_hd__mux2_2 _22463_ (.A0(mem_la_wdata[9]),
    .A1(mem_wdata[9]),
    .S(_19179_),
    .X(_03545_));
 sky130_fd_sc_hd__mux2_2 _22464_ (.A0(mem_la_wdata[8]),
    .A1(mem_wdata[8]),
    .S(_19179_),
    .X(_03544_));
 sky130_fd_sc_hd__buf_1 _22465_ (.A(_19174_),
    .X(_19180_));
 sky130_fd_sc_hd__mux2_2 _22466_ (.A0(_19149_),
    .A1(mem_wdata[7]),
    .S(_19180_),
    .X(_03543_));
 sky130_fd_sc_hd__mux2_2 _22467_ (.A0(_19150_),
    .A1(mem_wdata[6]),
    .S(_19180_),
    .X(_03542_));
 sky130_fd_sc_hd__mux2_2 _22468_ (.A0(_19151_),
    .A1(mem_wdata[5]),
    .S(_19180_),
    .X(_03541_));
 sky130_fd_sc_hd__mux2_2 _22469_ (.A0(_19152_),
    .A1(mem_wdata[4]),
    .S(_19180_),
    .X(_03540_));
 sky130_fd_sc_hd__mux2_2 _22470_ (.A0(_19153_),
    .A1(mem_wdata[3]),
    .S(_19180_),
    .X(_03539_));
 sky130_fd_sc_hd__mux2_2 _22471_ (.A0(_19154_),
    .A1(mem_wdata[2]),
    .S(_19180_),
    .X(_03538_));
 sky130_fd_sc_hd__mux2_2 _22472_ (.A0(_19155_),
    .A1(mem_wdata[1]),
    .S(_19175_),
    .X(_03537_));
 sky130_fd_sc_hd__mux2_2 _22473_ (.A0(_19156_),
    .A1(mem_wdata[0]),
    .S(_19175_),
    .X(_03536_));
 sky130_fd_sc_hd__nand2_2 _22474_ (.A(_19164_),
    .B(_19082_),
    .Y(_19181_));
 sky130_fd_sc_hd__buf_1 _22475_ (.A(_19181_),
    .X(_19182_));
 sky130_fd_sc_hd__buf_1 _22476_ (.A(_19182_),
    .X(_19183_));
 sky130_fd_sc_hd__mux2_2 _22477_ (.A0(_19068_),
    .A1(\cpuregs[7][31] ),
    .S(_19183_),
    .X(_03535_));
 sky130_fd_sc_hd__mux2_2 _22478_ (.A0(_19086_),
    .A1(\cpuregs[7][30] ),
    .S(_19183_),
    .X(_03534_));
 sky130_fd_sc_hd__mux2_2 _22479_ (.A0(_19087_),
    .A1(\cpuregs[7][29] ),
    .S(_19183_),
    .X(_03533_));
 sky130_fd_sc_hd__mux2_2 _22480_ (.A0(_19088_),
    .A1(\cpuregs[7][28] ),
    .S(_19183_),
    .X(_03532_));
 sky130_fd_sc_hd__mux2_2 _22481_ (.A0(_19089_),
    .A1(\cpuregs[7][27] ),
    .S(_19183_),
    .X(_03531_));
 sky130_fd_sc_hd__mux2_2 _22482_ (.A0(_19090_),
    .A1(\cpuregs[7][26] ),
    .S(_19183_),
    .X(_03530_));
 sky130_fd_sc_hd__buf_1 _22483_ (.A(_19182_),
    .X(_19184_));
 sky130_fd_sc_hd__mux2_2 _22484_ (.A0(_19091_),
    .A1(\cpuregs[7][25] ),
    .S(_19184_),
    .X(_03529_));
 sky130_fd_sc_hd__mux2_2 _22485_ (.A0(_19093_),
    .A1(\cpuregs[7][24] ),
    .S(_19184_),
    .X(_03528_));
 sky130_fd_sc_hd__mux2_2 _22486_ (.A0(_19094_),
    .A1(\cpuregs[7][23] ),
    .S(_19184_),
    .X(_03527_));
 sky130_fd_sc_hd__mux2_2 _22487_ (.A0(_19095_),
    .A1(\cpuregs[7][22] ),
    .S(_19184_),
    .X(_03526_));
 sky130_fd_sc_hd__mux2_2 _22488_ (.A0(_19096_),
    .A1(\cpuregs[7][21] ),
    .S(_19184_),
    .X(_03525_));
 sky130_fd_sc_hd__mux2_2 _22489_ (.A0(_19097_),
    .A1(\cpuregs[7][20] ),
    .S(_19184_),
    .X(_03524_));
 sky130_fd_sc_hd__buf_1 _22490_ (.A(_19182_),
    .X(_19185_));
 sky130_fd_sc_hd__mux2_2 _22491_ (.A0(_19098_),
    .A1(\cpuregs[7][19] ),
    .S(_19185_),
    .X(_03523_));
 sky130_fd_sc_hd__mux2_2 _22492_ (.A0(_19100_),
    .A1(\cpuregs[7][18] ),
    .S(_19185_),
    .X(_03522_));
 sky130_fd_sc_hd__mux2_2 _22493_ (.A0(_19101_),
    .A1(\cpuregs[7][17] ),
    .S(_19185_),
    .X(_03521_));
 sky130_fd_sc_hd__mux2_2 _22494_ (.A0(_19102_),
    .A1(\cpuregs[7][16] ),
    .S(_19185_),
    .X(_03520_));
 sky130_fd_sc_hd__mux2_2 _22495_ (.A0(_19103_),
    .A1(\cpuregs[7][15] ),
    .S(_19185_),
    .X(_03519_));
 sky130_fd_sc_hd__mux2_2 _22496_ (.A0(_19104_),
    .A1(\cpuregs[7][14] ),
    .S(_19185_),
    .X(_03518_));
 sky130_fd_sc_hd__buf_1 _22497_ (.A(_19182_),
    .X(_19186_));
 sky130_fd_sc_hd__mux2_2 _22498_ (.A0(_19105_),
    .A1(\cpuregs[7][13] ),
    .S(_19186_),
    .X(_03517_));
 sky130_fd_sc_hd__mux2_2 _22499_ (.A0(_19107_),
    .A1(\cpuregs[7][12] ),
    .S(_19186_),
    .X(_03516_));
 sky130_fd_sc_hd__mux2_2 _22500_ (.A0(_19108_),
    .A1(\cpuregs[7][11] ),
    .S(_19186_),
    .X(_03515_));
 sky130_fd_sc_hd__mux2_2 _22501_ (.A0(_19109_),
    .A1(\cpuregs[7][10] ),
    .S(_19186_),
    .X(_03514_));
 sky130_fd_sc_hd__mux2_2 _22502_ (.A0(_19110_),
    .A1(\cpuregs[7][9] ),
    .S(_19186_),
    .X(_03513_));
 sky130_fd_sc_hd__mux2_2 _22503_ (.A0(_19111_),
    .A1(\cpuregs[7][8] ),
    .S(_19186_),
    .X(_03512_));
 sky130_fd_sc_hd__buf_1 _22504_ (.A(_19181_),
    .X(_19187_));
 sky130_fd_sc_hd__mux2_2 _22505_ (.A0(_19112_),
    .A1(\cpuregs[7][7] ),
    .S(_19187_),
    .X(_03511_));
 sky130_fd_sc_hd__mux2_2 _22506_ (.A0(_19114_),
    .A1(\cpuregs[7][6] ),
    .S(_19187_),
    .X(_03510_));
 sky130_fd_sc_hd__mux2_2 _22507_ (.A0(_19115_),
    .A1(\cpuregs[7][5] ),
    .S(_19187_),
    .X(_03509_));
 sky130_fd_sc_hd__mux2_2 _22508_ (.A0(_19116_),
    .A1(\cpuregs[7][4] ),
    .S(_19187_),
    .X(_03508_));
 sky130_fd_sc_hd__mux2_2 _22509_ (.A0(_19117_),
    .A1(\cpuregs[7][3] ),
    .S(_19187_),
    .X(_03507_));
 sky130_fd_sc_hd__mux2_2 _22510_ (.A0(_19118_),
    .A1(\cpuregs[7][2] ),
    .S(_19187_),
    .X(_03506_));
 sky130_fd_sc_hd__mux2_2 _22511_ (.A0(_19119_),
    .A1(\cpuregs[7][1] ),
    .S(_19182_),
    .X(_03505_));
 sky130_fd_sc_hd__mux2_2 _22512_ (.A0(_19120_),
    .A1(\cpuregs[7][0] ),
    .S(_19182_),
    .X(_03504_));
 sky130_fd_sc_hd__buf_1 _22513_ (.A(_18193_),
    .X(_19188_));
 sky130_fd_sc_hd__or2_2 _22514_ (.A(is_beq_bne_blt_bge_bltu_bgeu),
    .B(_18252_),
    .X(_19189_));
 sky130_fd_sc_hd__o2111a_2 _22515_ (.A1(instr_setq),
    .A2(_19188_),
    .B1(_18637_),
    .C1(_18035_),
    .D1(_19189_),
    .X(_19190_));
 sky130_fd_sc_hd__mux2_2 _22516_ (.A0(\latched_rd[4] ),
    .A1(_20583_),
    .S(_19190_),
    .X(_03503_));
 sky130_fd_sc_hd__and3_2 _22517_ (.A(_19081_),
    .B(\latched_rd[2] ),
    .C(\latched_rd[3] ),
    .X(_19191_));
 sky130_fd_sc_hd__nand2_2 _22518_ (.A(_19164_),
    .B(_19191_),
    .Y(_19192_));
 sky130_fd_sc_hd__buf_1 _22519_ (.A(_19192_),
    .X(_19193_));
 sky130_fd_sc_hd__buf_1 _22520_ (.A(_19193_),
    .X(_19194_));
 sky130_fd_sc_hd__mux2_2 _22521_ (.A0(_19068_),
    .A1(\cpuregs[15][31] ),
    .S(_19194_),
    .X(_03502_));
 sky130_fd_sc_hd__mux2_2 _22522_ (.A0(_19086_),
    .A1(\cpuregs[15][30] ),
    .S(_19194_),
    .X(_03501_));
 sky130_fd_sc_hd__mux2_2 _22523_ (.A0(_19087_),
    .A1(\cpuregs[15][29] ),
    .S(_19194_),
    .X(_03500_));
 sky130_fd_sc_hd__mux2_2 _22524_ (.A0(_19088_),
    .A1(\cpuregs[15][28] ),
    .S(_19194_),
    .X(_03499_));
 sky130_fd_sc_hd__mux2_2 _22525_ (.A0(_19089_),
    .A1(\cpuregs[15][27] ),
    .S(_19194_),
    .X(_03498_));
 sky130_fd_sc_hd__mux2_2 _22526_ (.A0(_19090_),
    .A1(\cpuregs[15][26] ),
    .S(_19194_),
    .X(_03497_));
 sky130_fd_sc_hd__buf_1 _22527_ (.A(_19193_),
    .X(_19195_));
 sky130_fd_sc_hd__mux2_2 _22528_ (.A0(_19091_),
    .A1(\cpuregs[15][25] ),
    .S(_19195_),
    .X(_03496_));
 sky130_fd_sc_hd__mux2_2 _22529_ (.A0(_19093_),
    .A1(\cpuregs[15][24] ),
    .S(_19195_),
    .X(_03495_));
 sky130_fd_sc_hd__mux2_2 _22530_ (.A0(_19094_),
    .A1(\cpuregs[15][23] ),
    .S(_19195_),
    .X(_03494_));
 sky130_fd_sc_hd__mux2_2 _22531_ (.A0(_19095_),
    .A1(\cpuregs[15][22] ),
    .S(_19195_),
    .X(_03493_));
 sky130_fd_sc_hd__mux2_2 _22532_ (.A0(_19096_),
    .A1(\cpuregs[15][21] ),
    .S(_19195_),
    .X(_03492_));
 sky130_fd_sc_hd__mux2_2 _22533_ (.A0(_19097_),
    .A1(\cpuregs[15][20] ),
    .S(_19195_),
    .X(_03491_));
 sky130_fd_sc_hd__buf_1 _22534_ (.A(_19193_),
    .X(_19196_));
 sky130_fd_sc_hd__mux2_2 _22535_ (.A0(_19098_),
    .A1(\cpuregs[15][19] ),
    .S(_19196_),
    .X(_03490_));
 sky130_fd_sc_hd__mux2_2 _22536_ (.A0(_19100_),
    .A1(\cpuregs[15][18] ),
    .S(_19196_),
    .X(_03489_));
 sky130_fd_sc_hd__mux2_2 _22537_ (.A0(_19101_),
    .A1(\cpuregs[15][17] ),
    .S(_19196_),
    .X(_03488_));
 sky130_fd_sc_hd__mux2_2 _22538_ (.A0(_19102_),
    .A1(\cpuregs[15][16] ),
    .S(_19196_),
    .X(_03487_));
 sky130_fd_sc_hd__mux2_2 _22539_ (.A0(_19103_),
    .A1(\cpuregs[15][15] ),
    .S(_19196_),
    .X(_03486_));
 sky130_fd_sc_hd__mux2_2 _22540_ (.A0(_19104_),
    .A1(\cpuregs[15][14] ),
    .S(_19196_),
    .X(_03485_));
 sky130_fd_sc_hd__buf_1 _22541_ (.A(_19193_),
    .X(_19197_));
 sky130_fd_sc_hd__mux2_2 _22542_ (.A0(_19105_),
    .A1(\cpuregs[15][13] ),
    .S(_19197_),
    .X(_03484_));
 sky130_fd_sc_hd__mux2_2 _22543_ (.A0(_19107_),
    .A1(\cpuregs[15][12] ),
    .S(_19197_),
    .X(_03483_));
 sky130_fd_sc_hd__mux2_2 _22544_ (.A0(_19108_),
    .A1(\cpuregs[15][11] ),
    .S(_19197_),
    .X(_03482_));
 sky130_fd_sc_hd__mux2_2 _22545_ (.A0(_19109_),
    .A1(\cpuregs[15][10] ),
    .S(_19197_),
    .X(_03481_));
 sky130_fd_sc_hd__mux2_2 _22546_ (.A0(_19110_),
    .A1(\cpuregs[15][9] ),
    .S(_19197_),
    .X(_03480_));
 sky130_fd_sc_hd__mux2_2 _22547_ (.A0(_19111_),
    .A1(\cpuregs[15][8] ),
    .S(_19197_),
    .X(_03479_));
 sky130_fd_sc_hd__buf_1 _22548_ (.A(_19192_),
    .X(_19198_));
 sky130_fd_sc_hd__mux2_2 _22549_ (.A0(_19112_),
    .A1(\cpuregs[15][7] ),
    .S(_19198_),
    .X(_03478_));
 sky130_fd_sc_hd__mux2_2 _22550_ (.A0(_19114_),
    .A1(\cpuregs[15][6] ),
    .S(_19198_),
    .X(_03477_));
 sky130_fd_sc_hd__mux2_2 _22551_ (.A0(_19115_),
    .A1(\cpuregs[15][5] ),
    .S(_19198_),
    .X(_03476_));
 sky130_fd_sc_hd__mux2_2 _22552_ (.A0(_19116_),
    .A1(\cpuregs[15][4] ),
    .S(_19198_),
    .X(_03475_));
 sky130_fd_sc_hd__mux2_2 _22553_ (.A0(_19117_),
    .A1(\cpuregs[15][3] ),
    .S(_19198_),
    .X(_03474_));
 sky130_fd_sc_hd__mux2_2 _22554_ (.A0(_19118_),
    .A1(\cpuregs[15][2] ),
    .S(_19198_),
    .X(_03473_));
 sky130_fd_sc_hd__mux2_2 _22555_ (.A0(_19119_),
    .A1(\cpuregs[15][1] ),
    .S(_19193_),
    .X(_03472_));
 sky130_fd_sc_hd__mux2_2 _22556_ (.A0(_19120_),
    .A1(\cpuregs[15][0] ),
    .S(_19193_),
    .X(_03471_));
 sky130_fd_sc_hd__buf_1 _22557_ (.A(\cpuregs_wrdata[31] ),
    .X(_19199_));
 sky130_fd_sc_hd__nand2_2 _22558_ (.A(_19164_),
    .B(_19123_),
    .Y(_19200_));
 sky130_fd_sc_hd__buf_1 _22559_ (.A(_19200_),
    .X(_19201_));
 sky130_fd_sc_hd__buf_1 _22560_ (.A(_19201_),
    .X(_19202_));
 sky130_fd_sc_hd__mux2_2 _22561_ (.A0(_19199_),
    .A1(\cpuregs[11][31] ),
    .S(_19202_),
    .X(_03470_));
 sky130_fd_sc_hd__buf_1 _22562_ (.A(\cpuregs_wrdata[30] ),
    .X(_19203_));
 sky130_fd_sc_hd__mux2_2 _22563_ (.A0(_19203_),
    .A1(\cpuregs[11][30] ),
    .S(_19202_),
    .X(_03469_));
 sky130_fd_sc_hd__buf_1 _22564_ (.A(\cpuregs_wrdata[29] ),
    .X(_19204_));
 sky130_fd_sc_hd__mux2_2 _22565_ (.A0(_19204_),
    .A1(\cpuregs[11][29] ),
    .S(_19202_),
    .X(_03468_));
 sky130_fd_sc_hd__buf_1 _22566_ (.A(\cpuregs_wrdata[28] ),
    .X(_19205_));
 sky130_fd_sc_hd__mux2_2 _22567_ (.A0(_19205_),
    .A1(\cpuregs[11][28] ),
    .S(_19202_),
    .X(_03467_));
 sky130_fd_sc_hd__buf_1 _22568_ (.A(\cpuregs_wrdata[27] ),
    .X(_19206_));
 sky130_fd_sc_hd__mux2_2 _22569_ (.A0(_19206_),
    .A1(\cpuregs[11][27] ),
    .S(_19202_),
    .X(_03466_));
 sky130_fd_sc_hd__buf_1 _22570_ (.A(\cpuregs_wrdata[26] ),
    .X(_19207_));
 sky130_fd_sc_hd__mux2_2 _22571_ (.A0(_19207_),
    .A1(\cpuregs[11][26] ),
    .S(_19202_),
    .X(_03465_));
 sky130_fd_sc_hd__buf_1 _22572_ (.A(\cpuregs_wrdata[25] ),
    .X(_19208_));
 sky130_fd_sc_hd__buf_1 _22573_ (.A(_19201_),
    .X(_19209_));
 sky130_fd_sc_hd__mux2_2 _22574_ (.A0(_19208_),
    .A1(\cpuregs[11][25] ),
    .S(_19209_),
    .X(_03464_));
 sky130_fd_sc_hd__buf_1 _22575_ (.A(\cpuregs_wrdata[24] ),
    .X(_19210_));
 sky130_fd_sc_hd__mux2_2 _22576_ (.A0(_19210_),
    .A1(\cpuregs[11][24] ),
    .S(_19209_),
    .X(_03463_));
 sky130_fd_sc_hd__buf_1 _22577_ (.A(\cpuregs_wrdata[23] ),
    .X(_19211_));
 sky130_fd_sc_hd__mux2_2 _22578_ (.A0(_19211_),
    .A1(\cpuregs[11][23] ),
    .S(_19209_),
    .X(_03462_));
 sky130_fd_sc_hd__buf_1 _22579_ (.A(\cpuregs_wrdata[22] ),
    .X(_19212_));
 sky130_fd_sc_hd__mux2_2 _22580_ (.A0(_19212_),
    .A1(\cpuregs[11][22] ),
    .S(_19209_),
    .X(_03461_));
 sky130_fd_sc_hd__buf_1 _22581_ (.A(\cpuregs_wrdata[21] ),
    .X(_19213_));
 sky130_fd_sc_hd__mux2_2 _22582_ (.A0(_19213_),
    .A1(\cpuregs[11][21] ),
    .S(_19209_),
    .X(_03460_));
 sky130_fd_sc_hd__buf_1 _22583_ (.A(\cpuregs_wrdata[20] ),
    .X(_19214_));
 sky130_fd_sc_hd__mux2_2 _22584_ (.A0(_19214_),
    .A1(\cpuregs[11][20] ),
    .S(_19209_),
    .X(_03459_));
 sky130_fd_sc_hd__buf_1 _22585_ (.A(\cpuregs_wrdata[19] ),
    .X(_19215_));
 sky130_fd_sc_hd__buf_1 _22586_ (.A(_19201_),
    .X(_19216_));
 sky130_fd_sc_hd__mux2_2 _22587_ (.A0(_19215_),
    .A1(\cpuregs[11][19] ),
    .S(_19216_),
    .X(_03458_));
 sky130_fd_sc_hd__buf_1 _22588_ (.A(\cpuregs_wrdata[18] ),
    .X(_19217_));
 sky130_fd_sc_hd__mux2_2 _22589_ (.A0(_19217_),
    .A1(\cpuregs[11][18] ),
    .S(_19216_),
    .X(_03457_));
 sky130_fd_sc_hd__buf_1 _22590_ (.A(\cpuregs_wrdata[17] ),
    .X(_19218_));
 sky130_fd_sc_hd__mux2_2 _22591_ (.A0(_19218_),
    .A1(\cpuregs[11][17] ),
    .S(_19216_),
    .X(_03456_));
 sky130_fd_sc_hd__buf_1 _22592_ (.A(\cpuregs_wrdata[16] ),
    .X(_19219_));
 sky130_fd_sc_hd__mux2_2 _22593_ (.A0(_19219_),
    .A1(\cpuregs[11][16] ),
    .S(_19216_),
    .X(_03455_));
 sky130_fd_sc_hd__buf_1 _22594_ (.A(\cpuregs_wrdata[15] ),
    .X(_19220_));
 sky130_fd_sc_hd__mux2_2 _22595_ (.A0(_19220_),
    .A1(\cpuregs[11][15] ),
    .S(_19216_),
    .X(_03454_));
 sky130_fd_sc_hd__buf_1 _22596_ (.A(\cpuregs_wrdata[14] ),
    .X(_19221_));
 sky130_fd_sc_hd__mux2_2 _22597_ (.A0(_19221_),
    .A1(\cpuregs[11][14] ),
    .S(_19216_),
    .X(_03453_));
 sky130_fd_sc_hd__buf_1 _22598_ (.A(\cpuregs_wrdata[13] ),
    .X(_19222_));
 sky130_fd_sc_hd__buf_1 _22599_ (.A(_19201_),
    .X(_19223_));
 sky130_fd_sc_hd__mux2_2 _22600_ (.A0(_19222_),
    .A1(\cpuregs[11][13] ),
    .S(_19223_),
    .X(_03452_));
 sky130_fd_sc_hd__buf_1 _22601_ (.A(\cpuregs_wrdata[12] ),
    .X(_19224_));
 sky130_fd_sc_hd__mux2_2 _22602_ (.A0(_19224_),
    .A1(\cpuregs[11][12] ),
    .S(_19223_),
    .X(_03451_));
 sky130_fd_sc_hd__buf_1 _22603_ (.A(\cpuregs_wrdata[11] ),
    .X(_19225_));
 sky130_fd_sc_hd__mux2_2 _22604_ (.A0(_19225_),
    .A1(\cpuregs[11][11] ),
    .S(_19223_),
    .X(_03450_));
 sky130_fd_sc_hd__buf_1 _22605_ (.A(\cpuregs_wrdata[10] ),
    .X(_19226_));
 sky130_fd_sc_hd__mux2_2 _22606_ (.A0(_19226_),
    .A1(\cpuregs[11][10] ),
    .S(_19223_),
    .X(_03449_));
 sky130_fd_sc_hd__buf_1 _22607_ (.A(\cpuregs_wrdata[9] ),
    .X(_19227_));
 sky130_fd_sc_hd__mux2_2 _22608_ (.A0(_19227_),
    .A1(\cpuregs[11][9] ),
    .S(_19223_),
    .X(_03448_));
 sky130_fd_sc_hd__buf_1 _22609_ (.A(\cpuregs_wrdata[8] ),
    .X(_19228_));
 sky130_fd_sc_hd__mux2_2 _22610_ (.A0(_19228_),
    .A1(\cpuregs[11][8] ),
    .S(_19223_),
    .X(_03447_));
 sky130_fd_sc_hd__buf_1 _22611_ (.A(\cpuregs_wrdata[7] ),
    .X(_19229_));
 sky130_fd_sc_hd__buf_1 _22612_ (.A(_19200_),
    .X(_19230_));
 sky130_fd_sc_hd__mux2_2 _22613_ (.A0(_19229_),
    .A1(\cpuregs[11][7] ),
    .S(_19230_),
    .X(_03446_));
 sky130_fd_sc_hd__buf_1 _22614_ (.A(\cpuregs_wrdata[6] ),
    .X(_19231_));
 sky130_fd_sc_hd__mux2_2 _22615_ (.A0(_19231_),
    .A1(\cpuregs[11][6] ),
    .S(_19230_),
    .X(_03445_));
 sky130_fd_sc_hd__buf_1 _22616_ (.A(\cpuregs_wrdata[5] ),
    .X(_19232_));
 sky130_fd_sc_hd__mux2_2 _22617_ (.A0(_19232_),
    .A1(\cpuregs[11][5] ),
    .S(_19230_),
    .X(_03444_));
 sky130_fd_sc_hd__buf_1 _22618_ (.A(\cpuregs_wrdata[4] ),
    .X(_19233_));
 sky130_fd_sc_hd__mux2_2 _22619_ (.A0(_19233_),
    .A1(\cpuregs[11][4] ),
    .S(_19230_),
    .X(_03443_));
 sky130_fd_sc_hd__buf_1 _22620_ (.A(\cpuregs_wrdata[3] ),
    .X(_19234_));
 sky130_fd_sc_hd__mux2_2 _22621_ (.A0(_19234_),
    .A1(\cpuregs[11][3] ),
    .S(_19230_),
    .X(_03442_));
 sky130_fd_sc_hd__buf_1 _22622_ (.A(\cpuregs_wrdata[2] ),
    .X(_19235_));
 sky130_fd_sc_hd__mux2_2 _22623_ (.A0(_19235_),
    .A1(\cpuregs[11][2] ),
    .S(_19230_),
    .X(_03441_));
 sky130_fd_sc_hd__buf_1 _22624_ (.A(\cpuregs_wrdata[1] ),
    .X(_19236_));
 sky130_fd_sc_hd__mux2_2 _22625_ (.A0(_19236_),
    .A1(\cpuregs[11][1] ),
    .S(_19201_),
    .X(_03440_));
 sky130_fd_sc_hd__buf_1 _22626_ (.A(\cpuregs_wrdata[0] ),
    .X(_19237_));
 sky130_fd_sc_hd__mux2_2 _22627_ (.A0(_19237_),
    .A1(\cpuregs[11][0] ),
    .S(_19201_),
    .X(_03439_));
 sky130_fd_sc_hd__inv_2 _22628_ (.A(_19074_),
    .Y(_19238_));
 sky130_fd_sc_hd__nand2_2 _22629_ (.A(_19164_),
    .B(_19238_),
    .Y(_19239_));
 sky130_fd_sc_hd__buf_1 _22630_ (.A(_19239_),
    .X(_19240_));
 sky130_fd_sc_hd__buf_1 _22631_ (.A(_19240_),
    .X(_19241_));
 sky130_fd_sc_hd__mux2_2 _22632_ (.A0(_19199_),
    .A1(\cpuregs[3][31] ),
    .S(_19241_),
    .X(_03438_));
 sky130_fd_sc_hd__mux2_2 _22633_ (.A0(_19203_),
    .A1(\cpuregs[3][30] ),
    .S(_19241_),
    .X(_03437_));
 sky130_fd_sc_hd__mux2_2 _22634_ (.A0(_19204_),
    .A1(\cpuregs[3][29] ),
    .S(_19241_),
    .X(_03436_));
 sky130_fd_sc_hd__mux2_2 _22635_ (.A0(_19205_),
    .A1(\cpuregs[3][28] ),
    .S(_19241_),
    .X(_03435_));
 sky130_fd_sc_hd__mux2_2 _22636_ (.A0(_19206_),
    .A1(\cpuregs[3][27] ),
    .S(_19241_),
    .X(_03434_));
 sky130_fd_sc_hd__mux2_2 _22637_ (.A0(_19207_),
    .A1(\cpuregs[3][26] ),
    .S(_19241_),
    .X(_03433_));
 sky130_fd_sc_hd__buf_1 _22638_ (.A(_19240_),
    .X(_19242_));
 sky130_fd_sc_hd__mux2_2 _22639_ (.A0(_19208_),
    .A1(\cpuregs[3][25] ),
    .S(_19242_),
    .X(_03432_));
 sky130_fd_sc_hd__mux2_2 _22640_ (.A0(_19210_),
    .A1(\cpuregs[3][24] ),
    .S(_19242_),
    .X(_03431_));
 sky130_fd_sc_hd__mux2_2 _22641_ (.A0(_19211_),
    .A1(\cpuregs[3][23] ),
    .S(_19242_),
    .X(_03430_));
 sky130_fd_sc_hd__mux2_2 _22642_ (.A0(_19212_),
    .A1(\cpuregs[3][22] ),
    .S(_19242_),
    .X(_03429_));
 sky130_fd_sc_hd__mux2_2 _22643_ (.A0(_19213_),
    .A1(\cpuregs[3][21] ),
    .S(_19242_),
    .X(_03428_));
 sky130_fd_sc_hd__mux2_2 _22644_ (.A0(_19214_),
    .A1(\cpuregs[3][20] ),
    .S(_19242_),
    .X(_03427_));
 sky130_fd_sc_hd__buf_1 _22645_ (.A(_19240_),
    .X(_19243_));
 sky130_fd_sc_hd__mux2_2 _22646_ (.A0(_19215_),
    .A1(\cpuregs[3][19] ),
    .S(_19243_),
    .X(_03426_));
 sky130_fd_sc_hd__mux2_2 _22647_ (.A0(_19217_),
    .A1(\cpuregs[3][18] ),
    .S(_19243_),
    .X(_03425_));
 sky130_fd_sc_hd__mux2_2 _22648_ (.A0(_19218_),
    .A1(\cpuregs[3][17] ),
    .S(_19243_),
    .X(_03424_));
 sky130_fd_sc_hd__mux2_2 _22649_ (.A0(_19219_),
    .A1(\cpuregs[3][16] ),
    .S(_19243_),
    .X(_03423_));
 sky130_fd_sc_hd__mux2_2 _22650_ (.A0(_19220_),
    .A1(\cpuregs[3][15] ),
    .S(_19243_),
    .X(_03422_));
 sky130_fd_sc_hd__mux2_2 _22651_ (.A0(_19221_),
    .A1(\cpuregs[3][14] ),
    .S(_19243_),
    .X(_03421_));
 sky130_fd_sc_hd__buf_1 _22652_ (.A(_19240_),
    .X(_19244_));
 sky130_fd_sc_hd__mux2_2 _22653_ (.A0(_19222_),
    .A1(\cpuregs[3][13] ),
    .S(_19244_),
    .X(_03420_));
 sky130_fd_sc_hd__mux2_2 _22654_ (.A0(_19224_),
    .A1(\cpuregs[3][12] ),
    .S(_19244_),
    .X(_03419_));
 sky130_fd_sc_hd__mux2_2 _22655_ (.A0(_19225_),
    .A1(\cpuregs[3][11] ),
    .S(_19244_),
    .X(_03418_));
 sky130_fd_sc_hd__mux2_2 _22656_ (.A0(_19226_),
    .A1(\cpuregs[3][10] ),
    .S(_19244_),
    .X(_03417_));
 sky130_fd_sc_hd__mux2_2 _22657_ (.A0(_19227_),
    .A1(\cpuregs[3][9] ),
    .S(_19244_),
    .X(_03416_));
 sky130_fd_sc_hd__mux2_2 _22658_ (.A0(_19228_),
    .A1(\cpuregs[3][8] ),
    .S(_19244_),
    .X(_03415_));
 sky130_fd_sc_hd__buf_1 _22659_ (.A(_19239_),
    .X(_19245_));
 sky130_fd_sc_hd__mux2_2 _22660_ (.A0(_19229_),
    .A1(\cpuregs[3][7] ),
    .S(_19245_),
    .X(_03414_));
 sky130_fd_sc_hd__mux2_2 _22661_ (.A0(_19231_),
    .A1(\cpuregs[3][6] ),
    .S(_19245_),
    .X(_03413_));
 sky130_fd_sc_hd__mux2_2 _22662_ (.A0(_19232_),
    .A1(\cpuregs[3][5] ),
    .S(_19245_),
    .X(_03412_));
 sky130_fd_sc_hd__mux2_2 _22663_ (.A0(_19233_),
    .A1(\cpuregs[3][4] ),
    .S(_19245_),
    .X(_03411_));
 sky130_fd_sc_hd__mux2_2 _22664_ (.A0(_19234_),
    .A1(\cpuregs[3][3] ),
    .S(_19245_),
    .X(_03410_));
 sky130_fd_sc_hd__mux2_2 _22665_ (.A0(_19235_),
    .A1(\cpuregs[3][2] ),
    .S(_19245_),
    .X(_03409_));
 sky130_fd_sc_hd__mux2_2 _22666_ (.A0(_19236_),
    .A1(\cpuregs[3][1] ),
    .S(_19240_),
    .X(_03408_));
 sky130_fd_sc_hd__mux2_2 _22667_ (.A0(_19237_),
    .A1(\cpuregs[3][0] ),
    .S(_19240_),
    .X(_03407_));
 sky130_fd_sc_hd__buf_1 _22668_ (.A(\cpuregs_wrdata[31] ),
    .X(_19246_));
 sky130_fd_sc_hd__and2_2 _22669_ (.A(_19121_),
    .B(_19238_),
    .X(_19247_));
 sky130_fd_sc_hd__buf_1 _22670_ (.A(_19247_),
    .X(_19248_));
 sky130_fd_sc_hd__buf_1 _22671_ (.A(_19248_),
    .X(_19249_));
 sky130_fd_sc_hd__mux2_2 _22672_ (.A0(\cpuregs[1][31] ),
    .A1(_19246_),
    .S(_19249_),
    .X(_03406_));
 sky130_fd_sc_hd__buf_1 _22673_ (.A(\cpuregs_wrdata[30] ),
    .X(_19250_));
 sky130_fd_sc_hd__mux2_2 _22674_ (.A0(\cpuregs[1][30] ),
    .A1(_19250_),
    .S(_19249_),
    .X(_03405_));
 sky130_fd_sc_hd__buf_1 _22675_ (.A(\cpuregs_wrdata[29] ),
    .X(_19251_));
 sky130_fd_sc_hd__mux2_2 _22676_ (.A0(\cpuregs[1][29] ),
    .A1(_19251_),
    .S(_19249_),
    .X(_03404_));
 sky130_fd_sc_hd__buf_1 _22677_ (.A(\cpuregs_wrdata[28] ),
    .X(_19252_));
 sky130_fd_sc_hd__mux2_2 _22678_ (.A0(\cpuregs[1][28] ),
    .A1(_19252_),
    .S(_19249_),
    .X(_03403_));
 sky130_fd_sc_hd__buf_1 _22679_ (.A(\cpuregs_wrdata[27] ),
    .X(_19253_));
 sky130_fd_sc_hd__mux2_2 _22680_ (.A0(\cpuregs[1][27] ),
    .A1(_19253_),
    .S(_19249_),
    .X(_03402_));
 sky130_fd_sc_hd__buf_1 _22681_ (.A(\cpuregs_wrdata[26] ),
    .X(_19254_));
 sky130_fd_sc_hd__mux2_2 _22682_ (.A0(\cpuregs[1][26] ),
    .A1(_19254_),
    .S(_19249_),
    .X(_03401_));
 sky130_fd_sc_hd__buf_1 _22683_ (.A(\cpuregs_wrdata[25] ),
    .X(_19255_));
 sky130_fd_sc_hd__buf_1 _22684_ (.A(_19248_),
    .X(_19256_));
 sky130_fd_sc_hd__mux2_2 _22685_ (.A0(\cpuregs[1][25] ),
    .A1(_19255_),
    .S(_19256_),
    .X(_03400_));
 sky130_fd_sc_hd__buf_1 _22686_ (.A(\cpuregs_wrdata[24] ),
    .X(_19257_));
 sky130_fd_sc_hd__mux2_2 _22687_ (.A0(\cpuregs[1][24] ),
    .A1(_19257_),
    .S(_19256_),
    .X(_03399_));
 sky130_fd_sc_hd__buf_1 _22688_ (.A(\cpuregs_wrdata[23] ),
    .X(_19258_));
 sky130_fd_sc_hd__mux2_2 _22689_ (.A0(\cpuregs[1][23] ),
    .A1(_19258_),
    .S(_19256_),
    .X(_03398_));
 sky130_fd_sc_hd__buf_1 _22690_ (.A(\cpuregs_wrdata[22] ),
    .X(_19259_));
 sky130_fd_sc_hd__mux2_2 _22691_ (.A0(\cpuregs[1][22] ),
    .A1(_19259_),
    .S(_19256_),
    .X(_03397_));
 sky130_fd_sc_hd__buf_1 _22692_ (.A(\cpuregs_wrdata[21] ),
    .X(_19260_));
 sky130_fd_sc_hd__mux2_2 _22693_ (.A0(\cpuregs[1][21] ),
    .A1(_19260_),
    .S(_19256_),
    .X(_03396_));
 sky130_fd_sc_hd__buf_1 _22694_ (.A(\cpuregs_wrdata[20] ),
    .X(_19261_));
 sky130_fd_sc_hd__mux2_2 _22695_ (.A0(\cpuregs[1][20] ),
    .A1(_19261_),
    .S(_19256_),
    .X(_03395_));
 sky130_fd_sc_hd__buf_1 _22696_ (.A(\cpuregs_wrdata[19] ),
    .X(_19262_));
 sky130_fd_sc_hd__buf_1 _22697_ (.A(_19248_),
    .X(_19263_));
 sky130_fd_sc_hd__mux2_2 _22698_ (.A0(\cpuregs[1][19] ),
    .A1(_19262_),
    .S(_19263_),
    .X(_03394_));
 sky130_fd_sc_hd__buf_1 _22699_ (.A(\cpuregs_wrdata[18] ),
    .X(_19264_));
 sky130_fd_sc_hd__mux2_2 _22700_ (.A0(\cpuregs[1][18] ),
    .A1(_19264_),
    .S(_19263_),
    .X(_03393_));
 sky130_fd_sc_hd__buf_1 _22701_ (.A(\cpuregs_wrdata[17] ),
    .X(_19265_));
 sky130_fd_sc_hd__mux2_2 _22702_ (.A0(\cpuregs[1][17] ),
    .A1(_19265_),
    .S(_19263_),
    .X(_03392_));
 sky130_fd_sc_hd__buf_1 _22703_ (.A(\cpuregs_wrdata[16] ),
    .X(_19266_));
 sky130_fd_sc_hd__mux2_2 _22704_ (.A0(\cpuregs[1][16] ),
    .A1(_19266_),
    .S(_19263_),
    .X(_03391_));
 sky130_fd_sc_hd__buf_1 _22705_ (.A(\cpuregs_wrdata[15] ),
    .X(_19267_));
 sky130_fd_sc_hd__mux2_2 _22706_ (.A0(\cpuregs[1][15] ),
    .A1(_19267_),
    .S(_19263_),
    .X(_03390_));
 sky130_fd_sc_hd__buf_1 _22707_ (.A(\cpuregs_wrdata[14] ),
    .X(_19268_));
 sky130_fd_sc_hd__mux2_2 _22708_ (.A0(\cpuregs[1][14] ),
    .A1(_19268_),
    .S(_19263_),
    .X(_03389_));
 sky130_fd_sc_hd__buf_1 _22709_ (.A(\cpuregs_wrdata[13] ),
    .X(_19269_));
 sky130_fd_sc_hd__buf_1 _22710_ (.A(_19248_),
    .X(_19270_));
 sky130_fd_sc_hd__mux2_2 _22711_ (.A0(\cpuregs[1][13] ),
    .A1(_19269_),
    .S(_19270_),
    .X(_03388_));
 sky130_fd_sc_hd__buf_1 _22712_ (.A(\cpuregs_wrdata[12] ),
    .X(_19271_));
 sky130_fd_sc_hd__mux2_2 _22713_ (.A0(\cpuregs[1][12] ),
    .A1(_19271_),
    .S(_19270_),
    .X(_03387_));
 sky130_fd_sc_hd__buf_1 _22714_ (.A(\cpuregs_wrdata[11] ),
    .X(_19272_));
 sky130_fd_sc_hd__mux2_2 _22715_ (.A0(\cpuregs[1][11] ),
    .A1(_19272_),
    .S(_19270_),
    .X(_03386_));
 sky130_fd_sc_hd__buf_1 _22716_ (.A(\cpuregs_wrdata[10] ),
    .X(_19273_));
 sky130_fd_sc_hd__mux2_2 _22717_ (.A0(\cpuregs[1][10] ),
    .A1(_19273_),
    .S(_19270_),
    .X(_03385_));
 sky130_fd_sc_hd__buf_1 _22718_ (.A(\cpuregs_wrdata[9] ),
    .X(_19274_));
 sky130_fd_sc_hd__mux2_2 _22719_ (.A0(\cpuregs[1][9] ),
    .A1(_19274_),
    .S(_19270_),
    .X(_03384_));
 sky130_fd_sc_hd__buf_1 _22720_ (.A(\cpuregs_wrdata[8] ),
    .X(_19275_));
 sky130_fd_sc_hd__mux2_2 _22721_ (.A0(\cpuregs[1][8] ),
    .A1(_19275_),
    .S(_19270_),
    .X(_03383_));
 sky130_fd_sc_hd__buf_1 _22722_ (.A(\cpuregs_wrdata[7] ),
    .X(_19276_));
 sky130_fd_sc_hd__buf_1 _22723_ (.A(_19247_),
    .X(_19277_));
 sky130_fd_sc_hd__mux2_2 _22724_ (.A0(\cpuregs[1][7] ),
    .A1(_19276_),
    .S(_19277_),
    .X(_03382_));
 sky130_fd_sc_hd__buf_1 _22725_ (.A(\cpuregs_wrdata[6] ),
    .X(_19278_));
 sky130_fd_sc_hd__mux2_2 _22726_ (.A0(\cpuregs[1][6] ),
    .A1(_19278_),
    .S(_19277_),
    .X(_03381_));
 sky130_fd_sc_hd__buf_1 _22727_ (.A(\cpuregs_wrdata[5] ),
    .X(_19279_));
 sky130_fd_sc_hd__mux2_2 _22728_ (.A0(\cpuregs[1][5] ),
    .A1(_19279_),
    .S(_19277_),
    .X(_03380_));
 sky130_fd_sc_hd__buf_1 _22729_ (.A(\cpuregs_wrdata[4] ),
    .X(_19280_));
 sky130_fd_sc_hd__mux2_2 _22730_ (.A0(\cpuregs[1][4] ),
    .A1(_19280_),
    .S(_19277_),
    .X(_03379_));
 sky130_fd_sc_hd__buf_1 _22731_ (.A(\cpuregs_wrdata[3] ),
    .X(_19281_));
 sky130_fd_sc_hd__mux2_2 _22732_ (.A0(\cpuregs[1][3] ),
    .A1(_19281_),
    .S(_19277_),
    .X(_03378_));
 sky130_fd_sc_hd__buf_1 _22733_ (.A(\cpuregs_wrdata[2] ),
    .X(_19282_));
 sky130_fd_sc_hd__mux2_2 _22734_ (.A0(\cpuregs[1][2] ),
    .A1(_19282_),
    .S(_19277_),
    .X(_03377_));
 sky130_fd_sc_hd__buf_1 _22735_ (.A(\cpuregs_wrdata[1] ),
    .X(_19283_));
 sky130_fd_sc_hd__mux2_2 _22736_ (.A0(\cpuregs[1][1] ),
    .A1(_19283_),
    .S(_19248_),
    .X(_03376_));
 sky130_fd_sc_hd__buf_1 _22737_ (.A(\cpuregs_wrdata[0] ),
    .X(_19284_));
 sky130_fd_sc_hd__mux2_2 _22738_ (.A0(\cpuregs[1][0] ),
    .A1(_19284_),
    .S(_19248_),
    .X(_03375_));
 sky130_fd_sc_hd__or3b_2 _22739_ (.A(_19071_),
    .B(_19078_),
    .C_N(_19191_),
    .X(_19285_));
 sky130_fd_sc_hd__buf_1 _22740_ (.A(_19285_),
    .X(_19286_));
 sky130_fd_sc_hd__buf_1 _22741_ (.A(_19286_),
    .X(_19287_));
 sky130_fd_sc_hd__mux2_2 _22742_ (.A0(_19199_),
    .A1(\cpuregs[12][31] ),
    .S(_19287_),
    .X(_03374_));
 sky130_fd_sc_hd__mux2_2 _22743_ (.A0(_19203_),
    .A1(\cpuregs[12][30] ),
    .S(_19287_),
    .X(_03373_));
 sky130_fd_sc_hd__mux2_2 _22744_ (.A0(_19204_),
    .A1(\cpuregs[12][29] ),
    .S(_19287_),
    .X(_03372_));
 sky130_fd_sc_hd__mux2_2 _22745_ (.A0(_19205_),
    .A1(\cpuregs[12][28] ),
    .S(_19287_),
    .X(_03371_));
 sky130_fd_sc_hd__mux2_2 _22746_ (.A0(_19206_),
    .A1(\cpuregs[12][27] ),
    .S(_19287_),
    .X(_03370_));
 sky130_fd_sc_hd__mux2_2 _22747_ (.A0(_19207_),
    .A1(\cpuregs[12][26] ),
    .S(_19287_),
    .X(_03369_));
 sky130_fd_sc_hd__buf_1 _22748_ (.A(_19286_),
    .X(_19288_));
 sky130_fd_sc_hd__mux2_2 _22749_ (.A0(_19208_),
    .A1(\cpuregs[12][25] ),
    .S(_19288_),
    .X(_03368_));
 sky130_fd_sc_hd__mux2_2 _22750_ (.A0(_19210_),
    .A1(\cpuregs[12][24] ),
    .S(_19288_),
    .X(_03367_));
 sky130_fd_sc_hd__mux2_2 _22751_ (.A0(_19211_),
    .A1(\cpuregs[12][23] ),
    .S(_19288_),
    .X(_03366_));
 sky130_fd_sc_hd__mux2_2 _22752_ (.A0(_19212_),
    .A1(\cpuregs[12][22] ),
    .S(_19288_),
    .X(_03365_));
 sky130_fd_sc_hd__mux2_2 _22753_ (.A0(_19213_),
    .A1(\cpuregs[12][21] ),
    .S(_19288_),
    .X(_03364_));
 sky130_fd_sc_hd__mux2_2 _22754_ (.A0(_19214_),
    .A1(\cpuregs[12][20] ),
    .S(_19288_),
    .X(_03363_));
 sky130_fd_sc_hd__buf_1 _22755_ (.A(_19286_),
    .X(_19289_));
 sky130_fd_sc_hd__mux2_2 _22756_ (.A0(_19215_),
    .A1(\cpuregs[12][19] ),
    .S(_19289_),
    .X(_03362_));
 sky130_fd_sc_hd__mux2_2 _22757_ (.A0(_19217_),
    .A1(\cpuregs[12][18] ),
    .S(_19289_),
    .X(_03361_));
 sky130_fd_sc_hd__mux2_2 _22758_ (.A0(_19218_),
    .A1(\cpuregs[12][17] ),
    .S(_19289_),
    .X(_03360_));
 sky130_fd_sc_hd__mux2_2 _22759_ (.A0(_19219_),
    .A1(\cpuregs[12][16] ),
    .S(_19289_),
    .X(_03359_));
 sky130_fd_sc_hd__mux2_2 _22760_ (.A0(_19220_),
    .A1(\cpuregs[12][15] ),
    .S(_19289_),
    .X(_03358_));
 sky130_fd_sc_hd__mux2_2 _22761_ (.A0(_19221_),
    .A1(\cpuregs[12][14] ),
    .S(_19289_),
    .X(_03357_));
 sky130_fd_sc_hd__buf_1 _22762_ (.A(_19286_),
    .X(_19290_));
 sky130_fd_sc_hd__mux2_2 _22763_ (.A0(_19222_),
    .A1(\cpuregs[12][13] ),
    .S(_19290_),
    .X(_03356_));
 sky130_fd_sc_hd__mux2_2 _22764_ (.A0(_19224_),
    .A1(\cpuregs[12][12] ),
    .S(_19290_),
    .X(_03355_));
 sky130_fd_sc_hd__mux2_2 _22765_ (.A0(_19225_),
    .A1(\cpuregs[12][11] ),
    .S(_19290_),
    .X(_03354_));
 sky130_fd_sc_hd__mux2_2 _22766_ (.A0(_19226_),
    .A1(\cpuregs[12][10] ),
    .S(_19290_),
    .X(_03353_));
 sky130_fd_sc_hd__mux2_2 _22767_ (.A0(_19227_),
    .A1(\cpuregs[12][9] ),
    .S(_19290_),
    .X(_03352_));
 sky130_fd_sc_hd__mux2_2 _22768_ (.A0(_19228_),
    .A1(\cpuregs[12][8] ),
    .S(_19290_),
    .X(_03351_));
 sky130_fd_sc_hd__buf_1 _22769_ (.A(_19285_),
    .X(_19291_));
 sky130_fd_sc_hd__mux2_2 _22770_ (.A0(_19229_),
    .A1(\cpuregs[12][7] ),
    .S(_19291_),
    .X(_03350_));
 sky130_fd_sc_hd__mux2_2 _22771_ (.A0(_19231_),
    .A1(\cpuregs[12][6] ),
    .S(_19291_),
    .X(_03349_));
 sky130_fd_sc_hd__mux2_2 _22772_ (.A0(_19232_),
    .A1(\cpuregs[12][5] ),
    .S(_19291_),
    .X(_03348_));
 sky130_fd_sc_hd__mux2_2 _22773_ (.A0(_19233_),
    .A1(\cpuregs[12][4] ),
    .S(_19291_),
    .X(_03347_));
 sky130_fd_sc_hd__mux2_2 _22774_ (.A0(_19234_),
    .A1(\cpuregs[12][3] ),
    .S(_19291_),
    .X(_03346_));
 sky130_fd_sc_hd__mux2_2 _22775_ (.A0(_19235_),
    .A1(\cpuregs[12][2] ),
    .S(_19291_),
    .X(_03345_));
 sky130_fd_sc_hd__mux2_2 _22776_ (.A0(_19236_),
    .A1(\cpuregs[12][1] ),
    .S(_19286_),
    .X(_03344_));
 sky130_fd_sc_hd__mux2_2 _22777_ (.A0(_19237_),
    .A1(\cpuregs[12][0] ),
    .S(_19286_),
    .X(_03343_));
 sky130_fd_sc_hd__or3_2 _22778_ (.A(\latched_rd[2] ),
    .B(\latched_rd[3] ),
    .C(_19071_),
    .X(_19292_));
 sky130_fd_sc_hd__nor2_2 _22779_ (.A(_19292_),
    .B(_19078_),
    .Y(_19293_));
 sky130_fd_sc_hd__buf_1 _22780_ (.A(_19293_),
    .X(_19294_));
 sky130_fd_sc_hd__buf_1 _22781_ (.A(_19294_),
    .X(_19295_));
 sky130_fd_sc_hd__mux2_2 _22782_ (.A0(\cpuregs[16][31] ),
    .A1(_19246_),
    .S(_19295_),
    .X(_03342_));
 sky130_fd_sc_hd__mux2_2 _22783_ (.A0(\cpuregs[16][30] ),
    .A1(_19250_),
    .S(_19295_),
    .X(_03341_));
 sky130_fd_sc_hd__mux2_2 _22784_ (.A0(\cpuregs[16][29] ),
    .A1(_19251_),
    .S(_19295_),
    .X(_03340_));
 sky130_fd_sc_hd__mux2_2 _22785_ (.A0(\cpuregs[16][28] ),
    .A1(_19252_),
    .S(_19295_),
    .X(_03339_));
 sky130_fd_sc_hd__mux2_2 _22786_ (.A0(\cpuregs[16][27] ),
    .A1(_19253_),
    .S(_19295_),
    .X(_03338_));
 sky130_fd_sc_hd__mux2_2 _22787_ (.A0(\cpuregs[16][26] ),
    .A1(_19254_),
    .S(_19295_),
    .X(_03337_));
 sky130_fd_sc_hd__buf_1 _22788_ (.A(_19294_),
    .X(_19296_));
 sky130_fd_sc_hd__mux2_2 _22789_ (.A0(\cpuregs[16][25] ),
    .A1(_19255_),
    .S(_19296_),
    .X(_03336_));
 sky130_fd_sc_hd__mux2_2 _22790_ (.A0(\cpuregs[16][24] ),
    .A1(_19257_),
    .S(_19296_),
    .X(_03335_));
 sky130_fd_sc_hd__mux2_2 _22791_ (.A0(\cpuregs[16][23] ),
    .A1(_19258_),
    .S(_19296_),
    .X(_03334_));
 sky130_fd_sc_hd__mux2_2 _22792_ (.A0(\cpuregs[16][22] ),
    .A1(_19259_),
    .S(_19296_),
    .X(_03333_));
 sky130_fd_sc_hd__mux2_2 _22793_ (.A0(\cpuregs[16][21] ),
    .A1(_19260_),
    .S(_19296_),
    .X(_03332_));
 sky130_fd_sc_hd__mux2_2 _22794_ (.A0(\cpuregs[16][20] ),
    .A1(_19261_),
    .S(_19296_),
    .X(_03331_));
 sky130_fd_sc_hd__buf_1 _22795_ (.A(_19294_),
    .X(_19297_));
 sky130_fd_sc_hd__mux2_2 _22796_ (.A0(\cpuregs[16][19] ),
    .A1(_19262_),
    .S(_19297_),
    .X(_03330_));
 sky130_fd_sc_hd__mux2_2 _22797_ (.A0(\cpuregs[16][18] ),
    .A1(_19264_),
    .S(_19297_),
    .X(_03329_));
 sky130_fd_sc_hd__mux2_2 _22798_ (.A0(\cpuregs[16][17] ),
    .A1(_19265_),
    .S(_19297_),
    .X(_03328_));
 sky130_fd_sc_hd__mux2_2 _22799_ (.A0(\cpuregs[16][16] ),
    .A1(_19266_),
    .S(_19297_),
    .X(_03327_));
 sky130_fd_sc_hd__mux2_2 _22800_ (.A0(\cpuregs[16][15] ),
    .A1(_19267_),
    .S(_19297_),
    .X(_03326_));
 sky130_fd_sc_hd__mux2_2 _22801_ (.A0(\cpuregs[16][14] ),
    .A1(_19268_),
    .S(_19297_),
    .X(_03325_));
 sky130_fd_sc_hd__buf_1 _22802_ (.A(_19294_),
    .X(_19298_));
 sky130_fd_sc_hd__mux2_2 _22803_ (.A0(\cpuregs[16][13] ),
    .A1(_19269_),
    .S(_19298_),
    .X(_03324_));
 sky130_fd_sc_hd__mux2_2 _22804_ (.A0(\cpuregs[16][12] ),
    .A1(_19271_),
    .S(_19298_),
    .X(_03323_));
 sky130_fd_sc_hd__mux2_2 _22805_ (.A0(\cpuregs[16][11] ),
    .A1(_19272_),
    .S(_19298_),
    .X(_03322_));
 sky130_fd_sc_hd__mux2_2 _22806_ (.A0(\cpuregs[16][10] ),
    .A1(_19273_),
    .S(_19298_),
    .X(_03321_));
 sky130_fd_sc_hd__mux2_2 _22807_ (.A0(\cpuregs[16][9] ),
    .A1(_19274_),
    .S(_19298_),
    .X(_03320_));
 sky130_fd_sc_hd__mux2_2 _22808_ (.A0(\cpuregs[16][8] ),
    .A1(_19275_),
    .S(_19298_),
    .X(_03319_));
 sky130_fd_sc_hd__buf_1 _22809_ (.A(_19293_),
    .X(_19299_));
 sky130_fd_sc_hd__mux2_2 _22810_ (.A0(\cpuregs[16][7] ),
    .A1(_19276_),
    .S(_19299_),
    .X(_03318_));
 sky130_fd_sc_hd__mux2_2 _22811_ (.A0(\cpuregs[16][6] ),
    .A1(_19278_),
    .S(_19299_),
    .X(_03317_));
 sky130_fd_sc_hd__mux2_2 _22812_ (.A0(\cpuregs[16][5] ),
    .A1(_19279_),
    .S(_19299_),
    .X(_03316_));
 sky130_fd_sc_hd__mux2_2 _22813_ (.A0(\cpuregs[16][4] ),
    .A1(_19280_),
    .S(_19299_),
    .X(_03315_));
 sky130_fd_sc_hd__mux2_2 _22814_ (.A0(\cpuregs[16][3] ),
    .A1(_19281_),
    .S(_19299_),
    .X(_03314_));
 sky130_fd_sc_hd__mux2_2 _22815_ (.A0(\cpuregs[16][2] ),
    .A1(_19282_),
    .S(_19299_),
    .X(_03313_));
 sky130_fd_sc_hd__mux2_2 _22816_ (.A0(\cpuregs[16][1] ),
    .A1(_19283_),
    .S(_19294_),
    .X(_03312_));
 sky130_fd_sc_hd__mux2_2 _22817_ (.A0(\cpuregs[16][0] ),
    .A1(_19284_),
    .S(_19294_),
    .X(_03311_));
 sky130_fd_sc_hd__and2_2 _22818_ (.A(_19121_),
    .B(_19165_),
    .X(_19300_));
 sky130_fd_sc_hd__buf_1 _22819_ (.A(_19300_),
    .X(_19301_));
 sky130_fd_sc_hd__buf_1 _22820_ (.A(_19301_),
    .X(_19302_));
 sky130_fd_sc_hd__mux2_2 _22821_ (.A0(\cpuregs[17][31] ),
    .A1(_19246_),
    .S(_19302_),
    .X(_03310_));
 sky130_fd_sc_hd__mux2_2 _22822_ (.A0(\cpuregs[17][30] ),
    .A1(_19250_),
    .S(_19302_),
    .X(_03309_));
 sky130_fd_sc_hd__mux2_2 _22823_ (.A0(\cpuregs[17][29] ),
    .A1(_19251_),
    .S(_19302_),
    .X(_03308_));
 sky130_fd_sc_hd__mux2_2 _22824_ (.A0(\cpuregs[17][28] ),
    .A1(_19252_),
    .S(_19302_),
    .X(_03307_));
 sky130_fd_sc_hd__mux2_2 _22825_ (.A0(\cpuregs[17][27] ),
    .A1(_19253_),
    .S(_19302_),
    .X(_03306_));
 sky130_fd_sc_hd__mux2_2 _22826_ (.A0(\cpuregs[17][26] ),
    .A1(_19254_),
    .S(_19302_),
    .X(_03305_));
 sky130_fd_sc_hd__buf_1 _22827_ (.A(_19301_),
    .X(_19303_));
 sky130_fd_sc_hd__mux2_2 _22828_ (.A0(\cpuregs[17][25] ),
    .A1(_19255_),
    .S(_19303_),
    .X(_03304_));
 sky130_fd_sc_hd__mux2_2 _22829_ (.A0(\cpuregs[17][24] ),
    .A1(_19257_),
    .S(_19303_),
    .X(_03303_));
 sky130_fd_sc_hd__mux2_2 _22830_ (.A0(\cpuregs[17][23] ),
    .A1(_19258_),
    .S(_19303_),
    .X(_03302_));
 sky130_fd_sc_hd__mux2_2 _22831_ (.A0(\cpuregs[17][22] ),
    .A1(_19259_),
    .S(_19303_),
    .X(_03301_));
 sky130_fd_sc_hd__mux2_2 _22832_ (.A0(\cpuregs[17][21] ),
    .A1(_19260_),
    .S(_19303_),
    .X(_03300_));
 sky130_fd_sc_hd__mux2_2 _22833_ (.A0(\cpuregs[17][20] ),
    .A1(_19261_),
    .S(_19303_),
    .X(_03299_));
 sky130_fd_sc_hd__buf_1 _22834_ (.A(_19301_),
    .X(_19304_));
 sky130_fd_sc_hd__mux2_2 _22835_ (.A0(\cpuregs[17][19] ),
    .A1(_19262_),
    .S(_19304_),
    .X(_03298_));
 sky130_fd_sc_hd__mux2_2 _22836_ (.A0(\cpuregs[17][18] ),
    .A1(_19264_),
    .S(_19304_),
    .X(_03297_));
 sky130_fd_sc_hd__mux2_2 _22837_ (.A0(\cpuregs[17][17] ),
    .A1(_19265_),
    .S(_19304_),
    .X(_03296_));
 sky130_fd_sc_hd__mux2_2 _22838_ (.A0(\cpuregs[17][16] ),
    .A1(_19266_),
    .S(_19304_),
    .X(_03295_));
 sky130_fd_sc_hd__mux2_2 _22839_ (.A0(\cpuregs[17][15] ),
    .A1(_19267_),
    .S(_19304_),
    .X(_03294_));
 sky130_fd_sc_hd__mux2_2 _22840_ (.A0(\cpuregs[17][14] ),
    .A1(_19268_),
    .S(_19304_),
    .X(_03293_));
 sky130_fd_sc_hd__buf_1 _22841_ (.A(_19301_),
    .X(_19305_));
 sky130_fd_sc_hd__mux2_2 _22842_ (.A0(\cpuregs[17][13] ),
    .A1(_19269_),
    .S(_19305_),
    .X(_03292_));
 sky130_fd_sc_hd__mux2_2 _22843_ (.A0(\cpuregs[17][12] ),
    .A1(_19271_),
    .S(_19305_),
    .X(_03291_));
 sky130_fd_sc_hd__mux2_2 _22844_ (.A0(\cpuregs[17][11] ),
    .A1(_19272_),
    .S(_19305_),
    .X(_03290_));
 sky130_fd_sc_hd__mux2_2 _22845_ (.A0(\cpuregs[17][10] ),
    .A1(_19273_),
    .S(_19305_),
    .X(_03289_));
 sky130_fd_sc_hd__mux2_2 _22846_ (.A0(\cpuregs[17][9] ),
    .A1(_19274_),
    .S(_19305_),
    .X(_03288_));
 sky130_fd_sc_hd__mux2_2 _22847_ (.A0(\cpuregs[17][8] ),
    .A1(_19275_),
    .S(_19305_),
    .X(_03287_));
 sky130_fd_sc_hd__buf_1 _22848_ (.A(_19300_),
    .X(_19306_));
 sky130_fd_sc_hd__mux2_2 _22849_ (.A0(\cpuregs[17][7] ),
    .A1(_19276_),
    .S(_19306_),
    .X(_03286_));
 sky130_fd_sc_hd__mux2_2 _22850_ (.A0(\cpuregs[17][6] ),
    .A1(_19278_),
    .S(_19306_),
    .X(_03285_));
 sky130_fd_sc_hd__mux2_2 _22851_ (.A0(\cpuregs[17][5] ),
    .A1(_19279_),
    .S(_19306_),
    .X(_03284_));
 sky130_fd_sc_hd__mux2_2 _22852_ (.A0(\cpuregs[17][4] ),
    .A1(_19280_),
    .S(_19306_),
    .X(_03283_));
 sky130_fd_sc_hd__mux2_2 _22853_ (.A0(\cpuregs[17][3] ),
    .A1(_19281_),
    .S(_19306_),
    .X(_03282_));
 sky130_fd_sc_hd__mux2_2 _22854_ (.A0(\cpuregs[17][2] ),
    .A1(_19282_),
    .S(_19306_),
    .X(_03281_));
 sky130_fd_sc_hd__mux2_2 _22855_ (.A0(\cpuregs[17][1] ),
    .A1(_19283_),
    .S(_19301_),
    .X(_03280_));
 sky130_fd_sc_hd__mux2_2 _22856_ (.A0(\cpuregs[17][0] ),
    .A1(_19284_),
    .S(_19301_),
    .X(_03279_));
 sky130_fd_sc_hd__buf_1 _22857_ (.A(\pcpi_mul.rs2[31] ),
    .X(_19307_));
 sky130_fd_sc_hd__buf_1 _22858_ (.A(_19307_),
    .X(_19308_));
 sky130_fd_sc_hd__buf_1 _22859_ (.A(_19308_),
    .X(_19309_));
 sky130_fd_sc_hd__buf_1 _22860_ (.A(_19309_),
    .X(_19310_));
 sky130_fd_sc_hd__mux2_2 _22861_ (.A0(pcpi_rs2[31]),
    .A1(_19310_),
    .S(_18172_),
    .X(_03278_));
 sky130_fd_sc_hd__buf_1 _22862_ (.A(\pcpi_mul.rs2[30] ),
    .X(_19311_));
 sky130_fd_sc_hd__buf_1 _22863_ (.A(_19311_),
    .X(_19312_));
 sky130_fd_sc_hd__buf_1 _22864_ (.A(_19312_),
    .X(_19313_));
 sky130_fd_sc_hd__buf_1 _22865_ (.A(_19313_),
    .X(_19314_));
 sky130_fd_sc_hd__mux2_2 _22866_ (.A0(pcpi_rs2[30]),
    .A1(_19314_),
    .S(_18172_),
    .X(_03277_));
 sky130_fd_sc_hd__buf_1 _22867_ (.A(\pcpi_mul.rs2[29] ),
    .X(_19315_));
 sky130_fd_sc_hd__buf_1 _22868_ (.A(_19315_),
    .X(_19316_));
 sky130_fd_sc_hd__buf_1 _22869_ (.A(_19316_),
    .X(_19317_));
 sky130_fd_sc_hd__buf_1 _22870_ (.A(_19317_),
    .X(_19318_));
 sky130_fd_sc_hd__mux2_2 _22871_ (.A0(_19134_),
    .A1(_19318_),
    .S(_18172_),
    .X(_03276_));
 sky130_fd_sc_hd__buf_1 _22872_ (.A(\pcpi_mul.rs2[28] ),
    .X(_19319_));
 sky130_fd_sc_hd__buf_1 _22873_ (.A(_19319_),
    .X(_19320_));
 sky130_fd_sc_hd__buf_1 _22874_ (.A(_19320_),
    .X(_19321_));
 sky130_fd_sc_hd__mux2_2 _22875_ (.A0(pcpi_rs2[28]),
    .A1(_19321_),
    .S(_18172_),
    .X(_03275_));
 sky130_fd_sc_hd__buf_1 _22876_ (.A(\pcpi_mul.rs2[27] ),
    .X(_19322_));
 sky130_fd_sc_hd__buf_1 _22877_ (.A(_19322_),
    .X(_19323_));
 sky130_fd_sc_hd__buf_1 _22878_ (.A(_19323_),
    .X(_19324_));
 sky130_fd_sc_hd__buf_1 _22879_ (.A(_19324_),
    .X(_19325_));
 sky130_fd_sc_hd__buf_1 _22880_ (.A(_18171_),
    .X(_19326_));
 sky130_fd_sc_hd__mux2_2 _22881_ (.A0(_19135_),
    .A1(_19325_),
    .S(_19326_),
    .X(_03274_));
 sky130_fd_sc_hd__buf_1 _22882_ (.A(\pcpi_mul.rs2[26] ),
    .X(_19327_));
 sky130_fd_sc_hd__buf_1 _22883_ (.A(_19327_),
    .X(_19328_));
 sky130_fd_sc_hd__buf_1 _22884_ (.A(_19328_),
    .X(_19329_));
 sky130_fd_sc_hd__mux2_2 _22885_ (.A0(pcpi_rs2[26]),
    .A1(_19329_),
    .S(_19326_),
    .X(_03273_));
 sky130_fd_sc_hd__buf_1 _22886_ (.A(\pcpi_mul.rs2[25] ),
    .X(_19330_));
 sky130_fd_sc_hd__buf_1 _22887_ (.A(_19330_),
    .X(_19331_));
 sky130_fd_sc_hd__buf_1 _22888_ (.A(_19331_),
    .X(_19332_));
 sky130_fd_sc_hd__mux2_2 _22889_ (.A0(_19137_),
    .A1(_19332_),
    .S(_19326_),
    .X(_03272_));
 sky130_fd_sc_hd__buf_1 _22890_ (.A(\pcpi_mul.rs2[24] ),
    .X(_19333_));
 sky130_fd_sc_hd__buf_1 _22891_ (.A(_19333_),
    .X(_19334_));
 sky130_fd_sc_hd__buf_1 _22892_ (.A(_19334_),
    .X(_19335_));
 sky130_fd_sc_hd__mux2_2 _22893_ (.A0(pcpi_rs2[24]),
    .A1(_19335_),
    .S(_19326_),
    .X(_03271_));
 sky130_fd_sc_hd__buf_1 _22894_ (.A(\pcpi_mul.rs2[23] ),
    .X(_19336_));
 sky130_fd_sc_hd__buf_1 _22895_ (.A(_19336_),
    .X(_19337_));
 sky130_fd_sc_hd__buf_1 _22896_ (.A(_19337_),
    .X(_19338_));
 sky130_fd_sc_hd__mux2_2 _22897_ (.A0(_19138_),
    .A1(_19338_),
    .S(_19326_),
    .X(_03270_));
 sky130_fd_sc_hd__buf_2 _22898_ (.A(\pcpi_mul.rs2[22] ),
    .X(_19339_));
 sky130_fd_sc_hd__buf_1 _22899_ (.A(_19339_),
    .X(_19340_));
 sky130_fd_sc_hd__buf_1 _22900_ (.A(_19340_),
    .X(_19341_));
 sky130_fd_sc_hd__mux2_2 _22901_ (.A0(pcpi_rs2[22]),
    .A1(_19341_),
    .S(_19326_),
    .X(_03269_));
 sky130_fd_sc_hd__buf_1 _22902_ (.A(\pcpi_mul.rs2[21] ),
    .X(_19342_));
 sky130_fd_sc_hd__buf_1 _22903_ (.A(_19342_),
    .X(_19343_));
 sky130_fd_sc_hd__buf_1 _22904_ (.A(_19343_),
    .X(_19344_));
 sky130_fd_sc_hd__buf_1 _22905_ (.A(_18171_),
    .X(_19345_));
 sky130_fd_sc_hd__mux2_2 _22906_ (.A0(_19139_),
    .A1(_19344_),
    .S(_19345_),
    .X(_03268_));
 sky130_fd_sc_hd__buf_1 _22907_ (.A(\pcpi_mul.rs2[20] ),
    .X(_19346_));
 sky130_fd_sc_hd__buf_1 _22908_ (.A(_19346_),
    .X(_19347_));
 sky130_fd_sc_hd__buf_1 _22909_ (.A(_19347_),
    .X(_19348_));
 sky130_fd_sc_hd__mux2_2 _22910_ (.A0(pcpi_rs2[20]),
    .A1(_19348_),
    .S(_19345_),
    .X(_03267_));
 sky130_fd_sc_hd__buf_1 _22911_ (.A(\pcpi_mul.rs2[19] ),
    .X(_19349_));
 sky130_fd_sc_hd__buf_1 _22912_ (.A(_19349_),
    .X(_19350_));
 sky130_fd_sc_hd__buf_1 _22913_ (.A(_19350_),
    .X(_19351_));
 sky130_fd_sc_hd__mux2_2 _22914_ (.A0(pcpi_rs2[19]),
    .A1(_19351_),
    .S(_19345_),
    .X(_03266_));
 sky130_fd_sc_hd__buf_1 _22915_ (.A(\pcpi_mul.rs2[18] ),
    .X(_19352_));
 sky130_fd_sc_hd__buf_1 _22916_ (.A(_19352_),
    .X(_19353_));
 sky130_fd_sc_hd__mux2_2 _22917_ (.A0(_19141_),
    .A1(_19353_),
    .S(_19345_),
    .X(_03265_));
 sky130_fd_sc_hd__buf_1 _22918_ (.A(\pcpi_mul.rs2[17] ),
    .X(_19354_));
 sky130_fd_sc_hd__buf_1 _22919_ (.A(_19354_),
    .X(_19355_));
 sky130_fd_sc_hd__mux2_2 _22920_ (.A0(pcpi_rs2[17]),
    .A1(_19355_),
    .S(_19345_),
    .X(_03264_));
 sky130_fd_sc_hd__buf_1 _22921_ (.A(\pcpi_mul.rs2[16] ),
    .X(_19356_));
 sky130_fd_sc_hd__buf_1 _22922_ (.A(_19356_),
    .X(_19357_));
 sky130_fd_sc_hd__buf_1 _22923_ (.A(_19357_),
    .X(_19358_));
 sky130_fd_sc_hd__mux2_2 _22924_ (.A0(pcpi_rs2[16]),
    .A1(_19358_),
    .S(_19345_),
    .X(_03263_));
 sky130_fd_sc_hd__buf_1 _22925_ (.A(\pcpi_mul.rs2[15] ),
    .X(_19359_));
 sky130_fd_sc_hd__buf_1 _22926_ (.A(_19359_),
    .X(_19360_));
 sky130_fd_sc_hd__buf_1 _22927_ (.A(_18171_),
    .X(_19361_));
 sky130_fd_sc_hd__mux2_2 _22928_ (.A0(_19142_),
    .A1(_19360_),
    .S(_19361_),
    .X(_03262_));
 sky130_fd_sc_hd__buf_1 _22929_ (.A(\pcpi_mul.rs2[14] ),
    .X(_19362_));
 sky130_fd_sc_hd__buf_1 _22930_ (.A(_19362_),
    .X(_19363_));
 sky130_fd_sc_hd__buf_1 _22931_ (.A(_19363_),
    .X(_19364_));
 sky130_fd_sc_hd__mux2_2 _22932_ (.A0(_19143_),
    .A1(_19364_),
    .S(_19361_),
    .X(_03261_));
 sky130_fd_sc_hd__buf_1 _22933_ (.A(\pcpi_mul.rs2[13] ),
    .X(_19365_));
 sky130_fd_sc_hd__buf_1 _22934_ (.A(_19365_),
    .X(_19366_));
 sky130_fd_sc_hd__mux2_2 _22935_ (.A0(_19145_),
    .A1(_19366_),
    .S(_19361_),
    .X(_03260_));
 sky130_fd_sc_hd__buf_1 _22936_ (.A(\pcpi_mul.rs2[12] ),
    .X(_19367_));
 sky130_fd_sc_hd__buf_1 _22937_ (.A(_19367_),
    .X(_19368_));
 sky130_fd_sc_hd__buf_1 _22938_ (.A(_19368_),
    .X(_19369_));
 sky130_fd_sc_hd__mux2_2 _22939_ (.A0(pcpi_rs2[12]),
    .A1(_19369_),
    .S(_19361_),
    .X(_03259_));
 sky130_fd_sc_hd__buf_1 _22940_ (.A(\pcpi_mul.rs2[11] ),
    .X(_19370_));
 sky130_fd_sc_hd__buf_1 _22941_ (.A(_19370_),
    .X(_19371_));
 sky130_fd_sc_hd__mux2_2 _22942_ (.A0(_19146_),
    .A1(_19371_),
    .S(_19361_),
    .X(_03258_));
 sky130_fd_sc_hd__buf_1 _22943_ (.A(\pcpi_mul.rs2[10] ),
    .X(_19372_));
 sky130_fd_sc_hd__buf_1 _22944_ (.A(_19372_),
    .X(_19373_));
 sky130_fd_sc_hd__buf_1 _22945_ (.A(_19373_),
    .X(_19374_));
 sky130_fd_sc_hd__mux2_2 _22946_ (.A0(pcpi_rs2[10]),
    .A1(_19374_),
    .S(_19361_),
    .X(_03257_));
 sky130_fd_sc_hd__buf_1 _22947_ (.A(\pcpi_mul.rs2[9] ),
    .X(_19375_));
 sky130_fd_sc_hd__buf_1 _22948_ (.A(_19375_),
    .X(_19376_));
 sky130_fd_sc_hd__buf_1 _22949_ (.A(_19376_),
    .X(_19377_));
 sky130_fd_sc_hd__buf_1 _22950_ (.A(_18171_),
    .X(_19378_));
 sky130_fd_sc_hd__mux2_2 _22951_ (.A0(_19147_),
    .A1(_19377_),
    .S(_19378_),
    .X(_03256_));
 sky130_fd_sc_hd__buf_1 _22952_ (.A(\pcpi_mul.rs2[8] ),
    .X(_19379_));
 sky130_fd_sc_hd__buf_1 _22953_ (.A(_19379_),
    .X(_19380_));
 sky130_fd_sc_hd__buf_1 _22954_ (.A(_19380_),
    .X(_19381_));
 sky130_fd_sc_hd__mux2_2 _22955_ (.A0(pcpi_rs2[8]),
    .A1(_19381_),
    .S(_19378_),
    .X(_03255_));
 sky130_fd_sc_hd__buf_2 _22956_ (.A(\pcpi_mul.rs2[7] ),
    .X(_19382_));
 sky130_fd_sc_hd__buf_1 _22957_ (.A(_19382_),
    .X(_19383_));
 sky130_fd_sc_hd__buf_1 _22958_ (.A(_19383_),
    .X(_19384_));
 sky130_fd_sc_hd__mux2_2 _22959_ (.A0(_19149_),
    .A1(_19384_),
    .S(_19378_),
    .X(_03254_));
 sky130_fd_sc_hd__buf_1 _22960_ (.A(\pcpi_mul.rs2[6] ),
    .X(_19385_));
 sky130_fd_sc_hd__buf_1 _22961_ (.A(_19385_),
    .X(_19386_));
 sky130_fd_sc_hd__mux2_2 _22962_ (.A0(_19150_),
    .A1(_19386_),
    .S(_19378_),
    .X(_03253_));
 sky130_fd_sc_hd__buf_1 _22963_ (.A(\pcpi_mul.rs2[5] ),
    .X(_19387_));
 sky130_fd_sc_hd__buf_1 _22964_ (.A(_19387_),
    .X(_19388_));
 sky130_fd_sc_hd__buf_1 _22965_ (.A(_19388_),
    .X(_19389_));
 sky130_fd_sc_hd__mux2_2 _22966_ (.A0(_19151_),
    .A1(_19389_),
    .S(_19378_),
    .X(_03252_));
 sky130_fd_sc_hd__buf_1 _22967_ (.A(\pcpi_mul.rs2[4] ),
    .X(_19390_));
 sky130_fd_sc_hd__buf_1 _22968_ (.A(_19390_),
    .X(_19391_));
 sky130_fd_sc_hd__buf_1 _22969_ (.A(_19391_),
    .X(_19392_));
 sky130_fd_sc_hd__mux2_2 _22970_ (.A0(_19152_),
    .A1(_19392_),
    .S(_19378_),
    .X(_03251_));
 sky130_fd_sc_hd__buf_1 _22971_ (.A(\pcpi_mul.rs2[3] ),
    .X(_19393_));
 sky130_fd_sc_hd__buf_1 _22972_ (.A(_19393_),
    .X(_19394_));
 sky130_fd_sc_hd__buf_1 _22973_ (.A(_19394_),
    .X(_19395_));
 sky130_fd_sc_hd__buf_1 _22974_ (.A(_18174_),
    .X(_19396_));
 sky130_fd_sc_hd__mux2_2 _22975_ (.A0(_19153_),
    .A1(_19395_),
    .S(_19396_),
    .X(_03250_));
 sky130_fd_sc_hd__buf_1 _22976_ (.A(\pcpi_mul.rs2[2] ),
    .X(_19397_));
 sky130_fd_sc_hd__buf_1 _22977_ (.A(_19397_),
    .X(_19398_));
 sky130_fd_sc_hd__buf_1 _22978_ (.A(_19398_),
    .X(_19399_));
 sky130_fd_sc_hd__mux2_2 _22979_ (.A0(_19154_),
    .A1(_19399_),
    .S(_19396_),
    .X(_03249_));
 sky130_fd_sc_hd__buf_1 _22980_ (.A(\pcpi_mul.rs2[1] ),
    .X(_19400_));
 sky130_fd_sc_hd__buf_1 _22981_ (.A(_19400_),
    .X(_19401_));
 sky130_fd_sc_hd__buf_1 _22982_ (.A(_19401_),
    .X(_19402_));
 sky130_fd_sc_hd__mux2_2 _22983_ (.A0(_19155_),
    .A1(_19402_),
    .S(_19396_),
    .X(_03248_));
 sky130_fd_sc_hd__buf_1 _22984_ (.A(\pcpi_mul.rs2[0] ),
    .X(_19403_));
 sky130_fd_sc_hd__buf_1 _22985_ (.A(_19403_),
    .X(_19404_));
 sky130_fd_sc_hd__mux2_2 _22986_ (.A0(_19156_),
    .A1(_19404_),
    .S(_19396_),
    .X(_03247_));
 sky130_fd_sc_hd__mux2_2 _22987_ (.A0(mem_wstrb[3]),
    .A1(_02541_),
    .S(_18053_),
    .X(_03246_));
 sky130_fd_sc_hd__mux2_2 _22988_ (.A0(mem_wstrb[2]),
    .A1(_02540_),
    .S(_18053_),
    .X(_03245_));
 sky130_fd_sc_hd__mux2_2 _22989_ (.A0(mem_wstrb[1]),
    .A1(_02539_),
    .S(_18052_),
    .X(_03244_));
 sky130_fd_sc_hd__mux2_2 _22990_ (.A0(mem_wstrb[0]),
    .A1(_02538_),
    .S(_18052_),
    .X(_03243_));
 sky130_fd_sc_hd__and4_2 _22991_ (.A(_18060_),
    .B(_18064_),
    .C(_18063_),
    .D(_18062_),
    .X(_19405_));
 sky130_fd_sc_hd__buf_1 _22992_ (.A(_18343_),
    .X(_19406_));
 sky130_fd_sc_hd__a32o_2 _22993_ (.A1(_19405_),
    .A2(_00329_),
    .A3(_00328_),
    .B1(is_alu_reg_reg),
    .B2(_19406_),
    .X(_03242_));
 sky130_fd_sc_hd__inv_2 _22994_ (.A(_00329_),
    .Y(_19407_));
 sky130_fd_sc_hd__a32o_2 _22995_ (.A1(_19405_),
    .A2(_19407_),
    .A3(_00328_),
    .B1(is_alu_reg_imm),
    .B2(_19406_),
    .X(_03241_));
 sky130_fd_sc_hd__and2_2 _22996_ (.A(_19121_),
    .B(_19191_),
    .X(_19408_));
 sky130_fd_sc_hd__buf_1 _22997_ (.A(_19408_),
    .X(_19409_));
 sky130_fd_sc_hd__buf_1 _22998_ (.A(_19409_),
    .X(_19410_));
 sky130_fd_sc_hd__mux2_2 _22999_ (.A0(\cpuregs[13][31] ),
    .A1(\cpuregs_wrdata[31] ),
    .S(_19410_),
    .X(_03240_));
 sky130_fd_sc_hd__mux2_2 _23000_ (.A0(\cpuregs[13][30] ),
    .A1(\cpuregs_wrdata[30] ),
    .S(_19410_),
    .X(_03239_));
 sky130_fd_sc_hd__mux2_2 _23001_ (.A0(\cpuregs[13][29] ),
    .A1(\cpuregs_wrdata[29] ),
    .S(_19410_),
    .X(_03238_));
 sky130_fd_sc_hd__mux2_2 _23002_ (.A0(\cpuregs[13][28] ),
    .A1(\cpuregs_wrdata[28] ),
    .S(_19410_),
    .X(_03237_));
 sky130_fd_sc_hd__mux2_2 _23003_ (.A0(\cpuregs[13][27] ),
    .A1(\cpuregs_wrdata[27] ),
    .S(_19410_),
    .X(_03236_));
 sky130_fd_sc_hd__mux2_2 _23004_ (.A0(\cpuregs[13][26] ),
    .A1(\cpuregs_wrdata[26] ),
    .S(_19410_),
    .X(_03235_));
 sky130_fd_sc_hd__buf_1 _23005_ (.A(_19409_),
    .X(_19411_));
 sky130_fd_sc_hd__mux2_2 _23006_ (.A0(\cpuregs[13][25] ),
    .A1(\cpuregs_wrdata[25] ),
    .S(_19411_),
    .X(_03234_));
 sky130_fd_sc_hd__mux2_2 _23007_ (.A0(\cpuregs[13][24] ),
    .A1(\cpuregs_wrdata[24] ),
    .S(_19411_),
    .X(_03233_));
 sky130_fd_sc_hd__mux2_2 _23008_ (.A0(\cpuregs[13][23] ),
    .A1(\cpuregs_wrdata[23] ),
    .S(_19411_),
    .X(_03232_));
 sky130_fd_sc_hd__mux2_2 _23009_ (.A0(\cpuregs[13][22] ),
    .A1(\cpuregs_wrdata[22] ),
    .S(_19411_),
    .X(_03231_));
 sky130_fd_sc_hd__mux2_2 _23010_ (.A0(\cpuregs[13][21] ),
    .A1(\cpuregs_wrdata[21] ),
    .S(_19411_),
    .X(_03230_));
 sky130_fd_sc_hd__mux2_2 _23011_ (.A0(\cpuregs[13][20] ),
    .A1(\cpuregs_wrdata[20] ),
    .S(_19411_),
    .X(_03229_));
 sky130_fd_sc_hd__buf_1 _23012_ (.A(_19409_),
    .X(_19412_));
 sky130_fd_sc_hd__mux2_2 _23013_ (.A0(\cpuregs[13][19] ),
    .A1(\cpuregs_wrdata[19] ),
    .S(_19412_),
    .X(_03228_));
 sky130_fd_sc_hd__mux2_2 _23014_ (.A0(\cpuregs[13][18] ),
    .A1(\cpuregs_wrdata[18] ),
    .S(_19412_),
    .X(_03227_));
 sky130_fd_sc_hd__mux2_2 _23015_ (.A0(\cpuregs[13][17] ),
    .A1(\cpuregs_wrdata[17] ),
    .S(_19412_),
    .X(_03226_));
 sky130_fd_sc_hd__mux2_2 _23016_ (.A0(\cpuregs[13][16] ),
    .A1(\cpuregs_wrdata[16] ),
    .S(_19412_),
    .X(_03225_));
 sky130_fd_sc_hd__mux2_2 _23017_ (.A0(\cpuregs[13][15] ),
    .A1(\cpuregs_wrdata[15] ),
    .S(_19412_),
    .X(_03224_));
 sky130_fd_sc_hd__mux2_2 _23018_ (.A0(\cpuregs[13][14] ),
    .A1(\cpuregs_wrdata[14] ),
    .S(_19412_),
    .X(_03223_));
 sky130_fd_sc_hd__buf_1 _23019_ (.A(_19409_),
    .X(_19413_));
 sky130_fd_sc_hd__mux2_2 _23020_ (.A0(\cpuregs[13][13] ),
    .A1(\cpuregs_wrdata[13] ),
    .S(_19413_),
    .X(_03222_));
 sky130_fd_sc_hd__mux2_2 _23021_ (.A0(\cpuregs[13][12] ),
    .A1(\cpuregs_wrdata[12] ),
    .S(_19413_),
    .X(_03221_));
 sky130_fd_sc_hd__mux2_2 _23022_ (.A0(\cpuregs[13][11] ),
    .A1(\cpuregs_wrdata[11] ),
    .S(_19413_),
    .X(_03220_));
 sky130_fd_sc_hd__mux2_2 _23023_ (.A0(\cpuregs[13][10] ),
    .A1(\cpuregs_wrdata[10] ),
    .S(_19413_),
    .X(_03219_));
 sky130_fd_sc_hd__mux2_2 _23024_ (.A0(\cpuregs[13][9] ),
    .A1(\cpuregs_wrdata[9] ),
    .S(_19413_),
    .X(_03218_));
 sky130_fd_sc_hd__mux2_2 _23025_ (.A0(\cpuregs[13][8] ),
    .A1(\cpuregs_wrdata[8] ),
    .S(_19413_),
    .X(_03217_));
 sky130_fd_sc_hd__buf_1 _23026_ (.A(_19408_),
    .X(_19414_));
 sky130_fd_sc_hd__mux2_2 _23027_ (.A0(\cpuregs[13][7] ),
    .A1(\cpuregs_wrdata[7] ),
    .S(_19414_),
    .X(_03216_));
 sky130_fd_sc_hd__mux2_2 _23028_ (.A0(\cpuregs[13][6] ),
    .A1(\cpuregs_wrdata[6] ),
    .S(_19414_),
    .X(_03215_));
 sky130_fd_sc_hd__mux2_2 _23029_ (.A0(\cpuregs[13][5] ),
    .A1(\cpuregs_wrdata[5] ),
    .S(_19414_),
    .X(_03214_));
 sky130_fd_sc_hd__mux2_2 _23030_ (.A0(\cpuregs[13][4] ),
    .A1(\cpuregs_wrdata[4] ),
    .S(_19414_),
    .X(_03213_));
 sky130_fd_sc_hd__mux2_2 _23031_ (.A0(\cpuregs[13][3] ),
    .A1(\cpuregs_wrdata[3] ),
    .S(_19414_),
    .X(_03212_));
 sky130_fd_sc_hd__mux2_2 _23032_ (.A0(\cpuregs[13][2] ),
    .A1(\cpuregs_wrdata[2] ),
    .S(_19414_),
    .X(_03211_));
 sky130_fd_sc_hd__mux2_2 _23033_ (.A0(\cpuregs[13][1] ),
    .A1(\cpuregs_wrdata[1] ),
    .S(_19409_),
    .X(_03210_));
 sky130_fd_sc_hd__mux2_2 _23034_ (.A0(\cpuregs[13][0] ),
    .A1(\cpuregs_wrdata[0] ),
    .S(_19409_),
    .X(_03209_));
 sky130_fd_sc_hd__buf_1 _23035_ (.A(is_sb_sh_sw),
    .X(_19415_));
 sky130_fd_sc_hd__a32o_2 _23036_ (.A1(_19405_),
    .A2(_00329_),
    .A3(_18341_),
    .B1(_19415_),
    .B2(_19406_),
    .X(_03208_));
 sky130_fd_sc_hd__nor2_2 _23037_ (.A(instr_jalr),
    .B(_18877_),
    .Y(_19416_));
 sky130_fd_sc_hd__inv_2 _23038_ (.A(is_alu_reg_imm),
    .Y(_19417_));
 sky130_fd_sc_hd__a31o_2 _23039_ (.A1(_18399_),
    .A2(_18402_),
    .A3(_00335_),
    .B1(_19417_),
    .X(_19418_));
 sky130_fd_sc_hd__buf_1 _23040_ (.A(_18353_),
    .X(_19419_));
 sky130_fd_sc_hd__o2bb2a_2 _23041_ (.A1_N(_19416_),
    .A2_N(_19418_),
    .B1(is_jalr_addi_slti_sltiu_xori_ori_andi),
    .B2(_19419_),
    .X(_03207_));
 sky130_fd_sc_hd__o2111a_2 _23042_ (.A1(_18364_),
    .A2(_18379_),
    .B1(_18363_),
    .C1(_18365_),
    .D1(_18362_),
    .X(_19420_));
 sky130_fd_sc_hd__nor2_2 _23043_ (.A(\mem_rdata_q[13] ),
    .B(_18415_),
    .Y(_19421_));
 sky130_fd_sc_hd__buf_1 _23044_ (.A(is_slli_srli_srai),
    .X(_19422_));
 sky130_fd_sc_hd__buf_1 _23045_ (.A(_18392_),
    .X(_19423_));
 sky130_fd_sc_hd__a32o_2 _23046_ (.A1(_19420_),
    .A2(_18398_),
    .A3(_19421_),
    .B1(_19422_),
    .B2(_19423_),
    .X(_03206_));
 sky130_fd_sc_hd__a22o_2 _23047_ (.A1(is_lb_lh_lw_lbu_lhu),
    .A2(_18343_),
    .B1(_19405_),
    .B2(_18066_),
    .X(_03205_));
 sky130_fd_sc_hd__buf_1 _23048_ (.A(\decoded_imm_uj[20] ),
    .X(_19424_));
 sky130_fd_sc_hd__buf_1 _23049_ (.A(_19424_),
    .X(_19425_));
 sky130_fd_sc_hd__buf_1 _23050_ (.A(_19425_),
    .X(_19426_));
 sky130_fd_sc_hd__mux2_2 _23051_ (.A0(_19426_),
    .A1(\mem_rdata_latched[31] ),
    .S(_18077_),
    .X(_03204_));
 sky130_fd_sc_hd__mux2_2 _23052_ (.A0(\decoded_imm_uj[19] ),
    .A1(\mem_rdata_latched[19] ),
    .S(_18077_),
    .X(_03203_));
 sky130_fd_sc_hd__inv_2 _23053_ (.A(\decoded_imm_uj[18] ),
    .Y(_19427_));
 sky130_fd_sc_hd__o21ai_2 _23054_ (.A1(_19427_),
    .A2(_20587_),
    .B1(_18345_),
    .Y(_03202_));
 sky130_fd_sc_hd__inv_2 _23055_ (.A(\decoded_imm_uj[17] ),
    .Y(_19428_));
 sky130_fd_sc_hd__o21ai_2 _23056_ (.A1(_19428_),
    .A2(_20587_),
    .B1(_18346_),
    .Y(_03201_));
 sky130_fd_sc_hd__inv_2 _23057_ (.A(\decoded_imm_uj[16] ),
    .Y(_19429_));
 sky130_fd_sc_hd__o21ai_2 _23058_ (.A1(_19429_),
    .A2(_20587_),
    .B1(_18347_),
    .Y(_03200_));
 sky130_fd_sc_hd__inv_2 _23059_ (.A(\decoded_imm_uj[15] ),
    .Y(_19430_));
 sky130_fd_sc_hd__o21ai_2 _23060_ (.A1(_19430_),
    .A2(_20587_),
    .B1(_18348_),
    .Y(_03199_));
 sky130_fd_sc_hd__buf_1 _23061_ (.A(_18060_),
    .X(_19431_));
 sky130_fd_sc_hd__mux2_2 _23062_ (.A0(\decoded_imm_uj[14] ),
    .A1(\mem_rdata_latched[14] ),
    .S(_19431_),
    .X(_03198_));
 sky130_fd_sc_hd__mux2_2 _23063_ (.A0(\decoded_imm_uj[13] ),
    .A1(\mem_rdata_latched[13] ),
    .S(_19431_),
    .X(_03197_));
 sky130_fd_sc_hd__mux2_2 _23064_ (.A0(\decoded_imm_uj[12] ),
    .A1(\mem_rdata_latched[12] ),
    .S(_19431_),
    .X(_03196_));
 sky130_fd_sc_hd__mux2_2 _23065_ (.A0(\decoded_imm_uj[11] ),
    .A1(\mem_rdata_latched[20] ),
    .S(_19431_),
    .X(_03195_));
 sky130_fd_sc_hd__mux2_2 _23066_ (.A0(\decoded_imm_uj[10] ),
    .A1(\mem_rdata_latched[30] ),
    .S(_19431_),
    .X(_03194_));
 sky130_fd_sc_hd__mux2_2 _23067_ (.A0(\decoded_imm_uj[9] ),
    .A1(\mem_rdata_latched[29] ),
    .S(_19431_),
    .X(_03193_));
 sky130_fd_sc_hd__buf_1 _23068_ (.A(_18060_),
    .X(_19432_));
 sky130_fd_sc_hd__mux2_2 _23069_ (.A0(\decoded_imm_uj[8] ),
    .A1(\mem_rdata_latched[28] ),
    .S(_19432_),
    .X(_03192_));
 sky130_fd_sc_hd__nor2_2 _23070_ (.A(_18068_),
    .B(_18343_),
    .Y(_19433_));
 sky130_fd_sc_hd__a21o_2 _23071_ (.A1(\decoded_imm_uj[7] ),
    .A2(_00337_),
    .B1(_19433_),
    .X(_03191_));
 sky130_fd_sc_hd__mux2_2 _23072_ (.A0(\decoded_imm_uj[6] ),
    .A1(\mem_rdata_latched[26] ),
    .S(_19432_),
    .X(_03190_));
 sky130_fd_sc_hd__mux2_2 _23073_ (.A0(\decoded_imm_uj[5] ),
    .A1(\mem_rdata_latched[25] ),
    .S(_19432_),
    .X(_03189_));
 sky130_fd_sc_hd__mux2_2 _23074_ (.A0(\decoded_imm_uj[4] ),
    .A1(\mem_rdata_latched[24] ),
    .S(_19432_),
    .X(_03188_));
 sky130_fd_sc_hd__mux2_2 _23075_ (.A0(\decoded_imm_uj[3] ),
    .A1(\mem_rdata_latched[23] ),
    .S(_19432_),
    .X(_03187_));
 sky130_fd_sc_hd__mux2_2 _23076_ (.A0(\decoded_imm_uj[2] ),
    .A1(\mem_rdata_latched[22] ),
    .S(_19432_),
    .X(_03186_));
 sky130_fd_sc_hd__buf_1 _23077_ (.A(_18060_),
    .X(_19434_));
 sky130_fd_sc_hd__mux2_2 _23078_ (.A0(\decoded_imm_uj[1] ),
    .A1(\mem_rdata_latched[21] ),
    .S(_19434_),
    .X(_03185_));
 sky130_fd_sc_hd__or3_2 _23079_ (.A(is_alu_reg_imm),
    .B(is_lb_lh_lw_lbu_lhu),
    .C(instr_jalr),
    .X(_19435_));
 sky130_fd_sc_hd__buf_1 _23080_ (.A(_19435_),
    .X(_19436_));
 sky130_fd_sc_hd__a22o_2 _23081_ (.A1(_19415_),
    .A2(\mem_rdata_q[7] ),
    .B1(_19436_),
    .B2(\mem_rdata_q[20] ),
    .X(_19437_));
 sky130_fd_sc_hd__mux2_2 _23082_ (.A0(_19437_),
    .A1(\decoded_imm[0] ),
    .S(_18386_),
    .X(_03184_));
 sky130_fd_sc_hd__mux2_2 _23083_ (.A0(\decoded_rd[4] ),
    .A1(\mem_rdata_latched[11] ),
    .S(_19434_),
    .X(_03183_));
 sky130_fd_sc_hd__mux2_2 _23084_ (.A0(\decoded_rd[3] ),
    .A1(\mem_rdata_latched[10] ),
    .S(_19434_),
    .X(_03182_));
 sky130_fd_sc_hd__mux2_2 _23085_ (.A0(\decoded_rd[2] ),
    .A1(\mem_rdata_latched[9] ),
    .S(_19434_),
    .X(_03181_));
 sky130_fd_sc_hd__mux2_2 _23086_ (.A0(\decoded_rd[1] ),
    .A1(\mem_rdata_latched[8] ),
    .S(_19434_),
    .X(_03180_));
 sky130_fd_sc_hd__mux2_2 _23087_ (.A0(\decoded_rd[0] ),
    .A1(\mem_rdata_latched[7] ),
    .S(_19434_),
    .X(_03179_));
 sky130_fd_sc_hd__buf_1 _23088_ (.A(instr_timer),
    .X(_19438_));
 sky130_fd_sc_hd__buf_1 _23089_ (.A(_19438_),
    .X(_19439_));
 sky130_fd_sc_hd__buf_1 _23090_ (.A(_18385_),
    .X(_19440_));
 sky130_fd_sc_hd__inv_2 _23091_ (.A(\mem_rdata_q[3] ),
    .Y(_19441_));
 sky130_fd_sc_hd__or4_2 _23092_ (.A(\mem_rdata_q[6] ),
    .B(\mem_rdata_q[5] ),
    .C(\mem_rdata_q[4] ),
    .D(_19441_),
    .X(_19442_));
 sky130_fd_sc_hd__inv_2 _23093_ (.A(\mem_rdata_q[2] ),
    .Y(_19443_));
 sky130_fd_sc_hd__and4b_2 _23094_ (.A_N(_19442_),
    .B(_19443_),
    .C(\mem_rdata_q[1] ),
    .D(\mem_rdata_q[0] ),
    .X(_19444_));
 sky130_fd_sc_hd__buf_1 _23095_ (.A(\mem_rdata_q[25] ),
    .X(_19445_));
 sky130_fd_sc_hd__and3_2 _23096_ (.A(_18366_),
    .B(_19445_),
    .C(_18359_),
    .X(_19446_));
 sky130_fd_sc_hd__buf_1 _23097_ (.A(_18352_),
    .X(_19447_));
 sky130_fd_sc_hd__and3_2 _23098_ (.A(_19446_),
    .B(\mem_rdata_q[27] ),
    .C(_19447_),
    .X(_19448_));
 sky130_fd_sc_hd__a22o_2 _23099_ (.A1(_19439_),
    .A2(_19440_),
    .B1(_19444_),
    .B2(_19448_),
    .X(_03178_));
 sky130_fd_sc_hd__a32o_2 _23100_ (.A1(_19433_),
    .A2(_18067_),
    .A3(_18075_),
    .B1(instr_waitirq),
    .B2(_19406_),
    .X(_03177_));
 sky130_fd_sc_hd__buf_1 _23101_ (.A(decoder_trigger),
    .X(_19449_));
 sky130_fd_sc_hd__and3_2 _23102_ (.A(_18360_),
    .B(_18375_),
    .C(_19449_),
    .X(_19450_));
 sky130_fd_sc_hd__inv_2 _23103_ (.A(\mem_rdata_q[28] ),
    .Y(_19451_));
 sky130_fd_sc_hd__buf_1 _23104_ (.A(\mem_rdata_q[26] ),
    .X(_19452_));
 sky130_fd_sc_hd__and4_2 _23105_ (.A(_18366_),
    .B(_19451_),
    .C(_19452_),
    .D(_19445_),
    .X(_19453_));
 sky130_fd_sc_hd__buf_1 _23106_ (.A(_18198_),
    .X(_19454_));
 sky130_fd_sc_hd__a32o_2 _23107_ (.A1(_19444_),
    .A2(_19450_),
    .A3(_19453_),
    .B1(_19454_),
    .B2(_19423_),
    .X(_03176_));
 sky130_fd_sc_hd__o21ai_2 _23108_ (.A1(_18033_),
    .A2(_18061_),
    .B1(_18074_),
    .Y(_03175_));
 sky130_fd_sc_hd__a32o_2 _23109_ (.A1(_19444_),
    .A2(_19446_),
    .A3(_19450_),
    .B1(instr_setq),
    .B2(_19423_),
    .X(_03174_));
 sky130_fd_sc_hd__a22o_2 _23110_ (.A1(instr_getq),
    .A2(_19440_),
    .B1(_19444_),
    .B2(_18388_),
    .X(_03173_));
 sky130_fd_sc_hd__buf_1 _23111_ (.A(\mem_rdata_q[24] ),
    .X(_19455_));
 sky130_fd_sc_hd__or4_2 _23112_ (.A(_19455_),
    .B(\mem_rdata_q[21] ),
    .C(\mem_rdata_q[11] ),
    .D(\mem_rdata_q[10] ),
    .X(_19456_));
 sky130_fd_sc_hd__or3_2 _23113_ (.A(\mem_rdata_q[17] ),
    .B(\mem_rdata_q[16] ),
    .C(\mem_rdata_q[15] ),
    .X(_19457_));
 sky130_fd_sc_hd__or4_2 _23114_ (.A(\mem_rdata_q[9] ),
    .B(\mem_rdata_q[8] ),
    .C(\mem_rdata_q[7] ),
    .D(_18409_),
    .X(_19458_));
 sky130_fd_sc_hd__nor2_2 _23115_ (.A(_19457_),
    .B(_19458_),
    .Y(_19459_));
 sky130_fd_sc_hd__nor2_2 _23116_ (.A(\mem_rdata_q[19] ),
    .B(\mem_rdata_q[18] ),
    .Y(_19460_));
 sky130_fd_sc_hd__and3b_2 _23117_ (.A_N(_19456_),
    .B(_19459_),
    .C(_19460_),
    .X(_19461_));
 sky130_fd_sc_hd__and3_2 _23118_ (.A(_19441_),
    .B(_19443_),
    .C(\mem_rdata_q[4] ),
    .X(_19462_));
 sky130_fd_sc_hd__nor2_2 _23119_ (.A(\mem_rdata_q[23] ),
    .B(\mem_rdata_q[22] ),
    .Y(_19463_));
 sky130_fd_sc_hd__and4_2 _23120_ (.A(\mem_rdata_q[6] ),
    .B(\mem_rdata_q[5] ),
    .C(\mem_rdata_q[1] ),
    .D(\mem_rdata_q[0] ),
    .X(_19464_));
 sky130_fd_sc_hd__and3_2 _23121_ (.A(_19462_),
    .B(_19463_),
    .C(_19464_),
    .X(_19465_));
 sky130_fd_sc_hd__a32o_2 _23122_ (.A1(_19461_),
    .A2(_18388_),
    .A3(_19465_),
    .B1(instr_ecall_ebreak),
    .B2(_19440_),
    .X(_03172_));
 sky130_fd_sc_hd__inv_2 _23123_ (.A(\mem_rdata_q[20] ),
    .Y(_19466_));
 sky130_fd_sc_hd__and3_2 _23124_ (.A(_19466_),
    .B(_18375_),
    .C(_19449_),
    .X(_19467_));
 sky130_fd_sc_hd__nand3_2 _23125_ (.A(_19465_),
    .B(\mem_rdata_q[21] ),
    .C(_19467_),
    .Y(_19468_));
 sky130_fd_sc_hd__nand2_2 _23126_ (.A(_18365_),
    .B(_19451_),
    .Y(_19469_));
 sky130_fd_sc_hd__nand2_2 _23127_ (.A(\mem_rdata_q[31] ),
    .B(\mem_rdata_q[30] ),
    .Y(_19470_));
 sky130_fd_sc_hd__or4_2 _23128_ (.A(\mem_rdata_q[26] ),
    .B(_19445_),
    .C(\mem_rdata_q[24] ),
    .D(_18360_),
    .X(_19471_));
 sky130_fd_sc_hd__or3b_2 _23129_ (.A(_18402_),
    .B(_19457_),
    .C_N(_19460_),
    .X(_19472_));
 sky130_fd_sc_hd__or4_2 _23130_ (.A(_19469_),
    .B(_19470_),
    .C(_19471_),
    .D(_19472_),
    .X(_19473_));
 sky130_fd_sc_hd__buf_1 _23131_ (.A(instr_rdinstrh),
    .X(_19474_));
 sky130_fd_sc_hd__buf_1 _23132_ (.A(_18427_),
    .X(_19475_));
 sky130_fd_sc_hd__a2bb2o_2 _23133_ (.A1_N(_19468_),
    .A2_N(_19473_),
    .B1(_19474_),
    .B2(_19475_),
    .X(_03171_));
 sky130_fd_sc_hd__or4_2 _23134_ (.A(\mem_rdata_q[27] ),
    .B(\mem_rdata_q[25] ),
    .C(_19470_),
    .D(_19469_),
    .X(_19476_));
 sky130_fd_sc_hd__or4_2 _23135_ (.A(_19452_),
    .B(_19455_),
    .C(_19476_),
    .D(_19472_),
    .X(_19477_));
 sky130_fd_sc_hd__buf_1 _23136_ (.A(instr_rdinstr),
    .X(_19478_));
 sky130_fd_sc_hd__a2bb2o_2 _23137_ (.A1_N(_19468_),
    .A2_N(_19477_),
    .B1(_19478_),
    .B2(_19475_),
    .X(_03170_));
 sky130_fd_sc_hd__inv_2 _23138_ (.A(\mem_rdata_q[21] ),
    .Y(_19479_));
 sky130_fd_sc_hd__and3_2 _23139_ (.A(_19479_),
    .B(_18375_),
    .C(_19449_),
    .X(_19480_));
 sky130_fd_sc_hd__nand2_2 _23140_ (.A(_19465_),
    .B(_19480_),
    .Y(_19481_));
 sky130_fd_sc_hd__buf_1 _23141_ (.A(instr_rdcycleh),
    .X(_19482_));
 sky130_fd_sc_hd__a2bb2o_2 _23142_ (.A1_N(_19481_),
    .A2_N(_19473_),
    .B1(_19482_),
    .B2(_19475_),
    .X(_03169_));
 sky130_fd_sc_hd__a2bb2o_2 _23143_ (.A1_N(_19481_),
    .A2_N(_19477_),
    .B1(instr_rdcycle),
    .B2(_19475_),
    .X(_03168_));
 sky130_fd_sc_hd__nor2_2 _23144_ (.A(_19417_),
    .B(_18381_),
    .Y(_19483_));
 sky130_fd_sc_hd__a22o_2 _23145_ (.A1(instr_srai),
    .A2(_18877_),
    .B1(_18378_),
    .B2(_19483_),
    .X(_03167_));
 sky130_fd_sc_hd__a22o_2 _23146_ (.A1(instr_srli),
    .A2(_18877_),
    .B1(_18388_),
    .B2(_19483_),
    .X(_03166_));
 sky130_fd_sc_hd__a32o_2 _23147_ (.A1(_18388_),
    .A2(is_alu_reg_imm),
    .A3(_18405_),
    .B1(instr_slli),
    .B2(_19440_),
    .X(_03165_));
 sky130_fd_sc_hd__and3_2 _23148_ (.A(_18375_),
    .B(_19415_),
    .C(_19449_),
    .X(_19484_));
 sky130_fd_sc_hd__a22o_2 _23149_ (.A1(instr_sw),
    .A2(_18877_),
    .B1(_18403_),
    .B2(_19484_),
    .X(_03164_));
 sky130_fd_sc_hd__a22o_2 _23150_ (.A1(_18405_),
    .A2(_19484_),
    .B1(_19475_),
    .B2(instr_sh),
    .X(_03163_));
 sky130_fd_sc_hd__a22o_2 _23151_ (.A1(_18408_),
    .A2(_19484_),
    .B1(instr_sb),
    .B2(_19440_),
    .X(_03162_));
 sky130_fd_sc_hd__and3_2 _23152_ (.A(_18375_),
    .B(is_lb_lh_lw_lbu_lhu),
    .C(_19449_),
    .X(_19485_));
 sky130_fd_sc_hd__a22o_2 _23153_ (.A1(_18380_),
    .A2(_19485_),
    .B1(_19423_),
    .B2(instr_lhu),
    .X(_03161_));
 sky130_fd_sc_hd__a22o_2 _23154_ (.A1(_18393_),
    .A2(_19485_),
    .B1(_19423_),
    .B2(instr_lbu),
    .X(_03160_));
 sky130_fd_sc_hd__a22o_2 _23155_ (.A1(instr_lw),
    .A2(_18877_),
    .B1(_18403_),
    .B2(_19485_),
    .X(_03159_));
 sky130_fd_sc_hd__a22o_2 _23156_ (.A1(_18405_),
    .A2(_19485_),
    .B1(_19423_),
    .B2(instr_lh),
    .X(_03158_));
 sky130_fd_sc_hd__a22o_2 _23157_ (.A1(_18408_),
    .A2(_19485_),
    .B1(instr_lb),
    .B2(_19440_),
    .X(_03157_));
 sky130_fd_sc_hd__nor3_2 _23158_ (.A(\mem_rdata_latched[14] ),
    .B(\mem_rdata_latched[13] ),
    .C(\mem_rdata_latched[12] ),
    .Y(_19486_));
 sky130_fd_sc_hd__and3_2 _23159_ (.A(_00325_),
    .B(_00324_),
    .C(_00326_),
    .X(_19487_));
 sky130_fd_sc_hd__and2_2 _23160_ (.A(_19487_),
    .B(_18064_),
    .X(_19488_));
 sky130_fd_sc_hd__nor2_2 _23161_ (.A(_02063_),
    .B(_18059_),
    .Y(_19489_));
 sky130_fd_sc_hd__a41o_2 _23162_ (.A1(_18061_),
    .A2(_18342_),
    .A3(_19486_),
    .A4(_19488_),
    .B1(_19489_),
    .X(_03156_));
 sky130_fd_sc_hd__nor2_2 _23163_ (.A(_00323_),
    .B(_18059_),
    .Y(_19490_));
 sky130_fd_sc_hd__a41o_2 _23164_ (.A1(_00327_),
    .A2(_18061_),
    .A3(_18342_),
    .A4(_19487_),
    .B1(_19490_),
    .X(_03155_));
 sky130_fd_sc_hd__and3_2 _23165_ (.A(_18059_),
    .B(_18063_),
    .C(_19488_),
    .X(_19491_));
 sky130_fd_sc_hd__a32o_2 _23166_ (.A1(_19491_),
    .A2(_19407_),
    .A3(_00328_),
    .B1(instr_auipc),
    .B2(_19406_),
    .X(_03154_));
 sky130_fd_sc_hd__buf_1 _23167_ (.A(instr_lui),
    .X(_19492_));
 sky130_fd_sc_hd__a32o_2 _23168_ (.A1(_19491_),
    .A2(_00329_),
    .A3(_00328_),
    .B1(_19492_),
    .B2(_19406_),
    .X(_03153_));
 sky130_fd_sc_hd__buf_1 _23169_ (.A(\mem_rdata_q[31] ),
    .X(_19493_));
 sky130_fd_sc_hd__buf_1 _23170_ (.A(_19447_),
    .X(_19494_));
 sky130_fd_sc_hd__mux2_2 _23171_ (.A0(pcpi_insn[31]),
    .A1(_19493_),
    .S(_19494_),
    .X(_03152_));
 sky130_fd_sc_hd__mux2_2 _23172_ (.A0(pcpi_insn[30]),
    .A1(\mem_rdata_q[30] ),
    .S(_19494_),
    .X(_03151_));
 sky130_fd_sc_hd__buf_1 _23173_ (.A(_19447_),
    .X(_19495_));
 sky130_fd_sc_hd__o21ba_2 _23174_ (.A1(pcpi_insn[29]),
    .A2(_19495_),
    .B1_N(_18376_),
    .X(_03150_));
 sky130_fd_sc_hd__mux2_2 _23175_ (.A0(pcpi_insn[28]),
    .A1(\mem_rdata_q[28] ),
    .S(_19494_),
    .X(_03149_));
 sky130_fd_sc_hd__o21ba_2 _23176_ (.A1(pcpi_insn[27]),
    .A2(_19495_),
    .B1_N(_19450_),
    .X(_03148_));
 sky130_fd_sc_hd__mux2_2 _23177_ (.A0(pcpi_insn[26]),
    .A1(_19452_),
    .S(_19494_),
    .X(_03147_));
 sky130_fd_sc_hd__mux2_2 _23178_ (.A0(pcpi_insn[25]),
    .A1(_19445_),
    .S(_19494_),
    .X(_03146_));
 sky130_fd_sc_hd__buf_1 _23179_ (.A(_19447_),
    .X(_19496_));
 sky130_fd_sc_hd__mux2_2 _23180_ (.A0(pcpi_insn[24]),
    .A1(_19455_),
    .S(_19496_),
    .X(_03145_));
 sky130_fd_sc_hd__mux2_2 _23181_ (.A0(pcpi_insn[23]),
    .A1(\mem_rdata_q[23] ),
    .S(_19496_),
    .X(_03144_));
 sky130_fd_sc_hd__mux2_2 _23182_ (.A0(pcpi_insn[22]),
    .A1(\mem_rdata_q[22] ),
    .S(_19496_),
    .X(_03143_));
 sky130_fd_sc_hd__o21ba_2 _23183_ (.A1(pcpi_insn[21]),
    .A2(_19495_),
    .B1_N(_19480_),
    .X(_03142_));
 sky130_fd_sc_hd__o21ba_2 _23184_ (.A1(pcpi_insn[20]),
    .A2(_19494_),
    .B1_N(_19467_),
    .X(_03141_));
 sky130_fd_sc_hd__mux2_2 _23185_ (.A0(pcpi_insn[19]),
    .A1(\mem_rdata_q[19] ),
    .S(_19496_),
    .X(_03140_));
 sky130_fd_sc_hd__mux2_2 _23186_ (.A0(pcpi_insn[18]),
    .A1(\mem_rdata_q[18] ),
    .S(_19496_),
    .X(_03139_));
 sky130_fd_sc_hd__mux2_2 _23187_ (.A0(pcpi_insn[17]),
    .A1(\mem_rdata_q[17] ),
    .S(_19496_),
    .X(_03138_));
 sky130_fd_sc_hd__buf_1 _23188_ (.A(_19447_),
    .X(_19497_));
 sky130_fd_sc_hd__mux2_2 _23189_ (.A0(pcpi_insn[16]),
    .A1(\mem_rdata_q[16] ),
    .S(_19497_),
    .X(_03137_));
 sky130_fd_sc_hd__mux2_2 _23190_ (.A0(pcpi_insn[15]),
    .A1(\mem_rdata_q[15] ),
    .S(_19497_),
    .X(_03136_));
 sky130_fd_sc_hd__mux2_2 _23191_ (.A0(pcpi_insn[14]),
    .A1(_18379_),
    .S(_19497_),
    .X(_03135_));
 sky130_fd_sc_hd__mux2_2 _23192_ (.A0(pcpi_insn[13]),
    .A1(\mem_rdata_q[13] ),
    .S(_19497_),
    .X(_03134_));
 sky130_fd_sc_hd__mux2_2 _23193_ (.A0(pcpi_insn[12]),
    .A1(_18398_),
    .S(_19497_),
    .X(_03133_));
 sky130_fd_sc_hd__mux2_2 _23194_ (.A0(pcpi_insn[11]),
    .A1(\mem_rdata_q[11] ),
    .S(_19497_),
    .X(_03132_));
 sky130_fd_sc_hd__buf_1 _23195_ (.A(_18352_),
    .X(_19498_));
 sky130_fd_sc_hd__mux2_2 _23196_ (.A0(pcpi_insn[10]),
    .A1(\mem_rdata_q[10] ),
    .S(_19498_),
    .X(_03131_));
 sky130_fd_sc_hd__mux2_2 _23197_ (.A0(pcpi_insn[9]),
    .A1(\mem_rdata_q[9] ),
    .S(_19498_),
    .X(_03130_));
 sky130_fd_sc_hd__mux2_2 _23198_ (.A0(pcpi_insn[8]),
    .A1(\mem_rdata_q[8] ),
    .S(_19498_),
    .X(_03129_));
 sky130_fd_sc_hd__mux2_2 _23199_ (.A0(pcpi_insn[7]),
    .A1(\mem_rdata_q[7] ),
    .S(_19498_),
    .X(_03128_));
 sky130_fd_sc_hd__mux2_2 _23200_ (.A0(pcpi_insn[6]),
    .A1(\mem_rdata_q[6] ),
    .S(_19498_),
    .X(_03127_));
 sky130_fd_sc_hd__mux2_2 _23201_ (.A0(pcpi_insn[5]),
    .A1(\mem_rdata_q[5] ),
    .S(_19498_),
    .X(_03126_));
 sky130_fd_sc_hd__buf_1 _23202_ (.A(_18352_),
    .X(_19499_));
 sky130_fd_sc_hd__mux2_2 _23203_ (.A0(pcpi_insn[4]),
    .A1(\mem_rdata_q[4] ),
    .S(_19499_),
    .X(_03125_));
 sky130_fd_sc_hd__mux2_2 _23204_ (.A0(pcpi_insn[3]),
    .A1(\mem_rdata_q[3] ),
    .S(_19499_),
    .X(_03124_));
 sky130_fd_sc_hd__mux2_2 _23205_ (.A0(pcpi_insn[2]),
    .A1(\mem_rdata_q[2] ),
    .S(_19499_),
    .X(_03123_));
 sky130_fd_sc_hd__mux2_2 _23206_ (.A0(pcpi_insn[1]),
    .A1(\mem_rdata_q[1] ),
    .S(_19499_),
    .X(_03122_));
 sky130_fd_sc_hd__mux2_2 _23207_ (.A0(pcpi_insn[0]),
    .A1(\mem_rdata_q[0] ),
    .S(_19499_),
    .X(_03121_));
 sky130_fd_sc_hd__inv_2 _23208_ (.A(\cpu_state[5] ),
    .Y(_19500_));
 sky130_fd_sc_hd__or3_2 _23209_ (.A(_00318_),
    .B(_00320_),
    .C(_18016_),
    .X(_19501_));
 sky130_fd_sc_hd__a31o_2 _23210_ (.A1(_18193_),
    .A2(_18205_),
    .A3(_19500_),
    .B1(_19501_),
    .X(_19502_));
 sky130_fd_sc_hd__buf_1 _23211_ (.A(_19502_),
    .X(_19503_));
 sky130_fd_sc_hd__buf_1 _23212_ (.A(_19503_),
    .X(_19504_));
 sky130_fd_sc_hd__mux2_2 _23213_ (.A0(_02499_),
    .A1(pcpi_rs1[31]),
    .S(_19504_),
    .X(_03120_));
 sky130_fd_sc_hd__buf_1 _23214_ (.A(pcpi_rs1[30]),
    .X(_19505_));
 sky130_fd_sc_hd__mux2_2 _23215_ (.A0(_02498_),
    .A1(_19505_),
    .S(_19504_),
    .X(_03119_));
 sky130_fd_sc_hd__buf_1 _23216_ (.A(pcpi_rs1[29]),
    .X(_19506_));
 sky130_fd_sc_hd__mux2_2 _23217_ (.A0(_02496_),
    .A1(_19506_),
    .S(_19504_),
    .X(_03118_));
 sky130_fd_sc_hd__buf_1 _23218_ (.A(pcpi_rs1[28]),
    .X(_19507_));
 sky130_fd_sc_hd__mux2_2 _23219_ (.A0(_02495_),
    .A1(_19507_),
    .S(_19504_),
    .X(_03117_));
 sky130_fd_sc_hd__mux2_2 _23220_ (.A0(_02494_),
    .A1(pcpi_rs1[27]),
    .S(_19504_),
    .X(_03116_));
 sky130_fd_sc_hd__buf_1 _23221_ (.A(pcpi_rs1[26]),
    .X(_19508_));
 sky130_fd_sc_hd__mux2_2 _23222_ (.A0(_02493_),
    .A1(_19508_),
    .S(_19504_),
    .X(_03115_));
 sky130_fd_sc_hd__buf_1 _23223_ (.A(pcpi_rs1[25]),
    .X(_19509_));
 sky130_fd_sc_hd__buf_1 _23224_ (.A(_19503_),
    .X(_19510_));
 sky130_fd_sc_hd__mux2_2 _23225_ (.A0(_02492_),
    .A1(_19509_),
    .S(_19510_),
    .X(_03114_));
 sky130_fd_sc_hd__buf_1 _23226_ (.A(pcpi_rs1[24]),
    .X(_19511_));
 sky130_fd_sc_hd__mux2_2 _23227_ (.A0(_02491_),
    .A1(_19511_),
    .S(_19510_),
    .X(_03113_));
 sky130_fd_sc_hd__buf_1 _23228_ (.A(pcpi_rs1[23]),
    .X(_19512_));
 sky130_fd_sc_hd__mux2_2 _23229_ (.A0(_02490_),
    .A1(_19512_),
    .S(_19510_),
    .X(_03112_));
 sky130_fd_sc_hd__buf_1 _23230_ (.A(pcpi_rs1[22]),
    .X(_19513_));
 sky130_fd_sc_hd__mux2_2 _23231_ (.A0(_02489_),
    .A1(_19513_),
    .S(_19510_),
    .X(_03111_));
 sky130_fd_sc_hd__buf_1 _23232_ (.A(pcpi_rs1[21]),
    .X(_19514_));
 sky130_fd_sc_hd__mux2_2 _23233_ (.A0(_02488_),
    .A1(_19514_),
    .S(_19510_),
    .X(_03110_));
 sky130_fd_sc_hd__mux2_2 _23234_ (.A0(_02487_),
    .A1(pcpi_rs1[20]),
    .S(_19510_),
    .X(_03109_));
 sky130_fd_sc_hd__buf_1 _23235_ (.A(pcpi_rs1[19]),
    .X(_19515_));
 sky130_fd_sc_hd__buf_1 _23236_ (.A(_19503_),
    .X(_19516_));
 sky130_fd_sc_hd__mux2_2 _23237_ (.A0(_02485_),
    .A1(_19515_),
    .S(_19516_),
    .X(_03108_));
 sky130_fd_sc_hd__buf_1 _23238_ (.A(pcpi_rs1[18]),
    .X(_19517_));
 sky130_fd_sc_hd__mux2_2 _23239_ (.A0(_02484_),
    .A1(_19517_),
    .S(_19516_),
    .X(_03107_));
 sky130_fd_sc_hd__buf_1 _23240_ (.A(pcpi_rs1[17]),
    .X(_19518_));
 sky130_fd_sc_hd__mux2_2 _23241_ (.A0(_02483_),
    .A1(_19518_),
    .S(_19516_),
    .X(_03106_));
 sky130_fd_sc_hd__buf_1 _23242_ (.A(pcpi_rs1[16]),
    .X(_19519_));
 sky130_fd_sc_hd__mux2_2 _23243_ (.A0(_02482_),
    .A1(_19519_),
    .S(_19516_),
    .X(_03105_));
 sky130_fd_sc_hd__buf_1 _23244_ (.A(pcpi_rs1[15]),
    .X(_19520_));
 sky130_fd_sc_hd__mux2_2 _23245_ (.A0(_02481_),
    .A1(_19520_),
    .S(_19516_),
    .X(_03104_));
 sky130_fd_sc_hd__mux2_2 _23246_ (.A0(_02480_),
    .A1(pcpi_rs1[14]),
    .S(_19516_),
    .X(_03103_));
 sky130_fd_sc_hd__buf_1 _23247_ (.A(pcpi_rs1[13]),
    .X(_19521_));
 sky130_fd_sc_hd__buf_1 _23248_ (.A(_19503_),
    .X(_19522_));
 sky130_fd_sc_hd__mux2_2 _23249_ (.A0(_02479_),
    .A1(_19521_),
    .S(_19522_),
    .X(_03102_));
 sky130_fd_sc_hd__buf_1 _23250_ (.A(pcpi_rs1[12]),
    .X(_19523_));
 sky130_fd_sc_hd__mux2_2 _23251_ (.A0(_02478_),
    .A1(_19523_),
    .S(_19522_),
    .X(_03101_));
 sky130_fd_sc_hd__buf_1 _23252_ (.A(pcpi_rs1[11]),
    .X(_19524_));
 sky130_fd_sc_hd__mux2_2 _23253_ (.A0(_02477_),
    .A1(_19524_),
    .S(_19522_),
    .X(_03100_));
 sky130_fd_sc_hd__mux2_2 _23254_ (.A0(_02476_),
    .A1(pcpi_rs1[10]),
    .S(_19522_),
    .X(_03099_));
 sky130_fd_sc_hd__buf_1 _23255_ (.A(pcpi_rs1[9]),
    .X(_19525_));
 sky130_fd_sc_hd__mux2_2 _23256_ (.A0(_02506_),
    .A1(_19525_),
    .S(_19522_),
    .X(_03098_));
 sky130_fd_sc_hd__buf_1 _23257_ (.A(pcpi_rs1[8]),
    .X(_19526_));
 sky130_fd_sc_hd__mux2_2 _23258_ (.A0(_02505_),
    .A1(_19526_),
    .S(_19522_),
    .X(_03097_));
 sky130_fd_sc_hd__buf_1 _23259_ (.A(_19502_),
    .X(_19527_));
 sky130_fd_sc_hd__mux2_2 _23260_ (.A0(_02504_),
    .A1(pcpi_rs1[7]),
    .S(_19527_),
    .X(_03096_));
 sky130_fd_sc_hd__buf_1 _23261_ (.A(pcpi_rs1[6]),
    .X(_19528_));
 sky130_fd_sc_hd__mux2_2 _23262_ (.A0(_02503_),
    .A1(_19528_),
    .S(_19527_),
    .X(_03095_));
 sky130_fd_sc_hd__buf_1 _23263_ (.A(pcpi_rs1[5]),
    .X(_19529_));
 sky130_fd_sc_hd__mux2_2 _23264_ (.A0(_02502_),
    .A1(_19529_),
    .S(_19527_),
    .X(_03094_));
 sky130_fd_sc_hd__buf_1 _23265_ (.A(pcpi_rs1[4]),
    .X(_19530_));
 sky130_fd_sc_hd__mux2_2 _23266_ (.A0(_02501_),
    .A1(_19530_),
    .S(_19527_),
    .X(_03093_));
 sky130_fd_sc_hd__buf_1 _23267_ (.A(pcpi_rs1[3]),
    .X(_19531_));
 sky130_fd_sc_hd__mux2_2 _23268_ (.A0(_02500_),
    .A1(_19531_),
    .S(_19527_),
    .X(_03092_));
 sky130_fd_sc_hd__buf_1 _23269_ (.A(pcpi_rs1[2]),
    .X(_19532_));
 sky130_fd_sc_hd__mux2_2 _23270_ (.A0(_02497_),
    .A1(_19532_),
    .S(_19527_),
    .X(_03091_));
 sky130_fd_sc_hd__buf_1 _23271_ (.A(pcpi_rs1[1]),
    .X(_19533_));
 sky130_fd_sc_hd__buf_1 _23272_ (.A(_19533_),
    .X(_19534_));
 sky130_fd_sc_hd__mux2_2 _23273_ (.A0(_02486_),
    .A1(_19534_),
    .S(_19503_),
    .X(_03090_));
 sky130_fd_sc_hd__buf_1 _23274_ (.A(pcpi_rs1[0]),
    .X(_19535_));
 sky130_fd_sc_hd__mux2_2 _23275_ (.A0(_02475_),
    .A1(_19535_),
    .S(_19503_),
    .X(_03089_));
 sky130_fd_sc_hd__mux2_2 _23276_ (.A0(mem_addr[31]),
    .A1(mem_la_addr[31]),
    .S(_18337_),
    .X(_03088_));
 sky130_fd_sc_hd__mux2_2 _23277_ (.A0(mem_addr[30]),
    .A1(mem_la_addr[30]),
    .S(_18337_),
    .X(_03087_));
 sky130_fd_sc_hd__mux2_2 _23278_ (.A0(mem_addr[29]),
    .A1(mem_la_addr[29]),
    .S(_18337_),
    .X(_03086_));
 sky130_fd_sc_hd__mux2_2 _23279_ (.A0(mem_addr[28]),
    .A1(mem_la_addr[28]),
    .S(_18337_),
    .X(_03085_));
 sky130_fd_sc_hd__mux2_2 _23280_ (.A0(mem_addr[27]),
    .A1(mem_la_addr[27]),
    .S(_18337_),
    .X(_03084_));
 sky130_fd_sc_hd__buf_1 _23281_ (.A(_18336_),
    .X(_19536_));
 sky130_fd_sc_hd__mux2_2 _23282_ (.A0(mem_addr[26]),
    .A1(mem_la_addr[26]),
    .S(_19536_),
    .X(_03083_));
 sky130_fd_sc_hd__mux2_2 _23283_ (.A0(mem_addr[25]),
    .A1(mem_la_addr[25]),
    .S(_19536_),
    .X(_03082_));
 sky130_fd_sc_hd__mux2_2 _23284_ (.A0(mem_addr[24]),
    .A1(mem_la_addr[24]),
    .S(_19536_),
    .X(_03081_));
 sky130_fd_sc_hd__mux2_2 _23285_ (.A0(mem_addr[23]),
    .A1(mem_la_addr[23]),
    .S(_19536_),
    .X(_03080_));
 sky130_fd_sc_hd__mux2_2 _23286_ (.A0(mem_addr[22]),
    .A1(mem_la_addr[22]),
    .S(_19536_),
    .X(_03079_));
 sky130_fd_sc_hd__mux2_2 _23287_ (.A0(mem_addr[21]),
    .A1(mem_la_addr[21]),
    .S(_19536_),
    .X(_03078_));
 sky130_fd_sc_hd__buf_1 _23288_ (.A(_18336_),
    .X(_19537_));
 sky130_fd_sc_hd__mux2_2 _23289_ (.A0(mem_addr[20]),
    .A1(mem_la_addr[20]),
    .S(_19537_),
    .X(_03077_));
 sky130_fd_sc_hd__mux2_2 _23290_ (.A0(mem_addr[19]),
    .A1(mem_la_addr[19]),
    .S(_19537_),
    .X(_03076_));
 sky130_fd_sc_hd__mux2_2 _23291_ (.A0(mem_addr[18]),
    .A1(mem_la_addr[18]),
    .S(_19537_),
    .X(_03075_));
 sky130_fd_sc_hd__mux2_2 _23292_ (.A0(mem_addr[17]),
    .A1(mem_la_addr[17]),
    .S(_19537_),
    .X(_03074_));
 sky130_fd_sc_hd__mux2_2 _23293_ (.A0(mem_addr[16]),
    .A1(mem_la_addr[16]),
    .S(_19537_),
    .X(_03073_));
 sky130_fd_sc_hd__mux2_2 _23294_ (.A0(mem_addr[15]),
    .A1(mem_la_addr[15]),
    .S(_19537_),
    .X(_03072_));
 sky130_fd_sc_hd__buf_1 _23295_ (.A(_18336_),
    .X(_19538_));
 sky130_fd_sc_hd__mux2_2 _23296_ (.A0(mem_addr[14]),
    .A1(mem_la_addr[14]),
    .S(_19538_),
    .X(_03071_));
 sky130_fd_sc_hd__mux2_2 _23297_ (.A0(mem_addr[13]),
    .A1(mem_la_addr[13]),
    .S(_19538_),
    .X(_03070_));
 sky130_fd_sc_hd__mux2_2 _23298_ (.A0(mem_addr[12]),
    .A1(mem_la_addr[12]),
    .S(_19538_),
    .X(_03069_));
 sky130_fd_sc_hd__mux2_2 _23299_ (.A0(mem_addr[11]),
    .A1(mem_la_addr[11]),
    .S(_19538_),
    .X(_03068_));
 sky130_fd_sc_hd__mux2_2 _23300_ (.A0(mem_addr[10]),
    .A1(mem_la_addr[10]),
    .S(_19538_),
    .X(_03067_));
 sky130_fd_sc_hd__mux2_2 _23301_ (.A0(mem_addr[9]),
    .A1(mem_la_addr[9]),
    .S(_19538_),
    .X(_03066_));
 sky130_fd_sc_hd__buf_1 _23302_ (.A(_18336_),
    .X(_19539_));
 sky130_fd_sc_hd__mux2_2 _23303_ (.A0(mem_addr[8]),
    .A1(mem_la_addr[8]),
    .S(_19539_),
    .X(_03065_));
 sky130_fd_sc_hd__mux2_2 _23304_ (.A0(mem_addr[7]),
    .A1(mem_la_addr[7]),
    .S(_19539_),
    .X(_03064_));
 sky130_fd_sc_hd__mux2_2 _23305_ (.A0(mem_addr[6]),
    .A1(mem_la_addr[6]),
    .S(_19539_),
    .X(_03063_));
 sky130_fd_sc_hd__mux2_2 _23306_ (.A0(mem_addr[5]),
    .A1(mem_la_addr[5]),
    .S(_19539_),
    .X(_03062_));
 sky130_fd_sc_hd__mux2_2 _23307_ (.A0(mem_addr[4]),
    .A1(mem_la_addr[4]),
    .S(_19539_),
    .X(_03061_));
 sky130_fd_sc_hd__mux2_2 _23308_ (.A0(mem_addr[3]),
    .A1(mem_la_addr[3]),
    .S(_19539_),
    .X(_03060_));
 sky130_fd_sc_hd__mux2_2 _23309_ (.A0(mem_addr[2]),
    .A1(mem_la_addr[2]),
    .S(_18336_),
    .X(_03059_));
 sky130_fd_sc_hd__buf_1 _23310_ (.A(\pcpi_mul.rs1[31] ),
    .X(_19540_));
 sky130_fd_sc_hd__buf_1 _23311_ (.A(_19540_),
    .X(_19541_));
 sky130_fd_sc_hd__buf_1 _23312_ (.A(_19541_),
    .X(_19542_));
 sky130_fd_sc_hd__buf_1 _23313_ (.A(_19542_),
    .X(_19543_));
 sky130_fd_sc_hd__a21o_2 _23314_ (.A1(_19543_),
    .A2(_18172_),
    .B1(_18176_),
    .X(_03058_));
 sky130_fd_sc_hd__buf_1 _23315_ (.A(\pcpi_mul.rs1[30] ),
    .X(_19544_));
 sky130_fd_sc_hd__buf_1 _23316_ (.A(_19544_),
    .X(_19545_));
 sky130_fd_sc_hd__buf_1 _23317_ (.A(_19545_),
    .X(_19546_));
 sky130_fd_sc_hd__buf_1 _23318_ (.A(_19546_),
    .X(_19547_));
 sky130_fd_sc_hd__mux2_2 _23319_ (.A0(_19505_),
    .A1(_19547_),
    .S(_19396_),
    .X(_03057_));
 sky130_fd_sc_hd__buf_1 _23320_ (.A(\pcpi_mul.rs1[29] ),
    .X(_19548_));
 sky130_fd_sc_hd__buf_1 _23321_ (.A(_19548_),
    .X(_19549_));
 sky130_fd_sc_hd__buf_1 _23322_ (.A(_19549_),
    .X(_19550_));
 sky130_fd_sc_hd__buf_1 _23323_ (.A(_19550_),
    .X(_19551_));
 sky130_fd_sc_hd__mux2_2 _23324_ (.A0(_19506_),
    .A1(_19551_),
    .S(_19396_),
    .X(_03056_));
 sky130_fd_sc_hd__buf_1 _23325_ (.A(\pcpi_mul.rs1[28] ),
    .X(_19552_));
 sky130_fd_sc_hd__buf_1 _23326_ (.A(_19552_),
    .X(_19553_));
 sky130_fd_sc_hd__buf_1 _23327_ (.A(_19553_),
    .X(_19554_));
 sky130_fd_sc_hd__buf_1 _23328_ (.A(_19554_),
    .X(_19555_));
 sky130_fd_sc_hd__buf_1 _23329_ (.A(_18174_),
    .X(_19556_));
 sky130_fd_sc_hd__mux2_2 _23330_ (.A0(_19507_),
    .A1(_19555_),
    .S(_19556_),
    .X(_03055_));
 sky130_fd_sc_hd__buf_1 _23331_ (.A(\pcpi_mul.rs1[27] ),
    .X(_19557_));
 sky130_fd_sc_hd__buf_1 _23332_ (.A(_19557_),
    .X(_19558_));
 sky130_fd_sc_hd__buf_1 _23333_ (.A(_19558_),
    .X(_19559_));
 sky130_fd_sc_hd__buf_1 _23334_ (.A(_19559_),
    .X(_19560_));
 sky130_fd_sc_hd__mux2_2 _23335_ (.A0(pcpi_rs1[27]),
    .A1(_19560_),
    .S(_19556_),
    .X(_03054_));
 sky130_fd_sc_hd__buf_1 _23336_ (.A(\pcpi_mul.rs1[26] ),
    .X(_19561_));
 sky130_fd_sc_hd__buf_1 _23337_ (.A(_19561_),
    .X(_19562_));
 sky130_fd_sc_hd__buf_1 _23338_ (.A(_19562_),
    .X(_19563_));
 sky130_fd_sc_hd__mux2_2 _23339_ (.A0(_19508_),
    .A1(_19563_),
    .S(_19556_),
    .X(_03053_));
 sky130_fd_sc_hd__buf_1 _23340_ (.A(\pcpi_mul.rs1[25] ),
    .X(_19564_));
 sky130_fd_sc_hd__buf_1 _23341_ (.A(_19564_),
    .X(_19565_));
 sky130_fd_sc_hd__buf_1 _23342_ (.A(_19565_),
    .X(_19566_));
 sky130_fd_sc_hd__mux2_2 _23343_ (.A0(_19509_),
    .A1(_19566_),
    .S(_19556_),
    .X(_03052_));
 sky130_fd_sc_hd__buf_1 _23344_ (.A(\pcpi_mul.rs1[24] ),
    .X(_19567_));
 sky130_fd_sc_hd__buf_1 _23345_ (.A(_19567_),
    .X(_19568_));
 sky130_fd_sc_hd__buf_1 _23346_ (.A(_19568_),
    .X(_19569_));
 sky130_fd_sc_hd__mux2_2 _23347_ (.A0(_19511_),
    .A1(_19569_),
    .S(_19556_),
    .X(_03051_));
 sky130_fd_sc_hd__buf_1 _23348_ (.A(\pcpi_mul.rs1[23] ),
    .X(_19570_));
 sky130_fd_sc_hd__buf_1 _23349_ (.A(_19570_),
    .X(_19571_));
 sky130_fd_sc_hd__buf_1 _23350_ (.A(_19571_),
    .X(_19572_));
 sky130_fd_sc_hd__mux2_2 _23351_ (.A0(_19512_),
    .A1(_19572_),
    .S(_19556_),
    .X(_03050_));
 sky130_fd_sc_hd__buf_1 _23352_ (.A(\pcpi_mul.rs1[22] ),
    .X(_19573_));
 sky130_fd_sc_hd__buf_1 _23353_ (.A(_19573_),
    .X(_19574_));
 sky130_fd_sc_hd__buf_1 _23354_ (.A(_19574_),
    .X(_19575_));
 sky130_fd_sc_hd__buf_1 _23355_ (.A(_18174_),
    .X(_19576_));
 sky130_fd_sc_hd__mux2_2 _23356_ (.A0(_19513_),
    .A1(_19575_),
    .S(_19576_),
    .X(_03049_));
 sky130_fd_sc_hd__buf_1 _23357_ (.A(\pcpi_mul.rs1[21] ),
    .X(_19577_));
 sky130_fd_sc_hd__buf_1 _23358_ (.A(_19577_),
    .X(_19578_));
 sky130_fd_sc_hd__buf_1 _23359_ (.A(_19578_),
    .X(_19579_));
 sky130_fd_sc_hd__mux2_2 _23360_ (.A0(_19514_),
    .A1(_19579_),
    .S(_19576_),
    .X(_03048_));
 sky130_fd_sc_hd__buf_1 _23361_ (.A(\pcpi_mul.rs1[20] ),
    .X(_19580_));
 sky130_fd_sc_hd__buf_1 _23362_ (.A(_19580_),
    .X(_19581_));
 sky130_fd_sc_hd__mux2_2 _23363_ (.A0(pcpi_rs1[20]),
    .A1(_19581_),
    .S(_19576_),
    .X(_03047_));
 sky130_fd_sc_hd__buf_1 _23364_ (.A(\pcpi_mul.rs1[19] ),
    .X(_19582_));
 sky130_fd_sc_hd__buf_1 _23365_ (.A(_19582_),
    .X(_19583_));
 sky130_fd_sc_hd__mux2_2 _23366_ (.A0(_19515_),
    .A1(_19583_),
    .S(_19576_),
    .X(_03046_));
 sky130_fd_sc_hd__buf_2 _23367_ (.A(\pcpi_mul.rs1[18] ),
    .X(_19584_));
 sky130_fd_sc_hd__buf_2 _23368_ (.A(_19584_),
    .X(_19585_));
 sky130_fd_sc_hd__buf_1 _23369_ (.A(_19585_),
    .X(_19586_));
 sky130_fd_sc_hd__mux2_2 _23370_ (.A0(_19517_),
    .A1(_19586_),
    .S(_19576_),
    .X(_03045_));
 sky130_fd_sc_hd__buf_1 _23371_ (.A(\pcpi_mul.rs1[17] ),
    .X(_19587_));
 sky130_fd_sc_hd__buf_1 _23372_ (.A(_19587_),
    .X(_19588_));
 sky130_fd_sc_hd__buf_1 _23373_ (.A(_19588_),
    .X(_19589_));
 sky130_fd_sc_hd__mux2_2 _23374_ (.A0(_19518_),
    .A1(_19589_),
    .S(_19576_),
    .X(_03044_));
 sky130_fd_sc_hd__buf_1 _23375_ (.A(\pcpi_mul.rs1[16] ),
    .X(_19590_));
 sky130_fd_sc_hd__buf_1 _23376_ (.A(_19590_),
    .X(_19591_));
 sky130_fd_sc_hd__buf_1 _23377_ (.A(_18174_),
    .X(_19592_));
 sky130_fd_sc_hd__mux2_2 _23378_ (.A0(_19519_),
    .A1(_19591_),
    .S(_19592_),
    .X(_03043_));
 sky130_fd_sc_hd__buf_1 _23379_ (.A(\pcpi_mul.rs1[15] ),
    .X(_19593_));
 sky130_fd_sc_hd__buf_1 _23380_ (.A(_19593_),
    .X(_19594_));
 sky130_fd_sc_hd__buf_1 _23381_ (.A(_19594_),
    .X(_19595_));
 sky130_fd_sc_hd__mux2_2 _23382_ (.A0(_19520_),
    .A1(_19595_),
    .S(_19592_),
    .X(_03042_));
 sky130_fd_sc_hd__buf_1 _23383_ (.A(\pcpi_mul.rs1[14] ),
    .X(_19596_));
 sky130_fd_sc_hd__buf_1 _23384_ (.A(_19596_),
    .X(_19597_));
 sky130_fd_sc_hd__buf_1 _23385_ (.A(_19597_),
    .X(_19598_));
 sky130_fd_sc_hd__mux2_2 _23386_ (.A0(pcpi_rs1[14]),
    .A1(_19598_),
    .S(_19592_),
    .X(_03041_));
 sky130_fd_sc_hd__buf_1 _23387_ (.A(\pcpi_mul.rs1[13] ),
    .X(_19599_));
 sky130_fd_sc_hd__buf_1 _23388_ (.A(_19599_),
    .X(_19600_));
 sky130_fd_sc_hd__buf_1 _23389_ (.A(_19600_),
    .X(_19601_));
 sky130_fd_sc_hd__mux2_2 _23390_ (.A0(_19521_),
    .A1(_19601_),
    .S(_19592_),
    .X(_03040_));
 sky130_fd_sc_hd__buf_2 _23391_ (.A(\pcpi_mul.rs1[12] ),
    .X(_19602_));
 sky130_fd_sc_hd__buf_1 _23392_ (.A(_19602_),
    .X(_19603_));
 sky130_fd_sc_hd__buf_1 _23393_ (.A(_19603_),
    .X(_19604_));
 sky130_fd_sc_hd__mux2_2 _23394_ (.A0(_19523_),
    .A1(_19604_),
    .S(_19592_),
    .X(_03039_));
 sky130_fd_sc_hd__buf_1 _23395_ (.A(\pcpi_mul.rs1[11] ),
    .X(_19605_));
 sky130_fd_sc_hd__buf_1 _23396_ (.A(_19605_),
    .X(_19606_));
 sky130_fd_sc_hd__buf_1 _23397_ (.A(_19606_),
    .X(_19607_));
 sky130_fd_sc_hd__mux2_2 _23398_ (.A0(_19524_),
    .A1(_19607_),
    .S(_19592_),
    .X(_03038_));
 sky130_fd_sc_hd__buf_1 _23399_ (.A(\pcpi_mul.rs1[10] ),
    .X(_19608_));
 sky130_fd_sc_hd__buf_1 _23400_ (.A(_19608_),
    .X(_19609_));
 sky130_fd_sc_hd__buf_1 _23401_ (.A(_19609_),
    .X(_19610_));
 sky130_fd_sc_hd__buf_1 _23402_ (.A(_18174_),
    .X(_19611_));
 sky130_fd_sc_hd__mux2_2 _23403_ (.A0(pcpi_rs1[10]),
    .A1(_19610_),
    .S(_19611_),
    .X(_03037_));
 sky130_fd_sc_hd__buf_1 _23404_ (.A(\pcpi_mul.rs1[9] ),
    .X(_19612_));
 sky130_fd_sc_hd__buf_1 _23405_ (.A(_19612_),
    .X(_19613_));
 sky130_fd_sc_hd__buf_1 _23406_ (.A(_19613_),
    .X(_19614_));
 sky130_fd_sc_hd__mux2_2 _23407_ (.A0(_19525_),
    .A1(_19614_),
    .S(_19611_),
    .X(_03036_));
 sky130_fd_sc_hd__buf_1 _23408_ (.A(\pcpi_mul.rs1[8] ),
    .X(_19615_));
 sky130_fd_sc_hd__buf_1 _23409_ (.A(_19615_),
    .X(_19616_));
 sky130_fd_sc_hd__buf_1 _23410_ (.A(_19616_),
    .X(_19617_));
 sky130_fd_sc_hd__mux2_2 _23411_ (.A0(_19526_),
    .A1(_19617_),
    .S(_19611_),
    .X(_03035_));
 sky130_fd_sc_hd__buf_1 _23412_ (.A(\pcpi_mul.rs1[7] ),
    .X(_19618_));
 sky130_fd_sc_hd__buf_1 _23413_ (.A(_19618_),
    .X(_19619_));
 sky130_fd_sc_hd__buf_1 _23414_ (.A(_19619_),
    .X(_19620_));
 sky130_fd_sc_hd__mux2_2 _23415_ (.A0(pcpi_rs1[7]),
    .A1(_19620_),
    .S(_19611_),
    .X(_03034_));
 sky130_fd_sc_hd__buf_1 _23416_ (.A(\pcpi_mul.rs1[6] ),
    .X(_19621_));
 sky130_fd_sc_hd__buf_1 _23417_ (.A(_19621_),
    .X(_19622_));
 sky130_fd_sc_hd__buf_1 _23418_ (.A(_19622_),
    .X(_19623_));
 sky130_fd_sc_hd__mux2_2 _23419_ (.A0(_19528_),
    .A1(_19623_),
    .S(_19611_),
    .X(_03033_));
 sky130_fd_sc_hd__buf_1 _23420_ (.A(\pcpi_mul.rs1[5] ),
    .X(_19624_));
 sky130_fd_sc_hd__buf_1 _23421_ (.A(_19624_),
    .X(_19625_));
 sky130_fd_sc_hd__buf_1 _23422_ (.A(_19625_),
    .X(_19626_));
 sky130_fd_sc_hd__mux2_2 _23423_ (.A0(_19529_),
    .A1(_19626_),
    .S(_19611_),
    .X(_03032_));
 sky130_fd_sc_hd__buf_1 _23424_ (.A(\pcpi_mul.rs1[4] ),
    .X(_19627_));
 sky130_fd_sc_hd__buf_1 _23425_ (.A(_19627_),
    .X(_19628_));
 sky130_fd_sc_hd__mux2_2 _23426_ (.A0(_19530_),
    .A1(_19628_),
    .S(_18175_),
    .X(_03031_));
 sky130_fd_sc_hd__buf_1 _23427_ (.A(\pcpi_mul.rs1[3] ),
    .X(_19629_));
 sky130_fd_sc_hd__buf_1 _23428_ (.A(_19629_),
    .X(_19630_));
 sky130_fd_sc_hd__buf_1 _23429_ (.A(_19630_),
    .X(_19631_));
 sky130_fd_sc_hd__mux2_2 _23430_ (.A0(_19531_),
    .A1(_19631_),
    .S(_18175_),
    .X(_03030_));
 sky130_fd_sc_hd__buf_1 _23431_ (.A(\pcpi_mul.rs1[2] ),
    .X(_19632_));
 sky130_fd_sc_hd__buf_1 _23432_ (.A(_19632_),
    .X(_19633_));
 sky130_fd_sc_hd__buf_1 _23433_ (.A(_19633_),
    .X(_19634_));
 sky130_fd_sc_hd__mux2_2 _23434_ (.A0(_19532_),
    .A1(_19634_),
    .S(_18175_),
    .X(_03029_));
 sky130_fd_sc_hd__buf_1 _23435_ (.A(\pcpi_mul.rs1[1] ),
    .X(_19635_));
 sky130_fd_sc_hd__buf_1 _23436_ (.A(_19635_),
    .X(_19636_));
 sky130_fd_sc_hd__buf_1 _23437_ (.A(_19636_),
    .X(_19637_));
 sky130_fd_sc_hd__buf_1 _23438_ (.A(_19637_),
    .X(_19638_));
 sky130_fd_sc_hd__mux2_2 _23439_ (.A0(_19534_),
    .A1(_19638_),
    .S(_18175_),
    .X(_03028_));
 sky130_fd_sc_hd__buf_1 _23440_ (.A(\pcpi_mul.rs1[0] ),
    .X(_19639_));
 sky130_fd_sc_hd__buf_1 _23441_ (.A(_19639_),
    .X(_19640_));
 sky130_fd_sc_hd__buf_1 _23442_ (.A(_19640_),
    .X(_19641_));
 sky130_fd_sc_hd__buf_1 _23443_ (.A(_19641_),
    .X(_19642_));
 sky130_fd_sc_hd__mux2_2 _23444_ (.A0(_19535_),
    .A1(_19642_),
    .S(_18175_),
    .X(_03027_));
 sky130_fd_sc_hd__nand2_2 _23445_ (.A(_19121_),
    .B(_19082_),
    .Y(_19643_));
 sky130_fd_sc_hd__buf_1 _23446_ (.A(_19643_),
    .X(_19644_));
 sky130_fd_sc_hd__buf_1 _23447_ (.A(_19644_),
    .X(_19645_));
 sky130_fd_sc_hd__mux2_2 _23448_ (.A0(_19199_),
    .A1(\cpuregs[5][31] ),
    .S(_19645_),
    .X(_03026_));
 sky130_fd_sc_hd__mux2_2 _23449_ (.A0(_19203_),
    .A1(\cpuregs[5][30] ),
    .S(_19645_),
    .X(_03025_));
 sky130_fd_sc_hd__mux2_2 _23450_ (.A0(_19204_),
    .A1(\cpuregs[5][29] ),
    .S(_19645_),
    .X(_03024_));
 sky130_fd_sc_hd__mux2_2 _23451_ (.A0(_19205_),
    .A1(\cpuregs[5][28] ),
    .S(_19645_),
    .X(_03023_));
 sky130_fd_sc_hd__mux2_2 _23452_ (.A0(_19206_),
    .A1(\cpuregs[5][27] ),
    .S(_19645_),
    .X(_03022_));
 sky130_fd_sc_hd__mux2_2 _23453_ (.A0(_19207_),
    .A1(\cpuregs[5][26] ),
    .S(_19645_),
    .X(_03021_));
 sky130_fd_sc_hd__buf_1 _23454_ (.A(_19644_),
    .X(_19646_));
 sky130_fd_sc_hd__mux2_2 _23455_ (.A0(_19208_),
    .A1(\cpuregs[5][25] ),
    .S(_19646_),
    .X(_03020_));
 sky130_fd_sc_hd__mux2_2 _23456_ (.A0(_19210_),
    .A1(\cpuregs[5][24] ),
    .S(_19646_),
    .X(_03019_));
 sky130_fd_sc_hd__mux2_2 _23457_ (.A0(_19211_),
    .A1(\cpuregs[5][23] ),
    .S(_19646_),
    .X(_03018_));
 sky130_fd_sc_hd__mux2_2 _23458_ (.A0(_19212_),
    .A1(\cpuregs[5][22] ),
    .S(_19646_),
    .X(_03017_));
 sky130_fd_sc_hd__mux2_2 _23459_ (.A0(_19213_),
    .A1(\cpuregs[5][21] ),
    .S(_19646_),
    .X(_03016_));
 sky130_fd_sc_hd__mux2_2 _23460_ (.A0(_19214_),
    .A1(\cpuregs[5][20] ),
    .S(_19646_),
    .X(_03015_));
 sky130_fd_sc_hd__buf_1 _23461_ (.A(_19644_),
    .X(_19647_));
 sky130_fd_sc_hd__mux2_2 _23462_ (.A0(_19215_),
    .A1(\cpuregs[5][19] ),
    .S(_19647_),
    .X(_03014_));
 sky130_fd_sc_hd__mux2_2 _23463_ (.A0(_19217_),
    .A1(\cpuregs[5][18] ),
    .S(_19647_),
    .X(_03013_));
 sky130_fd_sc_hd__mux2_2 _23464_ (.A0(_19218_),
    .A1(\cpuregs[5][17] ),
    .S(_19647_),
    .X(_03012_));
 sky130_fd_sc_hd__mux2_2 _23465_ (.A0(_19219_),
    .A1(\cpuregs[5][16] ),
    .S(_19647_),
    .X(_03011_));
 sky130_fd_sc_hd__mux2_2 _23466_ (.A0(_19220_),
    .A1(\cpuregs[5][15] ),
    .S(_19647_),
    .X(_03010_));
 sky130_fd_sc_hd__mux2_2 _23467_ (.A0(_19221_),
    .A1(\cpuregs[5][14] ),
    .S(_19647_),
    .X(_03009_));
 sky130_fd_sc_hd__buf_1 _23468_ (.A(_19644_),
    .X(_19648_));
 sky130_fd_sc_hd__mux2_2 _23469_ (.A0(_19222_),
    .A1(\cpuregs[5][13] ),
    .S(_19648_),
    .X(_03008_));
 sky130_fd_sc_hd__mux2_2 _23470_ (.A0(_19224_),
    .A1(\cpuregs[5][12] ),
    .S(_19648_),
    .X(_03007_));
 sky130_fd_sc_hd__mux2_2 _23471_ (.A0(_19225_),
    .A1(\cpuregs[5][11] ),
    .S(_19648_),
    .X(_03006_));
 sky130_fd_sc_hd__mux2_2 _23472_ (.A0(_19226_),
    .A1(\cpuregs[5][10] ),
    .S(_19648_),
    .X(_03005_));
 sky130_fd_sc_hd__mux2_2 _23473_ (.A0(_19227_),
    .A1(\cpuregs[5][9] ),
    .S(_19648_),
    .X(_03004_));
 sky130_fd_sc_hd__mux2_2 _23474_ (.A0(_19228_),
    .A1(\cpuregs[5][8] ),
    .S(_19648_),
    .X(_03003_));
 sky130_fd_sc_hd__buf_1 _23475_ (.A(_19643_),
    .X(_19649_));
 sky130_fd_sc_hd__mux2_2 _23476_ (.A0(_19229_),
    .A1(\cpuregs[5][7] ),
    .S(_19649_),
    .X(_03002_));
 sky130_fd_sc_hd__mux2_2 _23477_ (.A0(_19231_),
    .A1(\cpuregs[5][6] ),
    .S(_19649_),
    .X(_03001_));
 sky130_fd_sc_hd__mux2_2 _23478_ (.A0(_19232_),
    .A1(\cpuregs[5][5] ),
    .S(_19649_),
    .X(_03000_));
 sky130_fd_sc_hd__mux2_2 _23479_ (.A0(_19233_),
    .A1(\cpuregs[5][4] ),
    .S(_19649_),
    .X(_02999_));
 sky130_fd_sc_hd__mux2_2 _23480_ (.A0(_19234_),
    .A1(\cpuregs[5][3] ),
    .S(_19649_),
    .X(_02998_));
 sky130_fd_sc_hd__mux2_2 _23481_ (.A0(_19235_),
    .A1(\cpuregs[5][2] ),
    .S(_19649_),
    .X(_02997_));
 sky130_fd_sc_hd__mux2_2 _23482_ (.A0(_19236_),
    .A1(\cpuregs[5][1] ),
    .S(_19644_),
    .X(_02996_));
 sky130_fd_sc_hd__mux2_2 _23483_ (.A0(_19237_),
    .A1(\cpuregs[5][0] ),
    .S(_19644_),
    .X(_02995_));
 sky130_fd_sc_hd__nand2_2 _23484_ (.A(_19080_),
    .B(_19238_),
    .Y(_19650_));
 sky130_fd_sc_hd__buf_1 _23485_ (.A(_19650_),
    .X(_19651_));
 sky130_fd_sc_hd__buf_1 _23486_ (.A(_19651_),
    .X(_19652_));
 sky130_fd_sc_hd__mux2_2 _23487_ (.A0(_19199_),
    .A1(\cpuregs[2][31] ),
    .S(_19652_),
    .X(_02994_));
 sky130_fd_sc_hd__mux2_2 _23488_ (.A0(_19203_),
    .A1(\cpuregs[2][30] ),
    .S(_19652_),
    .X(_02993_));
 sky130_fd_sc_hd__mux2_2 _23489_ (.A0(_19204_),
    .A1(\cpuregs[2][29] ),
    .S(_19652_),
    .X(_02992_));
 sky130_fd_sc_hd__mux2_2 _23490_ (.A0(_19205_),
    .A1(\cpuregs[2][28] ),
    .S(_19652_),
    .X(_02991_));
 sky130_fd_sc_hd__mux2_2 _23491_ (.A0(_19206_),
    .A1(\cpuregs[2][27] ),
    .S(_19652_),
    .X(_02990_));
 sky130_fd_sc_hd__mux2_2 _23492_ (.A0(_19207_),
    .A1(\cpuregs[2][26] ),
    .S(_19652_),
    .X(_02989_));
 sky130_fd_sc_hd__buf_1 _23493_ (.A(_19651_),
    .X(_19653_));
 sky130_fd_sc_hd__mux2_2 _23494_ (.A0(_19208_),
    .A1(\cpuregs[2][25] ),
    .S(_19653_),
    .X(_02988_));
 sky130_fd_sc_hd__mux2_2 _23495_ (.A0(_19210_),
    .A1(\cpuregs[2][24] ),
    .S(_19653_),
    .X(_02987_));
 sky130_fd_sc_hd__mux2_2 _23496_ (.A0(_19211_),
    .A1(\cpuregs[2][23] ),
    .S(_19653_),
    .X(_02986_));
 sky130_fd_sc_hd__mux2_2 _23497_ (.A0(_19212_),
    .A1(\cpuregs[2][22] ),
    .S(_19653_),
    .X(_02985_));
 sky130_fd_sc_hd__mux2_2 _23498_ (.A0(_19213_),
    .A1(\cpuregs[2][21] ),
    .S(_19653_),
    .X(_02984_));
 sky130_fd_sc_hd__mux2_2 _23499_ (.A0(_19214_),
    .A1(\cpuregs[2][20] ),
    .S(_19653_),
    .X(_02983_));
 sky130_fd_sc_hd__buf_1 _23500_ (.A(_19651_),
    .X(_19654_));
 sky130_fd_sc_hd__mux2_2 _23501_ (.A0(_19215_),
    .A1(\cpuregs[2][19] ),
    .S(_19654_),
    .X(_02982_));
 sky130_fd_sc_hd__mux2_2 _23502_ (.A0(_19217_),
    .A1(\cpuregs[2][18] ),
    .S(_19654_),
    .X(_02981_));
 sky130_fd_sc_hd__mux2_2 _23503_ (.A0(_19218_),
    .A1(\cpuregs[2][17] ),
    .S(_19654_),
    .X(_02980_));
 sky130_fd_sc_hd__mux2_2 _23504_ (.A0(_19219_),
    .A1(\cpuregs[2][16] ),
    .S(_19654_),
    .X(_02979_));
 sky130_fd_sc_hd__mux2_2 _23505_ (.A0(_19220_),
    .A1(\cpuregs[2][15] ),
    .S(_19654_),
    .X(_02978_));
 sky130_fd_sc_hd__mux2_2 _23506_ (.A0(_19221_),
    .A1(\cpuregs[2][14] ),
    .S(_19654_),
    .X(_02977_));
 sky130_fd_sc_hd__buf_1 _23507_ (.A(_19651_),
    .X(_19655_));
 sky130_fd_sc_hd__mux2_2 _23508_ (.A0(_19222_),
    .A1(\cpuregs[2][13] ),
    .S(_19655_),
    .X(_02976_));
 sky130_fd_sc_hd__mux2_2 _23509_ (.A0(_19224_),
    .A1(\cpuregs[2][12] ),
    .S(_19655_),
    .X(_02975_));
 sky130_fd_sc_hd__mux2_2 _23510_ (.A0(_19225_),
    .A1(\cpuregs[2][11] ),
    .S(_19655_),
    .X(_02974_));
 sky130_fd_sc_hd__mux2_2 _23511_ (.A0(_19226_),
    .A1(\cpuregs[2][10] ),
    .S(_19655_),
    .X(_02973_));
 sky130_fd_sc_hd__mux2_2 _23512_ (.A0(_19227_),
    .A1(\cpuregs[2][9] ),
    .S(_19655_),
    .X(_02972_));
 sky130_fd_sc_hd__mux2_2 _23513_ (.A0(_19228_),
    .A1(\cpuregs[2][8] ),
    .S(_19655_),
    .X(_02971_));
 sky130_fd_sc_hd__buf_1 _23514_ (.A(_19650_),
    .X(_19656_));
 sky130_fd_sc_hd__mux2_2 _23515_ (.A0(_19229_),
    .A1(\cpuregs[2][7] ),
    .S(_19656_),
    .X(_02970_));
 sky130_fd_sc_hd__mux2_2 _23516_ (.A0(_19231_),
    .A1(\cpuregs[2][6] ),
    .S(_19656_),
    .X(_02969_));
 sky130_fd_sc_hd__mux2_2 _23517_ (.A0(_19232_),
    .A1(\cpuregs[2][5] ),
    .S(_19656_),
    .X(_02968_));
 sky130_fd_sc_hd__mux2_2 _23518_ (.A0(_19233_),
    .A1(\cpuregs[2][4] ),
    .S(_19656_),
    .X(_02967_));
 sky130_fd_sc_hd__mux2_2 _23519_ (.A0(_19234_),
    .A1(\cpuregs[2][3] ),
    .S(_19656_),
    .X(_02966_));
 sky130_fd_sc_hd__mux2_2 _23520_ (.A0(_19235_),
    .A1(\cpuregs[2][2] ),
    .S(_19656_),
    .X(_02965_));
 sky130_fd_sc_hd__mux2_2 _23521_ (.A0(_19236_),
    .A1(\cpuregs[2][1] ),
    .S(_19651_),
    .X(_02964_));
 sky130_fd_sc_hd__mux2_2 _23522_ (.A0(_19237_),
    .A1(\cpuregs[2][0] ),
    .S(_19651_),
    .X(_02963_));
 sky130_fd_sc_hd__buf_1 _23523_ (.A(_18007_),
    .X(_19657_));
 sky130_fd_sc_hd__buf_1 _23524_ (.A(_19657_),
    .X(mem_xfer));
 sky130_fd_sc_hd__mux2_2 _23525_ (.A0(_19493_),
    .A1(mem_rdata[31]),
    .S(mem_xfer),
    .X(_02962_));
 sky130_fd_sc_hd__mux2_2 _23526_ (.A0(\mem_rdata_q[30] ),
    .A1(mem_rdata[30]),
    .S(mem_xfer),
    .X(_02961_));
 sky130_fd_sc_hd__mux2_2 _23527_ (.A0(\mem_rdata_q[29] ),
    .A1(mem_rdata[29]),
    .S(mem_xfer),
    .X(_02960_));
 sky130_fd_sc_hd__mux2_2 _23528_ (.A0(\mem_rdata_q[28] ),
    .A1(mem_rdata[28]),
    .S(mem_xfer),
    .X(_02959_));
 sky130_fd_sc_hd__mux2_2 _23529_ (.A0(\mem_rdata_q[27] ),
    .A1(mem_rdata[27]),
    .S(mem_xfer),
    .X(_02958_));
 sky130_fd_sc_hd__buf_1 _23530_ (.A(_19657_),
    .X(_19658_));
 sky130_fd_sc_hd__mux2_2 _23531_ (.A0(_19452_),
    .A1(mem_rdata[26]),
    .S(_19658_),
    .X(_02957_));
 sky130_fd_sc_hd__mux2_2 _23532_ (.A0(_19445_),
    .A1(mem_rdata[25]),
    .S(_19658_),
    .X(_02956_));
 sky130_fd_sc_hd__mux2_2 _23533_ (.A0(_19455_),
    .A1(mem_rdata[24]),
    .S(_19658_),
    .X(_02955_));
 sky130_fd_sc_hd__mux2_2 _23534_ (.A0(\mem_rdata_q[23] ),
    .A1(mem_rdata[23]),
    .S(_19658_),
    .X(_02954_));
 sky130_fd_sc_hd__mux2_2 _23535_ (.A0(\mem_rdata_q[22] ),
    .A1(mem_rdata[22]),
    .S(_19658_),
    .X(_02953_));
 sky130_fd_sc_hd__mux2_2 _23536_ (.A0(\mem_rdata_q[21] ),
    .A1(mem_rdata[21]),
    .S(_19658_),
    .X(_02952_));
 sky130_fd_sc_hd__buf_1 _23537_ (.A(_19657_),
    .X(_19659_));
 sky130_fd_sc_hd__mux2_2 _23538_ (.A0(\mem_rdata_q[20] ),
    .A1(mem_rdata[20]),
    .S(_19659_),
    .X(_02951_));
 sky130_fd_sc_hd__mux2_2 _23539_ (.A0(\mem_rdata_q[19] ),
    .A1(mem_rdata[19]),
    .S(_19659_),
    .X(_02950_));
 sky130_fd_sc_hd__mux2_2 _23540_ (.A0(\mem_rdata_q[18] ),
    .A1(mem_rdata[18]),
    .S(_19659_),
    .X(_02949_));
 sky130_fd_sc_hd__mux2_2 _23541_ (.A0(\mem_rdata_q[17] ),
    .A1(mem_rdata[17]),
    .S(_19659_),
    .X(_02948_));
 sky130_fd_sc_hd__mux2_2 _23542_ (.A0(\mem_rdata_q[16] ),
    .A1(mem_rdata[16]),
    .S(_19659_),
    .X(_02947_));
 sky130_fd_sc_hd__mux2_2 _23543_ (.A0(\mem_rdata_q[15] ),
    .A1(mem_rdata[15]),
    .S(_19659_),
    .X(_02946_));
 sky130_fd_sc_hd__buf_1 _23544_ (.A(_18007_),
    .X(_19660_));
 sky130_fd_sc_hd__mux2_2 _23545_ (.A0(_18379_),
    .A1(mem_rdata[14]),
    .S(_19660_),
    .X(_02945_));
 sky130_fd_sc_hd__mux2_2 _23546_ (.A0(\mem_rdata_q[13] ),
    .A1(mem_rdata[13]),
    .S(_19660_),
    .X(_02944_));
 sky130_fd_sc_hd__mux2_2 _23547_ (.A0(_18398_),
    .A1(mem_rdata[12]),
    .S(_19660_),
    .X(_02943_));
 sky130_fd_sc_hd__mux2_2 _23548_ (.A0(\mem_rdata_q[11] ),
    .A1(mem_rdata[11]),
    .S(_19660_),
    .X(_02942_));
 sky130_fd_sc_hd__mux2_2 _23549_ (.A0(\mem_rdata_q[10] ),
    .A1(mem_rdata[10]),
    .S(_19660_),
    .X(_02941_));
 sky130_fd_sc_hd__mux2_2 _23550_ (.A0(\mem_rdata_q[9] ),
    .A1(mem_rdata[9]),
    .S(_19660_),
    .X(_02940_));
 sky130_fd_sc_hd__buf_1 _23551_ (.A(_18007_),
    .X(_19661_));
 sky130_fd_sc_hd__mux2_2 _23552_ (.A0(\mem_rdata_q[8] ),
    .A1(mem_rdata[8]),
    .S(_19661_),
    .X(_02939_));
 sky130_fd_sc_hd__mux2_2 _23553_ (.A0(\mem_rdata_q[7] ),
    .A1(mem_rdata[7]),
    .S(_19661_),
    .X(_02938_));
 sky130_fd_sc_hd__mux2_2 _23554_ (.A0(\mem_rdata_q[6] ),
    .A1(mem_rdata[6]),
    .S(_19661_),
    .X(_02937_));
 sky130_fd_sc_hd__mux2_2 _23555_ (.A0(\mem_rdata_q[5] ),
    .A1(mem_rdata[5]),
    .S(_19661_),
    .X(_02936_));
 sky130_fd_sc_hd__mux2_2 _23556_ (.A0(\mem_rdata_q[4] ),
    .A1(mem_rdata[4]),
    .S(_19661_),
    .X(_02935_));
 sky130_fd_sc_hd__mux2_2 _23557_ (.A0(\mem_rdata_q[3] ),
    .A1(mem_rdata[3]),
    .S(_19661_),
    .X(_02934_));
 sky130_fd_sc_hd__mux2_2 _23558_ (.A0(\mem_rdata_q[2] ),
    .A1(mem_rdata[2]),
    .S(_19657_),
    .X(_02933_));
 sky130_fd_sc_hd__mux2_2 _23559_ (.A0(\mem_rdata_q[1] ),
    .A1(mem_rdata[1]),
    .S(_19657_),
    .X(_02932_));
 sky130_fd_sc_hd__mux2_2 _23560_ (.A0(\mem_rdata_q[0] ),
    .A1(mem_rdata[0]),
    .S(_19657_),
    .X(_02931_));
 sky130_fd_sc_hd__nand2_2 _23561_ (.A(_19080_),
    .B(_19165_),
    .Y(_19662_));
 sky130_fd_sc_hd__buf_1 _23562_ (.A(_19662_),
    .X(_19663_));
 sky130_fd_sc_hd__buf_1 _23563_ (.A(_19663_),
    .X(_19664_));
 sky130_fd_sc_hd__mux2_2 _23564_ (.A0(_19199_),
    .A1(\cpuregs[18][31] ),
    .S(_19664_),
    .X(_02930_));
 sky130_fd_sc_hd__mux2_2 _23565_ (.A0(_19203_),
    .A1(\cpuregs[18][30] ),
    .S(_19664_),
    .X(_02929_));
 sky130_fd_sc_hd__mux2_2 _23566_ (.A0(_19204_),
    .A1(\cpuregs[18][29] ),
    .S(_19664_),
    .X(_02928_));
 sky130_fd_sc_hd__mux2_2 _23567_ (.A0(_19205_),
    .A1(\cpuregs[18][28] ),
    .S(_19664_),
    .X(_02927_));
 sky130_fd_sc_hd__mux2_2 _23568_ (.A0(_19206_),
    .A1(\cpuregs[18][27] ),
    .S(_19664_),
    .X(_02926_));
 sky130_fd_sc_hd__mux2_2 _23569_ (.A0(_19207_),
    .A1(\cpuregs[18][26] ),
    .S(_19664_),
    .X(_02925_));
 sky130_fd_sc_hd__buf_1 _23570_ (.A(_19663_),
    .X(_19665_));
 sky130_fd_sc_hd__mux2_2 _23571_ (.A0(_19208_),
    .A1(\cpuregs[18][25] ),
    .S(_19665_),
    .X(_02924_));
 sky130_fd_sc_hd__mux2_2 _23572_ (.A0(_19210_),
    .A1(\cpuregs[18][24] ),
    .S(_19665_),
    .X(_02923_));
 sky130_fd_sc_hd__mux2_2 _23573_ (.A0(_19211_),
    .A1(\cpuregs[18][23] ),
    .S(_19665_),
    .X(_02922_));
 sky130_fd_sc_hd__mux2_2 _23574_ (.A0(_19212_),
    .A1(\cpuregs[18][22] ),
    .S(_19665_),
    .X(_02921_));
 sky130_fd_sc_hd__mux2_2 _23575_ (.A0(_19213_),
    .A1(\cpuregs[18][21] ),
    .S(_19665_),
    .X(_02920_));
 sky130_fd_sc_hd__mux2_2 _23576_ (.A0(_19214_),
    .A1(\cpuregs[18][20] ),
    .S(_19665_),
    .X(_02919_));
 sky130_fd_sc_hd__buf_1 _23577_ (.A(_19663_),
    .X(_19666_));
 sky130_fd_sc_hd__mux2_2 _23578_ (.A0(_19215_),
    .A1(\cpuregs[18][19] ),
    .S(_19666_),
    .X(_02918_));
 sky130_fd_sc_hd__mux2_2 _23579_ (.A0(_19217_),
    .A1(\cpuregs[18][18] ),
    .S(_19666_),
    .X(_02917_));
 sky130_fd_sc_hd__mux2_2 _23580_ (.A0(_19218_),
    .A1(\cpuregs[18][17] ),
    .S(_19666_),
    .X(_02916_));
 sky130_fd_sc_hd__mux2_2 _23581_ (.A0(_19219_),
    .A1(\cpuregs[18][16] ),
    .S(_19666_),
    .X(_02915_));
 sky130_fd_sc_hd__mux2_2 _23582_ (.A0(_19220_),
    .A1(\cpuregs[18][15] ),
    .S(_19666_),
    .X(_02914_));
 sky130_fd_sc_hd__mux2_2 _23583_ (.A0(_19221_),
    .A1(\cpuregs[18][14] ),
    .S(_19666_),
    .X(_02913_));
 sky130_fd_sc_hd__buf_1 _23584_ (.A(_19663_),
    .X(_19667_));
 sky130_fd_sc_hd__mux2_2 _23585_ (.A0(_19222_),
    .A1(\cpuregs[18][13] ),
    .S(_19667_),
    .X(_02912_));
 sky130_fd_sc_hd__mux2_2 _23586_ (.A0(_19224_),
    .A1(\cpuregs[18][12] ),
    .S(_19667_),
    .X(_02911_));
 sky130_fd_sc_hd__mux2_2 _23587_ (.A0(_19225_),
    .A1(\cpuregs[18][11] ),
    .S(_19667_),
    .X(_02910_));
 sky130_fd_sc_hd__mux2_2 _23588_ (.A0(_19226_),
    .A1(\cpuregs[18][10] ),
    .S(_19667_),
    .X(_02909_));
 sky130_fd_sc_hd__mux2_2 _23589_ (.A0(_19227_),
    .A1(\cpuregs[18][9] ),
    .S(_19667_),
    .X(_02908_));
 sky130_fd_sc_hd__mux2_2 _23590_ (.A0(_19228_),
    .A1(\cpuregs[18][8] ),
    .S(_19667_),
    .X(_02907_));
 sky130_fd_sc_hd__buf_1 _23591_ (.A(_19662_),
    .X(_19668_));
 sky130_fd_sc_hd__mux2_2 _23592_ (.A0(_19229_),
    .A1(\cpuregs[18][7] ),
    .S(_19668_),
    .X(_02906_));
 sky130_fd_sc_hd__mux2_2 _23593_ (.A0(_19231_),
    .A1(\cpuregs[18][6] ),
    .S(_19668_),
    .X(_02905_));
 sky130_fd_sc_hd__mux2_2 _23594_ (.A0(_19232_),
    .A1(\cpuregs[18][5] ),
    .S(_19668_),
    .X(_02904_));
 sky130_fd_sc_hd__mux2_2 _23595_ (.A0(_19233_),
    .A1(\cpuregs[18][4] ),
    .S(_19668_),
    .X(_02903_));
 sky130_fd_sc_hd__mux2_2 _23596_ (.A0(_19234_),
    .A1(\cpuregs[18][3] ),
    .S(_19668_),
    .X(_02902_));
 sky130_fd_sc_hd__mux2_2 _23597_ (.A0(_19235_),
    .A1(\cpuregs[18][2] ),
    .S(_19668_),
    .X(_02901_));
 sky130_fd_sc_hd__mux2_2 _23598_ (.A0(_19236_),
    .A1(\cpuregs[18][1] ),
    .S(_19663_),
    .X(_02900_));
 sky130_fd_sc_hd__mux2_2 _23599_ (.A0(_19237_),
    .A1(\cpuregs[18][0] ),
    .S(_19663_),
    .X(_02899_));
 sky130_fd_sc_hd__nand2_2 _23600_ (.A(_19080_),
    .B(_19123_),
    .Y(_19669_));
 sky130_fd_sc_hd__buf_1 _23601_ (.A(_19669_),
    .X(_19670_));
 sky130_fd_sc_hd__buf_1 _23602_ (.A(_19670_),
    .X(_19671_));
 sky130_fd_sc_hd__mux2_2 _23603_ (.A0(_19246_),
    .A1(\cpuregs[10][31] ),
    .S(_19671_),
    .X(_02898_));
 sky130_fd_sc_hd__mux2_2 _23604_ (.A0(_19250_),
    .A1(\cpuregs[10][30] ),
    .S(_19671_),
    .X(_02897_));
 sky130_fd_sc_hd__mux2_2 _23605_ (.A0(_19251_),
    .A1(\cpuregs[10][29] ),
    .S(_19671_),
    .X(_02896_));
 sky130_fd_sc_hd__mux2_2 _23606_ (.A0(_19252_),
    .A1(\cpuregs[10][28] ),
    .S(_19671_),
    .X(_02895_));
 sky130_fd_sc_hd__mux2_2 _23607_ (.A0(_19253_),
    .A1(\cpuregs[10][27] ),
    .S(_19671_),
    .X(_02894_));
 sky130_fd_sc_hd__mux2_2 _23608_ (.A0(_19254_),
    .A1(\cpuregs[10][26] ),
    .S(_19671_),
    .X(_02893_));
 sky130_fd_sc_hd__buf_1 _23609_ (.A(_19670_),
    .X(_19672_));
 sky130_fd_sc_hd__mux2_2 _23610_ (.A0(_19255_),
    .A1(\cpuregs[10][25] ),
    .S(_19672_),
    .X(_02892_));
 sky130_fd_sc_hd__mux2_2 _23611_ (.A0(_19257_),
    .A1(\cpuregs[10][24] ),
    .S(_19672_),
    .X(_02891_));
 sky130_fd_sc_hd__mux2_2 _23612_ (.A0(_19258_),
    .A1(\cpuregs[10][23] ),
    .S(_19672_),
    .X(_02890_));
 sky130_fd_sc_hd__mux2_2 _23613_ (.A0(_19259_),
    .A1(\cpuregs[10][22] ),
    .S(_19672_),
    .X(_02889_));
 sky130_fd_sc_hd__mux2_2 _23614_ (.A0(_19260_),
    .A1(\cpuregs[10][21] ),
    .S(_19672_),
    .X(_02888_));
 sky130_fd_sc_hd__mux2_2 _23615_ (.A0(_19261_),
    .A1(\cpuregs[10][20] ),
    .S(_19672_),
    .X(_02887_));
 sky130_fd_sc_hd__buf_1 _23616_ (.A(_19670_),
    .X(_19673_));
 sky130_fd_sc_hd__mux2_2 _23617_ (.A0(_19262_),
    .A1(\cpuregs[10][19] ),
    .S(_19673_),
    .X(_02886_));
 sky130_fd_sc_hd__mux2_2 _23618_ (.A0(_19264_),
    .A1(\cpuregs[10][18] ),
    .S(_19673_),
    .X(_02885_));
 sky130_fd_sc_hd__mux2_2 _23619_ (.A0(_19265_),
    .A1(\cpuregs[10][17] ),
    .S(_19673_),
    .X(_02884_));
 sky130_fd_sc_hd__mux2_2 _23620_ (.A0(_19266_),
    .A1(\cpuregs[10][16] ),
    .S(_19673_),
    .X(_02883_));
 sky130_fd_sc_hd__mux2_2 _23621_ (.A0(_19267_),
    .A1(\cpuregs[10][15] ),
    .S(_19673_),
    .X(_02882_));
 sky130_fd_sc_hd__mux2_2 _23622_ (.A0(_19268_),
    .A1(\cpuregs[10][14] ),
    .S(_19673_),
    .X(_02881_));
 sky130_fd_sc_hd__buf_1 _23623_ (.A(_19670_),
    .X(_19674_));
 sky130_fd_sc_hd__mux2_2 _23624_ (.A0(_19269_),
    .A1(\cpuregs[10][13] ),
    .S(_19674_),
    .X(_02880_));
 sky130_fd_sc_hd__mux2_2 _23625_ (.A0(_19271_),
    .A1(\cpuregs[10][12] ),
    .S(_19674_),
    .X(_02879_));
 sky130_fd_sc_hd__mux2_2 _23626_ (.A0(_19272_),
    .A1(\cpuregs[10][11] ),
    .S(_19674_),
    .X(_02878_));
 sky130_fd_sc_hd__mux2_2 _23627_ (.A0(_19273_),
    .A1(\cpuregs[10][10] ),
    .S(_19674_),
    .X(_02877_));
 sky130_fd_sc_hd__mux2_2 _23628_ (.A0(_19274_),
    .A1(\cpuregs[10][9] ),
    .S(_19674_),
    .X(_02876_));
 sky130_fd_sc_hd__mux2_2 _23629_ (.A0(_19275_),
    .A1(\cpuregs[10][8] ),
    .S(_19674_),
    .X(_02875_));
 sky130_fd_sc_hd__buf_1 _23630_ (.A(_19669_),
    .X(_19675_));
 sky130_fd_sc_hd__mux2_2 _23631_ (.A0(_19276_),
    .A1(\cpuregs[10][7] ),
    .S(_19675_),
    .X(_02874_));
 sky130_fd_sc_hd__mux2_2 _23632_ (.A0(_19278_),
    .A1(\cpuregs[10][6] ),
    .S(_19675_),
    .X(_02873_));
 sky130_fd_sc_hd__mux2_2 _23633_ (.A0(_19279_),
    .A1(\cpuregs[10][5] ),
    .S(_19675_),
    .X(_02872_));
 sky130_fd_sc_hd__mux2_2 _23634_ (.A0(_19280_),
    .A1(\cpuregs[10][4] ),
    .S(_19675_),
    .X(_02871_));
 sky130_fd_sc_hd__mux2_2 _23635_ (.A0(_19281_),
    .A1(\cpuregs[10][3] ),
    .S(_19675_),
    .X(_02870_));
 sky130_fd_sc_hd__mux2_2 _23636_ (.A0(_19282_),
    .A1(\cpuregs[10][2] ),
    .S(_19675_),
    .X(_02869_));
 sky130_fd_sc_hd__mux2_2 _23637_ (.A0(_19283_),
    .A1(\cpuregs[10][1] ),
    .S(_19670_),
    .X(_02868_));
 sky130_fd_sc_hd__mux2_2 _23638_ (.A0(_19284_),
    .A1(\cpuregs[10][0] ),
    .S(_19670_),
    .X(_02867_));
 sky130_fd_sc_hd__buf_1 _23639_ (.A(\cpuregs[0][31] ),
    .X(_02866_));
 sky130_fd_sc_hd__buf_1 _23640_ (.A(\cpuregs[0][30] ),
    .X(_02865_));
 sky130_fd_sc_hd__buf_1 _23641_ (.A(\cpuregs[0][29] ),
    .X(_02864_));
 sky130_fd_sc_hd__buf_1 _23642_ (.A(\cpuregs[0][28] ),
    .X(_02863_));
 sky130_fd_sc_hd__buf_1 _23643_ (.A(\cpuregs[0][27] ),
    .X(_02862_));
 sky130_fd_sc_hd__buf_1 _23644_ (.A(\cpuregs[0][26] ),
    .X(_02861_));
 sky130_fd_sc_hd__buf_1 _23645_ (.A(\cpuregs[0][25] ),
    .X(_02860_));
 sky130_fd_sc_hd__buf_1 _23646_ (.A(\cpuregs[0][24] ),
    .X(_02859_));
 sky130_fd_sc_hd__buf_1 _23647_ (.A(\cpuregs[0][23] ),
    .X(_02858_));
 sky130_fd_sc_hd__buf_1 _23648_ (.A(\cpuregs[0][22] ),
    .X(_02857_));
 sky130_fd_sc_hd__buf_1 _23649_ (.A(\cpuregs[0][21] ),
    .X(_02856_));
 sky130_fd_sc_hd__buf_1 _23650_ (.A(\cpuregs[0][20] ),
    .X(_02855_));
 sky130_fd_sc_hd__buf_1 _23651_ (.A(\cpuregs[0][19] ),
    .X(_02854_));
 sky130_fd_sc_hd__buf_1 _23652_ (.A(\cpuregs[0][18] ),
    .X(_02853_));
 sky130_fd_sc_hd__buf_1 _23653_ (.A(\cpuregs[0][17] ),
    .X(_02852_));
 sky130_fd_sc_hd__buf_1 _23654_ (.A(\cpuregs[0][16] ),
    .X(_02851_));
 sky130_fd_sc_hd__buf_1 _23655_ (.A(\cpuregs[0][15] ),
    .X(_02850_));
 sky130_fd_sc_hd__buf_1 _23656_ (.A(\cpuregs[0][14] ),
    .X(_02849_));
 sky130_fd_sc_hd__buf_1 _23657_ (.A(\cpuregs[0][13] ),
    .X(_02848_));
 sky130_fd_sc_hd__buf_1 _23658_ (.A(\cpuregs[0][12] ),
    .X(_02847_));
 sky130_fd_sc_hd__buf_1 _23659_ (.A(\cpuregs[0][11] ),
    .X(_02846_));
 sky130_fd_sc_hd__buf_1 _23660_ (.A(\cpuregs[0][10] ),
    .X(_02845_));
 sky130_fd_sc_hd__buf_1 _23661_ (.A(\cpuregs[0][9] ),
    .X(_02844_));
 sky130_fd_sc_hd__buf_1 _23662_ (.A(\cpuregs[0][8] ),
    .X(_02843_));
 sky130_fd_sc_hd__buf_1 _23663_ (.A(\cpuregs[0][7] ),
    .X(_02842_));
 sky130_fd_sc_hd__buf_1 _23664_ (.A(\cpuregs[0][6] ),
    .X(_02841_));
 sky130_fd_sc_hd__buf_1 _23665_ (.A(\cpuregs[0][5] ),
    .X(_02840_));
 sky130_fd_sc_hd__buf_1 _23666_ (.A(\cpuregs[0][4] ),
    .X(_02839_));
 sky130_fd_sc_hd__buf_1 _23667_ (.A(\cpuregs[0][3] ),
    .X(_02838_));
 sky130_fd_sc_hd__buf_1 _23668_ (.A(\cpuregs[0][2] ),
    .X(_02837_));
 sky130_fd_sc_hd__buf_1 _23669_ (.A(\cpuregs[0][1] ),
    .X(_02836_));
 sky130_fd_sc_hd__buf_1 _23670_ (.A(\cpuregs[0][0] ),
    .X(_02835_));
 sky130_fd_sc_hd__nand2_2 _23671_ (.A(_19080_),
    .B(_19191_),
    .Y(_19676_));
 sky130_fd_sc_hd__buf_1 _23672_ (.A(_19676_),
    .X(_19677_));
 sky130_fd_sc_hd__buf_1 _23673_ (.A(_19677_),
    .X(_19678_));
 sky130_fd_sc_hd__mux2_2 _23674_ (.A0(_19246_),
    .A1(\cpuregs[14][31] ),
    .S(_19678_),
    .X(_02834_));
 sky130_fd_sc_hd__mux2_2 _23675_ (.A0(_19250_),
    .A1(\cpuregs[14][30] ),
    .S(_19678_),
    .X(_02833_));
 sky130_fd_sc_hd__mux2_2 _23676_ (.A0(_19251_),
    .A1(\cpuregs[14][29] ),
    .S(_19678_),
    .X(_02832_));
 sky130_fd_sc_hd__mux2_2 _23677_ (.A0(_19252_),
    .A1(\cpuregs[14][28] ),
    .S(_19678_),
    .X(_02831_));
 sky130_fd_sc_hd__mux2_2 _23678_ (.A0(_19253_),
    .A1(\cpuregs[14][27] ),
    .S(_19678_),
    .X(_02830_));
 sky130_fd_sc_hd__mux2_2 _23679_ (.A0(_19254_),
    .A1(\cpuregs[14][26] ),
    .S(_19678_),
    .X(_02829_));
 sky130_fd_sc_hd__buf_1 _23680_ (.A(_19677_),
    .X(_19679_));
 sky130_fd_sc_hd__mux2_2 _23681_ (.A0(_19255_),
    .A1(\cpuregs[14][25] ),
    .S(_19679_),
    .X(_02828_));
 sky130_fd_sc_hd__mux2_2 _23682_ (.A0(_19257_),
    .A1(\cpuregs[14][24] ),
    .S(_19679_),
    .X(_02827_));
 sky130_fd_sc_hd__mux2_2 _23683_ (.A0(_19258_),
    .A1(\cpuregs[14][23] ),
    .S(_19679_),
    .X(_02826_));
 sky130_fd_sc_hd__mux2_2 _23684_ (.A0(_19259_),
    .A1(\cpuregs[14][22] ),
    .S(_19679_),
    .X(_02825_));
 sky130_fd_sc_hd__mux2_2 _23685_ (.A0(_19260_),
    .A1(\cpuregs[14][21] ),
    .S(_19679_),
    .X(_02824_));
 sky130_fd_sc_hd__mux2_2 _23686_ (.A0(_19261_),
    .A1(\cpuregs[14][20] ),
    .S(_19679_),
    .X(_02823_));
 sky130_fd_sc_hd__buf_1 _23687_ (.A(_19677_),
    .X(_19680_));
 sky130_fd_sc_hd__mux2_2 _23688_ (.A0(_19262_),
    .A1(\cpuregs[14][19] ),
    .S(_19680_),
    .X(_02822_));
 sky130_fd_sc_hd__mux2_2 _23689_ (.A0(_19264_),
    .A1(\cpuregs[14][18] ),
    .S(_19680_),
    .X(_02821_));
 sky130_fd_sc_hd__mux2_2 _23690_ (.A0(_19265_),
    .A1(\cpuregs[14][17] ),
    .S(_19680_),
    .X(_02820_));
 sky130_fd_sc_hd__mux2_2 _23691_ (.A0(_19266_),
    .A1(\cpuregs[14][16] ),
    .S(_19680_),
    .X(_02819_));
 sky130_fd_sc_hd__mux2_2 _23692_ (.A0(_19267_),
    .A1(\cpuregs[14][15] ),
    .S(_19680_),
    .X(_02818_));
 sky130_fd_sc_hd__mux2_2 _23693_ (.A0(_19268_),
    .A1(\cpuregs[14][14] ),
    .S(_19680_),
    .X(_02817_));
 sky130_fd_sc_hd__buf_1 _23694_ (.A(_19677_),
    .X(_19681_));
 sky130_fd_sc_hd__mux2_2 _23695_ (.A0(_19269_),
    .A1(\cpuregs[14][13] ),
    .S(_19681_),
    .X(_02816_));
 sky130_fd_sc_hd__mux2_2 _23696_ (.A0(_19271_),
    .A1(\cpuregs[14][12] ),
    .S(_19681_),
    .X(_02815_));
 sky130_fd_sc_hd__mux2_2 _23697_ (.A0(_19272_),
    .A1(\cpuregs[14][11] ),
    .S(_19681_),
    .X(_02814_));
 sky130_fd_sc_hd__mux2_2 _23698_ (.A0(_19273_),
    .A1(\cpuregs[14][10] ),
    .S(_19681_),
    .X(_02813_));
 sky130_fd_sc_hd__mux2_2 _23699_ (.A0(_19274_),
    .A1(\cpuregs[14][9] ),
    .S(_19681_),
    .X(_02812_));
 sky130_fd_sc_hd__mux2_2 _23700_ (.A0(_19275_),
    .A1(\cpuregs[14][8] ),
    .S(_19681_),
    .X(_02811_));
 sky130_fd_sc_hd__buf_1 _23701_ (.A(_19676_),
    .X(_19682_));
 sky130_fd_sc_hd__mux2_2 _23702_ (.A0(_19276_),
    .A1(\cpuregs[14][7] ),
    .S(_19682_),
    .X(_02810_));
 sky130_fd_sc_hd__mux2_2 _23703_ (.A0(_19278_),
    .A1(\cpuregs[14][6] ),
    .S(_19682_),
    .X(_02809_));
 sky130_fd_sc_hd__mux2_2 _23704_ (.A0(_19279_),
    .A1(\cpuregs[14][5] ),
    .S(_19682_),
    .X(_02808_));
 sky130_fd_sc_hd__mux2_2 _23705_ (.A0(_19280_),
    .A1(\cpuregs[14][4] ),
    .S(_19682_),
    .X(_02807_));
 sky130_fd_sc_hd__mux2_2 _23706_ (.A0(_19281_),
    .A1(\cpuregs[14][3] ),
    .S(_19682_),
    .X(_02806_));
 sky130_fd_sc_hd__mux2_2 _23707_ (.A0(_19282_),
    .A1(\cpuregs[14][2] ),
    .S(_19682_),
    .X(_02805_));
 sky130_fd_sc_hd__mux2_2 _23708_ (.A0(_19283_),
    .A1(\cpuregs[14][1] ),
    .S(_19677_),
    .X(_02804_));
 sky130_fd_sc_hd__mux2_2 _23709_ (.A0(_19284_),
    .A1(\cpuregs[14][0] ),
    .S(_19677_),
    .X(_02803_));
 sky130_fd_sc_hd__or3_2 _23710_ (.A(_19071_),
    .B(_19122_),
    .C(_19078_),
    .X(_19683_));
 sky130_fd_sc_hd__buf_1 _23711_ (.A(_19683_),
    .X(_19684_));
 sky130_fd_sc_hd__buf_1 _23712_ (.A(_19684_),
    .X(_19685_));
 sky130_fd_sc_hd__mux2_2 _23713_ (.A0(_19246_),
    .A1(\cpuregs[8][31] ),
    .S(_19685_),
    .X(_02802_));
 sky130_fd_sc_hd__mux2_2 _23714_ (.A0(_19250_),
    .A1(\cpuregs[8][30] ),
    .S(_19685_),
    .X(_02801_));
 sky130_fd_sc_hd__mux2_2 _23715_ (.A0(_19251_),
    .A1(\cpuregs[8][29] ),
    .S(_19685_),
    .X(_02800_));
 sky130_fd_sc_hd__mux2_2 _23716_ (.A0(_19252_),
    .A1(\cpuregs[8][28] ),
    .S(_19685_),
    .X(_02799_));
 sky130_fd_sc_hd__mux2_2 _23717_ (.A0(_19253_),
    .A1(\cpuregs[8][27] ),
    .S(_19685_),
    .X(_02798_));
 sky130_fd_sc_hd__mux2_2 _23718_ (.A0(_19254_),
    .A1(\cpuregs[8][26] ),
    .S(_19685_),
    .X(_02797_));
 sky130_fd_sc_hd__buf_1 _23719_ (.A(_19684_),
    .X(_19686_));
 sky130_fd_sc_hd__mux2_2 _23720_ (.A0(_19255_),
    .A1(\cpuregs[8][25] ),
    .S(_19686_),
    .X(_02796_));
 sky130_fd_sc_hd__mux2_2 _23721_ (.A0(_19257_),
    .A1(\cpuregs[8][24] ),
    .S(_19686_),
    .X(_02795_));
 sky130_fd_sc_hd__mux2_2 _23722_ (.A0(_19258_),
    .A1(\cpuregs[8][23] ),
    .S(_19686_),
    .X(_02794_));
 sky130_fd_sc_hd__mux2_2 _23723_ (.A0(_19259_),
    .A1(\cpuregs[8][22] ),
    .S(_19686_),
    .X(_02793_));
 sky130_fd_sc_hd__mux2_2 _23724_ (.A0(_19260_),
    .A1(\cpuregs[8][21] ),
    .S(_19686_),
    .X(_02792_));
 sky130_fd_sc_hd__mux2_2 _23725_ (.A0(_19261_),
    .A1(\cpuregs[8][20] ),
    .S(_19686_),
    .X(_02791_));
 sky130_fd_sc_hd__buf_1 _23726_ (.A(_19684_),
    .X(_19687_));
 sky130_fd_sc_hd__mux2_2 _23727_ (.A0(_19262_),
    .A1(\cpuregs[8][19] ),
    .S(_19687_),
    .X(_02790_));
 sky130_fd_sc_hd__mux2_2 _23728_ (.A0(_19264_),
    .A1(\cpuregs[8][18] ),
    .S(_19687_),
    .X(_02789_));
 sky130_fd_sc_hd__mux2_2 _23729_ (.A0(_19265_),
    .A1(\cpuregs[8][17] ),
    .S(_19687_),
    .X(_02788_));
 sky130_fd_sc_hd__mux2_2 _23730_ (.A0(_19266_),
    .A1(\cpuregs[8][16] ),
    .S(_19687_),
    .X(_02787_));
 sky130_fd_sc_hd__mux2_2 _23731_ (.A0(_19267_),
    .A1(\cpuregs[8][15] ),
    .S(_19687_),
    .X(_02786_));
 sky130_fd_sc_hd__mux2_2 _23732_ (.A0(_19268_),
    .A1(\cpuregs[8][14] ),
    .S(_19687_),
    .X(_02785_));
 sky130_fd_sc_hd__buf_1 _23733_ (.A(_19684_),
    .X(_19688_));
 sky130_fd_sc_hd__mux2_2 _23734_ (.A0(_19269_),
    .A1(\cpuregs[8][13] ),
    .S(_19688_),
    .X(_02784_));
 sky130_fd_sc_hd__mux2_2 _23735_ (.A0(_19271_),
    .A1(\cpuregs[8][12] ),
    .S(_19688_),
    .X(_02783_));
 sky130_fd_sc_hd__mux2_2 _23736_ (.A0(_19272_),
    .A1(\cpuregs[8][11] ),
    .S(_19688_),
    .X(_02782_));
 sky130_fd_sc_hd__mux2_2 _23737_ (.A0(_19273_),
    .A1(\cpuregs[8][10] ),
    .S(_19688_),
    .X(_02781_));
 sky130_fd_sc_hd__mux2_2 _23738_ (.A0(_19274_),
    .A1(\cpuregs[8][9] ),
    .S(_19688_),
    .X(_02780_));
 sky130_fd_sc_hd__mux2_2 _23739_ (.A0(_19275_),
    .A1(\cpuregs[8][8] ),
    .S(_19688_),
    .X(_02779_));
 sky130_fd_sc_hd__buf_1 _23740_ (.A(_19683_),
    .X(_19689_));
 sky130_fd_sc_hd__mux2_2 _23741_ (.A0(_19276_),
    .A1(\cpuregs[8][7] ),
    .S(_19689_),
    .X(_02778_));
 sky130_fd_sc_hd__mux2_2 _23742_ (.A0(_19278_),
    .A1(\cpuregs[8][6] ),
    .S(_19689_),
    .X(_02777_));
 sky130_fd_sc_hd__mux2_2 _23743_ (.A0(_19279_),
    .A1(\cpuregs[8][5] ),
    .S(_19689_),
    .X(_02776_));
 sky130_fd_sc_hd__mux2_2 _23744_ (.A0(_19280_),
    .A1(\cpuregs[8][4] ),
    .S(_19689_),
    .X(_02775_));
 sky130_fd_sc_hd__mux2_2 _23745_ (.A0(_19281_),
    .A1(\cpuregs[8][3] ),
    .S(_19689_),
    .X(_02774_));
 sky130_fd_sc_hd__mux2_2 _23746_ (.A0(_19282_),
    .A1(\cpuregs[8][2] ),
    .S(_19689_),
    .X(_02773_));
 sky130_fd_sc_hd__mux2_2 _23747_ (.A0(_19283_),
    .A1(\cpuregs[8][1] ),
    .S(_19684_),
    .X(_02772_));
 sky130_fd_sc_hd__mux2_2 _23748_ (.A0(_19284_),
    .A1(\cpuregs[8][0] ),
    .S(_19684_),
    .X(_02771_));
 sky130_fd_sc_hd__nor2_2 _23749_ (.A(latched_branch),
    .B(_18240_),
    .Y(_00292_));
 sky130_fd_sc_hd__nor2_2 _23750_ (.A(latched_store),
    .B(_18037_),
    .Y(_19690_));
 sky130_fd_sc_hd__o311a_2 _23751_ (.A1(_18494_),
    .A2(_00292_),
    .A3(_19690_),
    .B1(_18407_),
    .C1(\reg_next_pc[0] ),
    .X(_02770_));
 sky130_fd_sc_hd__and2_2 _23752_ (.A(_18885_),
    .B(_00008_),
    .X(_02769_));
 sky130_fd_sc_hd__and2_2 _23753_ (.A(_18885_),
    .B(_20622_),
    .X(_02768_));
 sky130_fd_sc_hd__and2_2 _23754_ (.A(_18885_),
    .B(_00031_),
    .X(_02767_));
 sky130_fd_sc_hd__buf_1 _23755_ (.A(_18395_),
    .X(_19691_));
 sky130_fd_sc_hd__and2_2 _23756_ (.A(_19691_),
    .B(_00032_),
    .X(_02766_));
 sky130_fd_sc_hd__and2_2 _23757_ (.A(_19691_),
    .B(_00033_),
    .X(_02765_));
 sky130_fd_sc_hd__and2_2 _23758_ (.A(_19691_),
    .B(_00034_),
    .X(_02764_));
 sky130_fd_sc_hd__and2_2 _23759_ (.A(_19691_),
    .B(_00035_),
    .X(_02763_));
 sky130_fd_sc_hd__and2_2 _23760_ (.A(_19691_),
    .B(_00036_),
    .X(_02762_));
 sky130_fd_sc_hd__and2_2 _23761_ (.A(_19691_),
    .B(_00037_),
    .X(_02761_));
 sky130_fd_sc_hd__buf_1 _23762_ (.A(_18395_),
    .X(_19692_));
 sky130_fd_sc_hd__and2_2 _23763_ (.A(_19692_),
    .B(_00009_),
    .X(_02760_));
 sky130_fd_sc_hd__and2_2 _23764_ (.A(_19692_),
    .B(_00010_),
    .X(_02759_));
 sky130_fd_sc_hd__and2_2 _23765_ (.A(_19692_),
    .B(_00011_),
    .X(_02758_));
 sky130_fd_sc_hd__and2_2 _23766_ (.A(_19692_),
    .B(_00012_),
    .X(_02757_));
 sky130_fd_sc_hd__and2_2 _23767_ (.A(_19692_),
    .B(_00013_),
    .X(_02756_));
 sky130_fd_sc_hd__and2_2 _23768_ (.A(_19692_),
    .B(_00014_),
    .X(_02755_));
 sky130_fd_sc_hd__buf_1 _23769_ (.A(_18395_),
    .X(_19693_));
 sky130_fd_sc_hd__and2_2 _23770_ (.A(_19693_),
    .B(_00015_),
    .X(_02754_));
 sky130_fd_sc_hd__and2_2 _23771_ (.A(_19693_),
    .B(_00016_),
    .X(_02753_));
 sky130_fd_sc_hd__and2_2 _23772_ (.A(_19693_),
    .B(_00017_),
    .X(_02752_));
 sky130_fd_sc_hd__and2_2 _23773_ (.A(_19693_),
    .B(_00018_),
    .X(_02751_));
 sky130_fd_sc_hd__and2_2 _23774_ (.A(_19693_),
    .B(_00019_),
    .X(_02750_));
 sky130_fd_sc_hd__and2_2 _23775_ (.A(_19693_),
    .B(_00020_),
    .X(_02749_));
 sky130_fd_sc_hd__buf_1 _23776_ (.A(_18395_),
    .X(_19694_));
 sky130_fd_sc_hd__and2_2 _23777_ (.A(_19694_),
    .B(_00021_),
    .X(_02748_));
 sky130_fd_sc_hd__and2_2 _23778_ (.A(_19694_),
    .B(_00022_),
    .X(_02747_));
 sky130_fd_sc_hd__and2_2 _23779_ (.A(_19694_),
    .B(_00023_),
    .X(_02746_));
 sky130_fd_sc_hd__and2_2 _23780_ (.A(_19694_),
    .B(_00024_),
    .X(_02745_));
 sky130_fd_sc_hd__and2_2 _23781_ (.A(_19694_),
    .B(_00025_),
    .X(_02744_));
 sky130_fd_sc_hd__and2_2 _23782_ (.A(_19694_),
    .B(_00026_),
    .X(_02743_));
 sky130_fd_sc_hd__and2_2 _23783_ (.A(_18396_),
    .B(_00027_),
    .X(_02742_));
 sky130_fd_sc_hd__and2_2 _23784_ (.A(_18396_),
    .B(_00028_),
    .X(_02741_));
 sky130_fd_sc_hd__and2_2 _23785_ (.A(_18396_),
    .B(_00029_),
    .X(_02740_));
 sky130_fd_sc_hd__and2_2 _23786_ (.A(_18396_),
    .B(_00030_),
    .X(_02739_));
 sky130_fd_sc_hd__nand2_2 _23787_ (.A(_19436_),
    .B(\mem_rdata_q[21] ),
    .Y(_19695_));
 sky130_fd_sc_hd__buf_1 _23788_ (.A(_18262_),
    .X(_19696_));
 sky130_fd_sc_hd__nand2_2 _23789_ (.A(\decoded_imm_uj[1] ),
    .B(_19696_),
    .Y(_19697_));
 sky130_fd_sc_hd__nor2_2 _23790_ (.A(is_beq_bne_blt_bge_bltu_bgeu),
    .B(is_sb_sh_sw),
    .Y(_19698_));
 sky130_fd_sc_hd__inv_2 _23791_ (.A(_19698_),
    .Y(_19699_));
 sky130_fd_sc_hd__nand2_2 _23792_ (.A(_19699_),
    .B(\mem_rdata_q[8] ),
    .Y(_19700_));
 sky130_fd_sc_hd__a31o_2 _23793_ (.A1(_19695_),
    .A2(_19697_),
    .A3(_19700_),
    .B1(_18427_),
    .X(_19701_));
 sky130_fd_sc_hd__a21bo_2 _23794_ (.A1(\decoded_imm[1] ),
    .A2(_19475_),
    .B1_N(_19701_),
    .X(_02738_));
 sky130_fd_sc_hd__inv_2 _23795_ (.A(\decoded_imm[2] ),
    .Y(_19702_));
 sky130_fd_sc_hd__nand2_2 _23796_ (.A(_19436_),
    .B(\mem_rdata_q[22] ),
    .Y(_19703_));
 sky130_fd_sc_hd__nand2_2 _23797_ (.A(\decoded_imm_uj[2] ),
    .B(_18263_),
    .Y(_19704_));
 sky130_fd_sc_hd__nand2_2 _23798_ (.A(_19699_),
    .B(\mem_rdata_q[9] ),
    .Y(_19705_));
 sky130_fd_sc_hd__buf_1 _23799_ (.A(_18391_),
    .X(_19706_));
 sky130_fd_sc_hd__a31o_2 _23800_ (.A1(_19703_),
    .A2(_19704_),
    .A3(_19705_),
    .B1(_19706_),
    .X(_19707_));
 sky130_fd_sc_hd__o21ai_2 _23801_ (.A1(_19702_),
    .A2(_19419_),
    .B1(_19707_),
    .Y(_02737_));
 sky130_fd_sc_hd__inv_2 _23802_ (.A(\decoded_imm[3] ),
    .Y(_19708_));
 sky130_fd_sc_hd__nand2_2 _23803_ (.A(_19436_),
    .B(\mem_rdata_q[23] ),
    .Y(_19709_));
 sky130_fd_sc_hd__nand2_2 _23804_ (.A(\decoded_imm_uj[3] ),
    .B(_18263_),
    .Y(_19710_));
 sky130_fd_sc_hd__nand2_2 _23805_ (.A(_19699_),
    .B(\mem_rdata_q[10] ),
    .Y(_19711_));
 sky130_fd_sc_hd__a31o_2 _23806_ (.A1(_19709_),
    .A2(_19710_),
    .A3(_19711_),
    .B1(_19706_),
    .X(_19712_));
 sky130_fd_sc_hd__o21ai_2 _23807_ (.A1(_19708_),
    .A2(_19419_),
    .B1(_19712_),
    .Y(_02736_));
 sky130_fd_sc_hd__inv_2 _23808_ (.A(\decoded_imm[4] ),
    .Y(_19713_));
 sky130_fd_sc_hd__nand2_2 _23809_ (.A(_19436_),
    .B(_19455_),
    .Y(_19714_));
 sky130_fd_sc_hd__nand2_2 _23810_ (.A(\decoded_imm_uj[4] ),
    .B(_18263_),
    .Y(_19715_));
 sky130_fd_sc_hd__nand2_2 _23811_ (.A(_19699_),
    .B(\mem_rdata_q[11] ),
    .Y(_19716_));
 sky130_fd_sc_hd__a31o_2 _23812_ (.A1(_19714_),
    .A2(_19715_),
    .A3(_19716_),
    .B1(_19706_),
    .X(_19717_));
 sky130_fd_sc_hd__o21ai_2 _23813_ (.A1(_19713_),
    .A2(_19419_),
    .B1(_19717_),
    .Y(_02735_));
 sky130_fd_sc_hd__nor2_2 _23814_ (.A(_19699_),
    .B(_19435_),
    .Y(_19718_));
 sky130_fd_sc_hd__inv_2 _23815_ (.A(_19718_),
    .Y(_19719_));
 sky130_fd_sc_hd__a22o_2 _23816_ (.A1(\decoded_imm_uj[5] ),
    .A2(_18263_),
    .B1(_19719_),
    .B2(_19445_),
    .X(_19720_));
 sky130_fd_sc_hd__mux2_2 _23817_ (.A0(_19720_),
    .A1(\decoded_imm[5] ),
    .S(_18386_),
    .X(_02734_));
 sky130_fd_sc_hd__buf_1 _23818_ (.A(instr_jal),
    .X(_19721_));
 sky130_fd_sc_hd__a22o_2 _23819_ (.A1(\decoded_imm_uj[6] ),
    .A2(_19721_),
    .B1(_19719_),
    .B2(_19452_),
    .X(_19722_));
 sky130_fd_sc_hd__buf_1 _23820_ (.A(_18391_),
    .X(_19723_));
 sky130_fd_sc_hd__mux2_2 _23821_ (.A0(_19722_),
    .A1(\decoded_imm[6] ),
    .S(_19723_),
    .X(_02733_));
 sky130_fd_sc_hd__a22o_2 _23822_ (.A1(\decoded_imm_uj[7] ),
    .A2(_19721_),
    .B1(_19719_),
    .B2(\mem_rdata_q[27] ),
    .X(_19724_));
 sky130_fd_sc_hd__mux2_2 _23823_ (.A0(_19724_),
    .A1(\decoded_imm[7] ),
    .S(_19723_),
    .X(_02732_));
 sky130_fd_sc_hd__a22o_2 _23824_ (.A1(\decoded_imm_uj[8] ),
    .A2(_19721_),
    .B1(_19719_),
    .B2(\mem_rdata_q[28] ),
    .X(_19725_));
 sky130_fd_sc_hd__mux2_2 _23825_ (.A0(_19725_),
    .A1(\decoded_imm[8] ),
    .S(_19723_),
    .X(_02731_));
 sky130_fd_sc_hd__a22o_2 _23826_ (.A1(\decoded_imm_uj[9] ),
    .A2(_19721_),
    .B1(_19719_),
    .B2(\mem_rdata_q[29] ),
    .X(_19726_));
 sky130_fd_sc_hd__mux2_2 _23827_ (.A0(_19726_),
    .A1(\decoded_imm[9] ),
    .S(_19723_),
    .X(_02730_));
 sky130_fd_sc_hd__a22o_2 _23828_ (.A1(\decoded_imm_uj[10] ),
    .A2(_19721_),
    .B1(_19719_),
    .B2(\mem_rdata_q[30] ),
    .X(_19727_));
 sky130_fd_sc_hd__mux2_2 _23829_ (.A0(_19727_),
    .A1(\decoded_imm[10] ),
    .S(_19723_),
    .X(_02729_));
 sky130_fd_sc_hd__o21a_2 _23830_ (.A1(_19415_),
    .A2(_19435_),
    .B1(_19493_),
    .X(_19728_));
 sky130_fd_sc_hd__a221o_2 _23831_ (.A1(_18338_),
    .A2(\mem_rdata_q[7] ),
    .B1(\decoded_imm_uj[11] ),
    .B2(_18262_),
    .C1(_19728_),
    .X(_19729_));
 sky130_fd_sc_hd__mux2_2 _23832_ (.A0(_19729_),
    .A1(\decoded_imm[11] ),
    .S(_19723_),
    .X(_02728_));
 sky130_fd_sc_hd__inv_2 _23833_ (.A(_18218_),
    .Y(_19730_));
 sky130_fd_sc_hd__buf_1 _23834_ (.A(_19730_),
    .X(_19731_));
 sky130_fd_sc_hd__nor2_2 _23835_ (.A(_18363_),
    .B(_19718_),
    .Y(_19732_));
 sky130_fd_sc_hd__buf_1 _23836_ (.A(_19732_),
    .X(_19733_));
 sky130_fd_sc_hd__a221o_2 _23837_ (.A1(\decoded_imm_uj[12] ),
    .A2(_19696_),
    .B1(_18398_),
    .B2(_19731_),
    .C1(_19733_),
    .X(_19734_));
 sky130_fd_sc_hd__buf_1 _23838_ (.A(_18391_),
    .X(_19735_));
 sky130_fd_sc_hd__mux2_2 _23839_ (.A0(_19734_),
    .A1(\decoded_imm[12] ),
    .S(_19735_),
    .X(_02727_));
 sky130_fd_sc_hd__a221o_2 _23840_ (.A1(\decoded_imm_uj[13] ),
    .A2(_19696_),
    .B1(\mem_rdata_q[13] ),
    .B2(_19731_),
    .C1(_19733_),
    .X(_19736_));
 sky130_fd_sc_hd__mux2_2 _23841_ (.A0(_19736_),
    .A1(\decoded_imm[13] ),
    .S(_19735_),
    .X(_02726_));
 sky130_fd_sc_hd__buf_1 _23842_ (.A(_19730_),
    .X(_19737_));
 sky130_fd_sc_hd__a221o_2 _23843_ (.A1(\decoded_imm_uj[14] ),
    .A2(_19696_),
    .B1(_18379_),
    .B2(_19737_),
    .C1(_19733_),
    .X(_19738_));
 sky130_fd_sc_hd__mux2_2 _23844_ (.A0(_19738_),
    .A1(\decoded_imm[14] ),
    .S(_19735_),
    .X(_02725_));
 sky130_fd_sc_hd__a221o_2 _23845_ (.A1(\decoded_imm_uj[15] ),
    .A2(_19696_),
    .B1(\mem_rdata_q[15] ),
    .B2(_19737_),
    .C1(_19733_),
    .X(_19739_));
 sky130_fd_sc_hd__mux2_2 _23846_ (.A0(_19739_),
    .A1(\decoded_imm[15] ),
    .S(_19735_),
    .X(_02724_));
 sky130_fd_sc_hd__a221o_2 _23847_ (.A1(\decoded_imm_uj[16] ),
    .A2(_19696_),
    .B1(\mem_rdata_q[16] ),
    .B2(_19737_),
    .C1(_19733_),
    .X(_19740_));
 sky130_fd_sc_hd__mux2_2 _23848_ (.A0(_19740_),
    .A1(\decoded_imm[16] ),
    .S(_19735_),
    .X(_02723_));
 sky130_fd_sc_hd__a221o_2 _23849_ (.A1(\decoded_imm_uj[17] ),
    .A2(_18262_),
    .B1(\mem_rdata_q[17] ),
    .B2(_19737_),
    .C1(_19733_),
    .X(_19741_));
 sky130_fd_sc_hd__mux2_2 _23850_ (.A0(_19741_),
    .A1(\decoded_imm[17] ),
    .S(_19735_),
    .X(_02722_));
 sky130_fd_sc_hd__a221o_2 _23851_ (.A1(\decoded_imm_uj[18] ),
    .A2(_18262_),
    .B1(\mem_rdata_q[18] ),
    .B2(_19737_),
    .C1(_19732_),
    .X(_19742_));
 sky130_fd_sc_hd__mux2_2 _23852_ (.A0(_19742_),
    .A1(\decoded_imm[18] ),
    .S(_19706_),
    .X(_02721_));
 sky130_fd_sc_hd__a221o_2 _23853_ (.A1(\decoded_imm_uj[19] ),
    .A2(_18262_),
    .B1(\mem_rdata_q[19] ),
    .B2(_19737_),
    .C1(_19732_),
    .X(_19743_));
 sky130_fd_sc_hd__mux2_2 _23854_ (.A0(_19743_),
    .A1(\decoded_imm[19] ),
    .S(_19706_),
    .X(_02720_));
 sky130_fd_sc_hd__buf_1 _23855_ (.A(_18218_),
    .X(_19744_));
 sky130_fd_sc_hd__o21ai_2 _23856_ (.A1(_19466_),
    .A2(_19744_),
    .B1(_19499_),
    .Y(_19745_));
 sky130_fd_sc_hd__a22o_2 _23857_ (.A1(_19425_),
    .A2(instr_jal),
    .B1(_19699_),
    .B2(_19493_),
    .X(_19746_));
 sky130_fd_sc_hd__buf_1 _23858_ (.A(_19746_),
    .X(_19747_));
 sky130_fd_sc_hd__and2_2 _23859_ (.A(_19436_),
    .B(_19493_),
    .X(_19748_));
 sky130_fd_sc_hd__buf_1 _23860_ (.A(_19748_),
    .X(_19749_));
 sky130_fd_sc_hd__o32a_2 _23861_ (.A1(_19745_),
    .A2(_19747_),
    .A3(_19749_),
    .B1(\decoded_imm[20] ),
    .B2(_19419_),
    .X(_02719_));
 sky130_fd_sc_hd__buf_1 _23862_ (.A(_19447_),
    .X(_19750_));
 sky130_fd_sc_hd__o21ai_2 _23863_ (.A1(_19479_),
    .A2(_19744_),
    .B1(_19750_),
    .Y(_19751_));
 sky130_fd_sc_hd__o32a_2 _23864_ (.A1(_19751_),
    .A2(_19747_),
    .A3(_19749_),
    .B1(\decoded_imm[21] ),
    .B2(_19419_),
    .X(_02718_));
 sky130_fd_sc_hd__a21o_2 _23865_ (.A1(\mem_rdata_q[22] ),
    .A2(_19731_),
    .B1(_18385_),
    .X(_19752_));
 sky130_fd_sc_hd__buf_1 _23866_ (.A(_18353_),
    .X(_19753_));
 sky130_fd_sc_hd__o32a_2 _23867_ (.A1(_19747_),
    .A2(_19748_),
    .A3(_19752_),
    .B1(\decoded_imm[22] ),
    .B2(_19753_),
    .X(_02717_));
 sky130_fd_sc_hd__a21o_2 _23868_ (.A1(\mem_rdata_q[23] ),
    .A2(_19731_),
    .B1(_18385_),
    .X(_19754_));
 sky130_fd_sc_hd__o32a_2 _23869_ (.A1(_19747_),
    .A2(_19748_),
    .A3(_19754_),
    .B1(\decoded_imm[23] ),
    .B2(_19753_),
    .X(_02716_));
 sky130_fd_sc_hd__a21o_2 _23870_ (.A1(_19455_),
    .A2(_19731_),
    .B1(_18385_),
    .X(_19755_));
 sky130_fd_sc_hd__o32a_2 _23871_ (.A1(_19747_),
    .A2(_19748_),
    .A3(_19755_),
    .B1(\decoded_imm[24] ),
    .B2(_19753_),
    .X(_02715_));
 sky130_fd_sc_hd__o21ai_2 _23872_ (.A1(_18361_),
    .A2(_19744_),
    .B1(_19750_),
    .Y(_19756_));
 sky130_fd_sc_hd__o32a_2 _23873_ (.A1(_19756_),
    .A2(_19746_),
    .A3(_19749_),
    .B1(\decoded_imm[25] ),
    .B2(_19753_),
    .X(_02714_));
 sky130_fd_sc_hd__a21o_2 _23874_ (.A1(_19452_),
    .A2(_19731_),
    .B1(_18385_),
    .X(_19757_));
 sky130_fd_sc_hd__o32a_2 _23875_ (.A1(_19747_),
    .A2(_19748_),
    .A3(_19757_),
    .B1(\decoded_imm[26] ),
    .B2(_19753_),
    .X(_02713_));
 sky130_fd_sc_hd__o21ai_2 _23876_ (.A1(_18360_),
    .A2(_19744_),
    .B1(_19750_),
    .Y(_19758_));
 sky130_fd_sc_hd__o32a_2 _23877_ (.A1(_19758_),
    .A2(_19746_),
    .A3(_19749_),
    .B1(\decoded_imm[27] ),
    .B2(_19753_),
    .X(_02712_));
 sky130_fd_sc_hd__o21ai_2 _23878_ (.A1(_19451_),
    .A2(_19744_),
    .B1(_19750_),
    .Y(_19759_));
 sky130_fd_sc_hd__o32a_2 _23879_ (.A1(_19759_),
    .A2(_19746_),
    .A3(_19749_),
    .B1(\decoded_imm[28] ),
    .B2(_19495_),
    .X(_02711_));
 sky130_fd_sc_hd__o21ai_2 _23880_ (.A1(_18365_),
    .A2(_19744_),
    .B1(_19750_),
    .Y(_19760_));
 sky130_fd_sc_hd__o32a_2 _23881_ (.A1(_19760_),
    .A2(_19746_),
    .A3(_19749_),
    .B1(\decoded_imm[29] ),
    .B2(_19495_),
    .X(_02710_));
 sky130_fd_sc_hd__o21ai_2 _23882_ (.A1(_18364_),
    .A2(_18218_),
    .B1(_19750_),
    .Y(_19761_));
 sky130_fd_sc_hd__o32a_2 _23883_ (.A1(_19761_),
    .A2(_19746_),
    .A3(_19748_),
    .B1(\decoded_imm[30] ),
    .B2(_19495_),
    .X(_02709_));
 sky130_fd_sc_hd__nand2_2 _23884_ (.A(_19718_),
    .B(_18218_),
    .Y(_19762_));
 sky130_fd_sc_hd__a22o_2 _23885_ (.A1(_19426_),
    .A2(_19721_),
    .B1(_19762_),
    .B2(_19493_),
    .X(_19763_));
 sky130_fd_sc_hd__mux2_2 _23886_ (.A0(_19763_),
    .A1(\decoded_imm[31] ),
    .S(_19706_),
    .X(_02708_));
 sky130_fd_sc_hd__and2_2 _23887_ (.A(_18202_),
    .B(_20582_),
    .X(_19764_));
 sky130_fd_sc_hd__or4b_2 _23888_ (.A(_18017_),
    .B(_18250_),
    .C(_00331_),
    .D_N(_19189_),
    .X(_19765_));
 sky130_fd_sc_hd__buf_1 _23889_ (.A(_19765_),
    .X(_19766_));
 sky130_fd_sc_hd__mux2_2 _23890_ (.A0(_19764_),
    .A1(\latched_rd[0] ),
    .S(_19766_),
    .X(_02707_));
 sky130_fd_sc_hd__nor2_2 _23891_ (.A(_02542_),
    .B(_00308_),
    .Y(_19767_));
 sky130_fd_sc_hd__and2b_2 _23892_ (.A_N(_19766_),
    .B(\decoded_rd[1] ),
    .X(_19768_));
 sky130_fd_sc_hd__a22o_2 _23893_ (.A1(\latched_rd[1] ),
    .A2(_19766_),
    .B1(_19767_),
    .B2(_19768_),
    .X(_02706_));
 sky130_fd_sc_hd__and2b_2 _23894_ (.A_N(_19766_),
    .B(\decoded_rd[2] ),
    .X(_19769_));
 sky130_fd_sc_hd__a22o_2 _23895_ (.A1(\latched_rd[2] ),
    .A2(_19766_),
    .B1(_19767_),
    .B2(_19769_),
    .X(_02705_));
 sky130_fd_sc_hd__and2b_2 _23896_ (.A_N(_19765_),
    .B(\decoded_rd[3] ),
    .X(_19770_));
 sky130_fd_sc_hd__a22o_2 _23897_ (.A1(\latched_rd[3] ),
    .A2(_19766_),
    .B1(_19767_),
    .B2(_19770_),
    .X(_02704_));
 sky130_fd_sc_hd__buf_1 _23898_ (.A(_18193_),
    .X(_19771_));
 sky130_fd_sc_hd__nor2_2 _23899_ (.A(is_jalr_addi_slti_sltiu_xori_ori_andi),
    .B(is_slli_srli_srai),
    .Y(_01304_));
 sky130_fd_sc_hd__inv_2 _23900_ (.A(is_lui_auipc_jal),
    .Y(_19772_));
 sky130_fd_sc_hd__and2_2 _23901_ (.A(_01304_),
    .B(_19772_),
    .X(_19773_));
 sky130_fd_sc_hd__o32a_2 _23902_ (.A1(_19415_),
    .A2(_18227_),
    .A3(_00310_),
    .B1(_19771_),
    .B2(_19773_),
    .X(_19774_));
 sky130_fd_sc_hd__inv_2 _23903_ (.A(_19774_),
    .Y(_19775_));
 sky130_fd_sc_hd__and2_2 _23904_ (.A(_19775_),
    .B(_19133_),
    .X(_02703_));
 sky130_fd_sc_hd__inv_2 _23905_ (.A(mem_la_wdata[4]),
    .Y(_19776_));
 sky130_fd_sc_hd__buf_1 _23906_ (.A(_19776_),
    .X(_19777_));
 sky130_fd_sc_hd__buf_1 _23907_ (.A(_19777_),
    .X(_02327_));
 sky130_fd_sc_hd__and2_2 _23908_ (.A(_02327_),
    .B(_02558_),
    .X(_02702_));
 sky130_fd_sc_hd__and2_2 _23909_ (.A(_02327_),
    .B(_02557_),
    .X(_02701_));
 sky130_fd_sc_hd__and2_2 _23910_ (.A(_02327_),
    .B(_02556_),
    .X(_02700_));
 sky130_fd_sc_hd__and2_2 _23911_ (.A(_02327_),
    .B(_02555_),
    .X(_02699_));
 sky130_fd_sc_hd__and2_2 _23912_ (.A(_19777_),
    .B(_02554_),
    .X(_02698_));
 sky130_fd_sc_hd__and2_2 _23913_ (.A(_19777_),
    .B(_02553_),
    .X(_02697_));
 sky130_fd_sc_hd__and2_2 _23914_ (.A(_19777_),
    .B(_02552_),
    .X(_02696_));
 sky130_fd_sc_hd__and2_2 _23915_ (.A(_19777_),
    .B(_02551_),
    .X(_02695_));
 sky130_fd_sc_hd__buf_1 _23916_ (.A(_19153_),
    .X(_19778_));
 sky130_fd_sc_hd__inv_2 _23917_ (.A(_00122_),
    .Y(_19779_));
 sky130_fd_sc_hd__nor2_2 _23918_ (.A(_19778_),
    .B(_19779_),
    .Y(_02550_));
 sky130_fd_sc_hd__nor2_2 _23919_ (.A(_19152_),
    .B(_19153_),
    .Y(_19780_));
 sky130_fd_sc_hd__inv_2 _23920_ (.A(_19780_),
    .Y(_19781_));
 sky130_fd_sc_hd__nor2_2 _23921_ (.A(_19779_),
    .B(_19781_),
    .Y(_02694_));
 sky130_fd_sc_hd__inv_2 _23922_ (.A(_00116_),
    .Y(_19782_));
 sky130_fd_sc_hd__nor2_2 _23923_ (.A(_19778_),
    .B(_19782_),
    .Y(_02549_));
 sky130_fd_sc_hd__nor2_2 _23924_ (.A(_19782_),
    .B(_19781_),
    .Y(_02693_));
 sky130_fd_sc_hd__inv_2 _23925_ (.A(_00110_),
    .Y(_19783_));
 sky130_fd_sc_hd__nor2_2 _23926_ (.A(_19778_),
    .B(_19783_),
    .Y(_02548_));
 sky130_fd_sc_hd__nor2_2 _23927_ (.A(_19783_),
    .B(_19781_),
    .Y(_02692_));
 sky130_fd_sc_hd__inv_2 _23928_ (.A(_00104_),
    .Y(_19784_));
 sky130_fd_sc_hd__nor2_2 _23929_ (.A(_19778_),
    .B(_19784_),
    .Y(_02547_));
 sky130_fd_sc_hd__nor2_2 _23930_ (.A(_19784_),
    .B(_19781_),
    .Y(_02691_));
 sky130_fd_sc_hd__nor2_2 _23931_ (.A(mem_la_wdata[3]),
    .B(mem_la_wdata[2]),
    .Y(_19785_));
 sky130_fd_sc_hd__and2_2 _23932_ (.A(_19785_),
    .B(_00094_),
    .X(_02546_));
 sky130_fd_sc_hd__inv_2 _23933_ (.A(mem_la_wdata[2]),
    .Y(_19786_));
 sky130_fd_sc_hd__buf_1 _23934_ (.A(_19786_),
    .X(_02321_));
 sky130_fd_sc_hd__and3_2 _23935_ (.A(_19780_),
    .B(_02321_),
    .C(_00094_),
    .X(_02690_));
 sky130_fd_sc_hd__and2_2 _23936_ (.A(_19785_),
    .B(_00084_),
    .X(_02545_));
 sky130_fd_sc_hd__and3_2 _23937_ (.A(_19780_),
    .B(_19786_),
    .C(_00084_),
    .X(_02689_));
 sky130_fd_sc_hd__inv_2 _23938_ (.A(_19155_),
    .Y(_19787_));
 sky130_fd_sc_hd__buf_1 _23939_ (.A(_19787_),
    .X(_02318_));
 sky130_fd_sc_hd__and3_2 _23940_ (.A(_19785_),
    .B(_02318_),
    .C(_00066_),
    .X(_02544_));
 sky130_fd_sc_hd__and2_2 _23941_ (.A(_02318_),
    .B(_00066_),
    .X(_00067_));
 sky130_fd_sc_hd__and3_2 _23942_ (.A(_00067_),
    .B(_19786_),
    .C(_19780_),
    .X(_02688_));
 sky130_fd_sc_hd__nor2_2 _23943_ (.A(mem_la_wdata[1]),
    .B(mem_la_wdata[0]),
    .Y(_19788_));
 sky130_fd_sc_hd__and3_2 _23944_ (.A(_19785_),
    .B(_19788_),
    .C(_19535_),
    .X(_02543_));
 sky130_fd_sc_hd__inv_2 _23945_ (.A(pcpi_rs1[0]),
    .Y(_19789_));
 sky130_fd_sc_hd__buf_1 _23946_ (.A(_19789_),
    .X(_19790_));
 sky130_fd_sc_hd__nand2_2 _23947_ (.A(_19785_),
    .B(_19788_),
    .Y(_19791_));
 sky130_fd_sc_hd__nor2_2 _23948_ (.A(mem_la_wdata[4]),
    .B(_19791_),
    .Y(_19792_));
 sky130_fd_sc_hd__inv_2 _23949_ (.A(_19792_),
    .Y(_19793_));
 sky130_fd_sc_hd__nor2_2 _23950_ (.A(_19790_),
    .B(_19793_),
    .Y(_02687_));
 sky130_fd_sc_hd__o211a_2 _23951_ (.A1(\reg_pc[1] ),
    .A2(\reg_next_pc[0] ),
    .B1(_18024_),
    .C1(mem_do_rinst),
    .X(_00307_));
 sky130_fd_sc_hd__and3_2 _23952_ (.A(_18154_),
    .B(_18331_),
    .C(_18081_),
    .X(_00312_));
 sky130_fd_sc_hd__nor2_2 _23953_ (.A(_18016_),
    .B(_18011_),
    .Y(_00303_));
 sky130_fd_sc_hd__inv_2 _23954_ (.A(_00303_),
    .Y(_19794_));
 sky130_fd_sc_hd__nor2_2 _23955_ (.A(_00307_),
    .B(_19794_),
    .Y(_19795_));
 sky130_fd_sc_hd__inv_2 _23956_ (.A(\mem_wordsize[2] ),
    .Y(_19796_));
 sky130_fd_sc_hd__nor2_2 _23957_ (.A(_19789_),
    .B(_19796_),
    .Y(_00306_));
 sky130_fd_sc_hd__nor2_2 _23958_ (.A(irq_active),
    .B(\irq_mask[2] ),
    .Y(_19797_));
 sky130_fd_sc_hd__nand2_2 _23959_ (.A(_00306_),
    .B(_19797_),
    .Y(_19798_));
 sky130_fd_sc_hd__nor2_2 _23960_ (.A(irq_active),
    .B(\irq_mask[1] ),
    .Y(_19799_));
 sky130_fd_sc_hd__and3_2 _23961_ (.A(_18855_),
    .B(_18163_),
    .C(_19799_),
    .X(_19800_));
 sky130_fd_sc_hd__o211a_2 _23962_ (.A1(_18080_),
    .A2(_00309_),
    .B1(_18451_),
    .C1(_18147_),
    .X(_19801_));
 sky130_fd_sc_hd__a21oi_2 _23963_ (.A1(_18856_),
    .A2(_19800_),
    .B1(_19801_),
    .Y(_19802_));
 sky130_fd_sc_hd__inv_2 _23964_ (.A(\mem_wordsize[0] ),
    .Y(_19803_));
 sky130_fd_sc_hd__nor2_2 _23965_ (.A(_19533_),
    .B(pcpi_rs1[0]),
    .Y(_00304_));
 sky130_fd_sc_hd__nor2_2 _23966_ (.A(_19803_),
    .B(_00304_),
    .Y(_00305_));
 sky130_fd_sc_hd__nor2_2 _23967_ (.A(_00306_),
    .B(_00305_),
    .Y(_19804_));
 sky130_fd_sc_hd__buf_1 _23968_ (.A(_19797_),
    .X(_19805_));
 sky130_fd_sc_hd__o21ai_2 _23969_ (.A1(_19804_),
    .A2(_19805_),
    .B1(_03828_),
    .Y(_19806_));
 sky130_fd_sc_hd__o21ai_2 _23970_ (.A1(_19798_),
    .A2(_19802_),
    .B1(_19806_),
    .Y(_19807_));
 sky130_fd_sc_hd__o21ai_2 _23971_ (.A1(_18011_),
    .A2(_00307_),
    .B1(_03828_),
    .Y(_19808_));
 sky130_fd_sc_hd__nand2_2 _23972_ (.A(_18200_),
    .B(_18250_),
    .Y(_19809_));
 sky130_fd_sc_hd__or2_2 _23973_ (.A(_18011_),
    .B(_19804_),
    .X(_19810_));
 sky130_fd_sc_hd__inv_2 _23974_ (.A(_00307_),
    .Y(_19811_));
 sky130_fd_sc_hd__a21oi_2 _23975_ (.A1(_19810_),
    .A2(_19811_),
    .B1(_19805_),
    .Y(_19812_));
 sky130_fd_sc_hd__a21oi_2 _23976_ (.A1(_19808_),
    .A2(_19809_),
    .B1(_19812_),
    .Y(_19813_));
 sky130_fd_sc_hd__nor2_2 _23977_ (.A(_19794_),
    .B(_19804_),
    .Y(_19814_));
 sky130_fd_sc_hd__nor2_2 _23978_ (.A(_00307_),
    .B(_19814_),
    .Y(_19815_));
 sky130_fd_sc_hd__nor2_2 _23979_ (.A(_19805_),
    .B(_19815_),
    .Y(_19816_));
 sky130_fd_sc_hd__a211o_2 _23980_ (.A1(_18338_),
    .A2(_18014_),
    .B1(_18252_),
    .C1(_19816_),
    .X(_19817_));
 sky130_fd_sc_hd__or4b_2 _23981_ (.A(_18300_),
    .B(_00314_),
    .C(_19813_),
    .D_N(_19817_),
    .X(_19818_));
 sky130_fd_sc_hd__inv_2 _23982_ (.A(_00306_),
    .Y(_19819_));
 sky130_fd_sc_hd__inv_2 _23983_ (.A(_19797_),
    .Y(_19820_));
 sky130_fd_sc_hd__inv_2 _23984_ (.A(_00305_),
    .Y(_19821_));
 sky130_fd_sc_hd__nor2_2 _23985_ (.A(_19820_),
    .B(_19821_),
    .Y(_19822_));
 sky130_fd_sc_hd__nor2_2 _23986_ (.A(_19820_),
    .B(_19811_),
    .Y(_19823_));
 sky130_fd_sc_hd__nor2_2 _23987_ (.A(_19823_),
    .B(_19815_),
    .Y(_19824_));
 sky130_fd_sc_hd__inv_2 _23988_ (.A(_19824_),
    .Y(_19825_));
 sky130_fd_sc_hd__a31o_2 _23989_ (.A1(_19795_),
    .A2(_19819_),
    .A3(_19822_),
    .B1(_19825_),
    .X(_19826_));
 sky130_fd_sc_hd__a2bb2o_2 _23990_ (.A1_N(_18163_),
    .A2_N(_19816_),
    .B1(_19800_),
    .B2(_19826_),
    .X(_19827_));
 sky130_fd_sc_hd__and3_2 _23991_ (.A(_18856_),
    .B(_18637_),
    .C(_19827_),
    .X(_19828_));
 sky130_fd_sc_hd__nor2_2 _23992_ (.A(_19449_),
    .B(_18874_),
    .Y(_19829_));
 sky130_fd_sc_hd__o21a_2 _23993_ (.A1(_00309_),
    .A2(_19829_),
    .B1(_19823_),
    .X(_19830_));
 sky130_fd_sc_hd__o211a_2 _23994_ (.A1(_19821_),
    .A2(_19797_),
    .B1(_19819_),
    .C1(_19795_),
    .X(_19831_));
 sky130_fd_sc_hd__a32o_2 _23995_ (.A1(_18025_),
    .A2(_00308_),
    .A3(_19825_),
    .B1(_18875_),
    .B2(_19831_),
    .X(_19832_));
 sky130_fd_sc_hd__nor2_2 _23996_ (.A(_19798_),
    .B(_19794_),
    .Y(_19833_));
 sky130_fd_sc_hd__or3_2 _23997_ (.A(_00323_),
    .B(_18080_),
    .C(_18151_),
    .X(_19834_));
 sky130_fd_sc_hd__inv_2 _23998_ (.A(_19834_),
    .Y(_02062_));
 sky130_fd_sc_hd__o21a_2 _23999_ (.A1(_19823_),
    .A2(_19833_),
    .B1(_02062_),
    .X(_19835_));
 sky130_fd_sc_hd__a31o_2 _24000_ (.A1(_19822_),
    .A2(_00303_),
    .A3(_19819_),
    .B1(_19810_),
    .X(_19836_));
 sky130_fd_sc_hd__and3_2 _24001_ (.A(_18146_),
    .B(_19797_),
    .C(_19814_),
    .X(_19837_));
 sky130_fd_sc_hd__a31o_2 _24002_ (.A1(_02062_),
    .A2(_18024_),
    .A3(_19836_),
    .B1(_19837_),
    .X(_19838_));
 sky130_fd_sc_hd__a21oi_2 _24003_ (.A1(_18875_),
    .A2(_19794_),
    .B1(_19838_),
    .Y(_19839_));
 sky130_fd_sc_hd__nand2_2 _24004_ (.A(_19819_),
    .B(_19797_),
    .Y(_19840_));
 sky130_fd_sc_hd__a2111o_2 _24005_ (.A1(_19814_),
    .A2(_19840_),
    .B1(decoder_trigger),
    .C1(_00309_),
    .D1(_18874_),
    .X(_19841_));
 sky130_fd_sc_hd__a21oi_2 _24006_ (.A1(_19839_),
    .A2(_19841_),
    .B1(_00307_),
    .Y(_19842_));
 sky130_fd_sc_hd__o41a_2 _24007_ (.A1(_19830_),
    .A2(_19832_),
    .A3(_19835_),
    .A4(_19842_),
    .B1(_18452_),
    .X(_19843_));
 sky130_fd_sc_hd__a2111o_2 _24008_ (.A1(_19795_),
    .A2(_19807_),
    .B1(_19818_),
    .C1(_19828_),
    .D1(_19843_),
    .X(_00039_));
 sky130_fd_sc_hd__nor2_2 _24009_ (.A(_18048_),
    .B(_19816_),
    .Y(_19844_));
 sky130_fd_sc_hd__and2_2 _24010_ (.A(_18265_),
    .B(_19844_),
    .X(_00040_));
 sky130_fd_sc_hd__or2_2 _24011_ (.A(_18851_),
    .B(_18249_),
    .X(_19845_));
 sky130_fd_sc_hd__nand2_2 _24012_ (.A(_18878_),
    .B(_18029_),
    .Y(_19846_));
 sky130_fd_sc_hd__inv_2 _24013_ (.A(_19844_),
    .Y(_19847_));
 sky130_fd_sc_hd__a21oi_2 _24014_ (.A1(_19845_),
    .A2(_19846_),
    .B1(_19847_),
    .Y(_00044_));
 sky130_fd_sc_hd__nand3_2 _24015_ (.A(_18249_),
    .B(_18201_),
    .C(_19773_),
    .Y(_19848_));
 sky130_fd_sc_hd__a21oi_2 _24016_ (.A1(_18858_),
    .A2(_19848_),
    .B1(_19847_),
    .Y(_00041_));
 sky130_fd_sc_hd__and4b_2 _24017_ (.A_N(_19799_),
    .B(_18856_),
    .C(_18163_),
    .D(_18855_),
    .X(_19849_));
 sky130_fd_sc_hd__o31a_2 _24018_ (.A1(\cpu_state[0] ),
    .A2(_19812_),
    .A3(_19849_),
    .B1(_18879_),
    .X(_00038_));
 sky130_fd_sc_hd__nand2_2 _24019_ (.A(_18878_),
    .B(\cpu_state[5] ),
    .Y(_19850_));
 sky130_fd_sc_hd__buf_1 _24020_ (.A(_18257_),
    .X(_19851_));
 sky130_fd_sc_hd__buf_1 _24021_ (.A(_19851_),
    .X(_19852_));
 sky130_fd_sc_hd__nand2_2 _24022_ (.A(_19415_),
    .B(_19852_),
    .Y(_19853_));
 sky130_fd_sc_hd__a21oi_2 _24023_ (.A1(_19850_),
    .A2(_19853_),
    .B1(_19847_),
    .Y(_00043_));
 sky130_fd_sc_hd__o311a_2 _24024_ (.A1(mem_do_rinst),
    .A2(_18015_),
    .A3(mem_do_rdata),
    .B1(_18028_),
    .C1(_00290_),
    .X(mem_la_read));
 sky130_fd_sc_hd__nor2_2 _24025_ (.A(_00291_),
    .B(_19500_),
    .Y(_00317_));
 sky130_fd_sc_hd__o32a_2 _24026_ (.A1(_18191_),
    .A2(_18254_),
    .A3(_19816_),
    .B1(_00302_),
    .B2(_19847_),
    .X(_19854_));
 sky130_fd_sc_hd__a2bb2o_2 _24027_ (.A1_N(_18188_),
    .A2_N(_19854_),
    .B1(_19844_),
    .B2(_19775_),
    .X(_00042_));
 sky130_fd_sc_hd__nor2b_2 _24028_ (.A(pcpi_rs1[0]),
    .B_N(mem_la_wdata[0]),
    .Y(_19855_));
 sky130_fd_sc_hd__nor2_2 _24029_ (.A(mem_la_wdata[0]),
    .B(_19789_),
    .Y(_00048_));
 sky130_fd_sc_hd__nor2_2 _24030_ (.A(_19855_),
    .B(_00048_),
    .Y(_19856_));
 sky130_fd_sc_hd__inv_2 _24031_ (.A(_19856_),
    .Y(_02591_));
 sky130_fd_sc_hd__nor2_2 _24032_ (.A(mem_la_wdata[6]),
    .B(_19528_),
    .Y(_19857_));
 sky130_fd_sc_hd__inv_2 _24033_ (.A(mem_la_wdata[6]),
    .Y(_02333_));
 sky130_fd_sc_hd__inv_2 _24034_ (.A(_19528_),
    .Y(_19858_));
 sky130_fd_sc_hd__nor2_2 _24035_ (.A(_02333_),
    .B(_19858_),
    .Y(_19859_));
 sky130_fd_sc_hd__nor2_2 _24036_ (.A(_19857_),
    .B(_19859_),
    .Y(_19860_));
 sky130_fd_sc_hd__inv_2 _24037_ (.A(_19860_),
    .Y(_19861_));
 sky130_fd_sc_hd__inv_2 _24038_ (.A(mem_la_wdata[7]),
    .Y(_02336_));
 sky130_fd_sc_hd__inv_2 _24039_ (.A(pcpi_rs1[7]),
    .Y(_19862_));
 sky130_fd_sc_hd__nor2_2 _24040_ (.A(_02336_),
    .B(_19862_),
    .Y(_19863_));
 sky130_fd_sc_hd__nand2_2 _24041_ (.A(_02336_),
    .B(_19862_),
    .Y(_19864_));
 sky130_fd_sc_hd__or2b_2 _24042_ (.A(_19863_),
    .B_N(_19864_),
    .X(_19865_));
 sky130_fd_sc_hd__and3_2 _24043_ (.A(_19861_),
    .B(_19856_),
    .C(_19865_),
    .X(_19866_));
 sky130_fd_sc_hd__inv_2 _24044_ (.A(_19534_),
    .Y(_19867_));
 sky130_fd_sc_hd__nor2_2 _24045_ (.A(_19787_),
    .B(_19867_),
    .Y(_19868_));
 sky130_fd_sc_hd__nand2_2 _24046_ (.A(_02318_),
    .B(_19867_),
    .Y(_19869_));
 sky130_fd_sc_hd__or2b_2 _24047_ (.A(_19868_),
    .B_N(_19869_),
    .X(_19870_));
 sky130_fd_sc_hd__nand2_2 _24048_ (.A(_19866_),
    .B(_19870_),
    .Y(_19871_));
 sky130_fd_sc_hd__nor2_2 _24049_ (.A(_19142_),
    .B(_19520_),
    .Y(_19872_));
 sky130_fd_sc_hd__inv_2 _24050_ (.A(pcpi_rs2[15]),
    .Y(_02360_));
 sky130_fd_sc_hd__inv_2 _24051_ (.A(pcpi_rs1[15]),
    .Y(_19873_));
 sky130_fd_sc_hd__nor2_2 _24052_ (.A(_02360_),
    .B(_19873_),
    .Y(_19874_));
 sky130_fd_sc_hd__nor2_2 _24053_ (.A(_19872_),
    .B(_19874_),
    .Y(_19875_));
 sky130_fd_sc_hd__nor2_2 _24054_ (.A(_19145_),
    .B(_19521_),
    .Y(_19876_));
 sky130_fd_sc_hd__inv_2 _24055_ (.A(pcpi_rs2[13]),
    .Y(_02354_));
 sky130_fd_sc_hd__inv_2 _24056_ (.A(pcpi_rs1[13]),
    .Y(_19877_));
 sky130_fd_sc_hd__nor2_2 _24057_ (.A(_02354_),
    .B(_19877_),
    .Y(_19878_));
 sky130_fd_sc_hd__nor2_2 _24058_ (.A(_19876_),
    .B(_19878_),
    .Y(_19879_));
 sky130_fd_sc_hd__nor2_2 _24059_ (.A(pcpi_rs2[12]),
    .B(_19523_),
    .Y(_19880_));
 sky130_fd_sc_hd__inv_2 _24060_ (.A(pcpi_rs2[12]),
    .Y(_02351_));
 sky130_fd_sc_hd__inv_2 _24061_ (.A(pcpi_rs1[12]),
    .Y(_19881_));
 sky130_fd_sc_hd__nor2_2 _24062_ (.A(_02351_),
    .B(_19881_),
    .Y(_19882_));
 sky130_fd_sc_hd__nor2_2 _24063_ (.A(_19880_),
    .B(_19882_),
    .Y(_19883_));
 sky130_fd_sc_hd__nor2_2 _24064_ (.A(_19143_),
    .B(pcpi_rs1[14]),
    .Y(_19884_));
 sky130_fd_sc_hd__inv_2 _24065_ (.A(pcpi_rs2[14]),
    .Y(_02357_));
 sky130_fd_sc_hd__inv_2 _24066_ (.A(pcpi_rs1[14]),
    .Y(_19885_));
 sky130_fd_sc_hd__nor2_2 _24067_ (.A(_02357_),
    .B(_19885_),
    .Y(_19886_));
 sky130_fd_sc_hd__nor2_2 _24068_ (.A(_19884_),
    .B(_19886_),
    .Y(_19887_));
 sky130_fd_sc_hd__or4_2 _24069_ (.A(_19875_),
    .B(_19879_),
    .C(_19883_),
    .D(_19887_),
    .X(_19888_));
 sky130_fd_sc_hd__nor2_2 _24070_ (.A(_19146_),
    .B(_19524_),
    .Y(_19889_));
 sky130_fd_sc_hd__inv_2 _24071_ (.A(pcpi_rs2[11]),
    .Y(_02348_));
 sky130_fd_sc_hd__inv_2 _24072_ (.A(pcpi_rs1[11]),
    .Y(_19890_));
 sky130_fd_sc_hd__nor2_2 _24073_ (.A(_02348_),
    .B(_19890_),
    .Y(_19891_));
 sky130_fd_sc_hd__nor2_2 _24074_ (.A(_19889_),
    .B(_19891_),
    .Y(_19892_));
 sky130_fd_sc_hd__nor2_2 _24075_ (.A(_19147_),
    .B(_19525_),
    .Y(_19893_));
 sky130_fd_sc_hd__inv_2 _24076_ (.A(pcpi_rs2[9]),
    .Y(_02342_));
 sky130_fd_sc_hd__inv_2 _24077_ (.A(pcpi_rs1[9]),
    .Y(_19894_));
 sky130_fd_sc_hd__nor2_2 _24078_ (.A(_02342_),
    .B(_19894_),
    .Y(_19895_));
 sky130_fd_sc_hd__nor2_2 _24079_ (.A(_19893_),
    .B(_19895_),
    .Y(_19896_));
 sky130_fd_sc_hd__nor2_2 _24080_ (.A(pcpi_rs2[8]),
    .B(_19526_),
    .Y(_19897_));
 sky130_fd_sc_hd__inv_2 _24081_ (.A(pcpi_rs2[8]),
    .Y(_02339_));
 sky130_fd_sc_hd__inv_2 _24082_ (.A(pcpi_rs1[8]),
    .Y(_19898_));
 sky130_fd_sc_hd__nor2_2 _24083_ (.A(_02339_),
    .B(_19898_),
    .Y(_19899_));
 sky130_fd_sc_hd__nor2_2 _24084_ (.A(_19897_),
    .B(_19899_),
    .Y(_19900_));
 sky130_fd_sc_hd__nor2_2 _24085_ (.A(pcpi_rs2[10]),
    .B(pcpi_rs1[10]),
    .Y(_19901_));
 sky130_fd_sc_hd__inv_2 _24086_ (.A(pcpi_rs2[10]),
    .Y(_02345_));
 sky130_fd_sc_hd__inv_2 _24087_ (.A(pcpi_rs1[10]),
    .Y(_19902_));
 sky130_fd_sc_hd__nor2_2 _24088_ (.A(_02345_),
    .B(_19902_),
    .Y(_19903_));
 sky130_fd_sc_hd__nor2_2 _24089_ (.A(_19901_),
    .B(_19903_),
    .Y(_19904_));
 sky130_fd_sc_hd__or4_2 _24090_ (.A(_19892_),
    .B(_19896_),
    .C(_19900_),
    .D(_19904_),
    .X(_19905_));
 sky130_fd_sc_hd__nor2_2 _24091_ (.A(mem_la_wdata[4]),
    .B(_19530_),
    .Y(_19906_));
 sky130_fd_sc_hd__inv_2 _24092_ (.A(pcpi_rs1[4]),
    .Y(_19907_));
 sky130_fd_sc_hd__nor2_2 _24093_ (.A(_19776_),
    .B(_19907_),
    .Y(_19908_));
 sky130_fd_sc_hd__nor2_2 _24094_ (.A(_19906_),
    .B(_19908_),
    .Y(_19909_));
 sky130_fd_sc_hd__nor2_2 _24095_ (.A(mem_la_wdata[3]),
    .B(_19531_),
    .Y(_19910_));
 sky130_fd_sc_hd__inv_2 _24096_ (.A(mem_la_wdata[3]),
    .Y(_02324_));
 sky130_fd_sc_hd__inv_2 _24097_ (.A(pcpi_rs1[3]),
    .Y(_19911_));
 sky130_fd_sc_hd__nor2_2 _24098_ (.A(_02324_),
    .B(_19911_),
    .Y(_19912_));
 sky130_fd_sc_hd__nor2_2 _24099_ (.A(_19910_),
    .B(_19912_),
    .Y(_19913_));
 sky130_fd_sc_hd__nor2_2 _24100_ (.A(mem_la_wdata[2]),
    .B(_19532_),
    .Y(_19914_));
 sky130_fd_sc_hd__inv_2 _24101_ (.A(pcpi_rs1[2]),
    .Y(_19915_));
 sky130_fd_sc_hd__nor2_2 _24102_ (.A(_19786_),
    .B(_19915_),
    .Y(_19916_));
 sky130_fd_sc_hd__nor2_2 _24103_ (.A(_19914_),
    .B(_19916_),
    .Y(_19917_));
 sky130_fd_sc_hd__inv_2 _24104_ (.A(mem_la_wdata[5]),
    .Y(_02330_));
 sky130_fd_sc_hd__inv_2 _24105_ (.A(pcpi_rs1[5]),
    .Y(_19918_));
 sky130_fd_sc_hd__nand2_2 _24106_ (.A(_02330_),
    .B(_19918_),
    .Y(_19919_));
 sky130_fd_sc_hd__nand2_2 _24107_ (.A(mem_la_wdata[5]),
    .B(_19529_),
    .Y(_19920_));
 sky130_fd_sc_hd__nand2_2 _24108_ (.A(_19919_),
    .B(_19920_),
    .Y(_19921_));
 sky130_fd_sc_hd__inv_2 _24109_ (.A(_19921_),
    .Y(_19922_));
 sky130_fd_sc_hd__or4_2 _24110_ (.A(_19909_),
    .B(_19913_),
    .C(_19917_),
    .D(_19922_),
    .X(_19923_));
 sky130_fd_sc_hd__or4_2 _24111_ (.A(_19871_),
    .B(_19888_),
    .C(_19905_),
    .D(_19923_),
    .X(_19924_));
 sky130_fd_sc_hd__nor2_2 _24112_ (.A(_19139_),
    .B(_19514_),
    .Y(_19925_));
 sky130_fd_sc_hd__inv_2 _24113_ (.A(_19139_),
    .Y(_02378_));
 sky130_fd_sc_hd__inv_2 _24114_ (.A(pcpi_rs1[21]),
    .Y(_19926_));
 sky130_fd_sc_hd__nor2_2 _24115_ (.A(_02378_),
    .B(_19926_),
    .Y(_19927_));
 sky130_fd_sc_hd__nor2_2 _24116_ (.A(_19925_),
    .B(_19927_),
    .Y(_19928_));
 sky130_fd_sc_hd__nor2_2 _24117_ (.A(_19138_),
    .B(_19512_),
    .Y(_19929_));
 sky130_fd_sc_hd__inv_2 _24118_ (.A(pcpi_rs2[23]),
    .Y(_02384_));
 sky130_fd_sc_hd__inv_2 _24119_ (.A(pcpi_rs1[23]),
    .Y(_19930_));
 sky130_fd_sc_hd__nor2_2 _24120_ (.A(_02384_),
    .B(_19930_),
    .Y(_19931_));
 sky130_fd_sc_hd__nor2_2 _24121_ (.A(_19929_),
    .B(_19931_),
    .Y(_19932_));
 sky130_fd_sc_hd__nor2_2 _24122_ (.A(_19928_),
    .B(_19932_),
    .Y(_19933_));
 sky130_fd_sc_hd__nor2_2 _24123_ (.A(pcpi_rs2[22]),
    .B(_19513_),
    .Y(_19934_));
 sky130_fd_sc_hd__inv_2 _24124_ (.A(pcpi_rs2[22]),
    .Y(_02381_));
 sky130_fd_sc_hd__inv_2 _24125_ (.A(pcpi_rs1[22]),
    .Y(_19935_));
 sky130_fd_sc_hd__nor2_2 _24126_ (.A(_02381_),
    .B(_19935_),
    .Y(_19936_));
 sky130_fd_sc_hd__nor2_2 _24127_ (.A(_19934_),
    .B(_19936_),
    .Y(_19937_));
 sky130_fd_sc_hd__inv_2 _24128_ (.A(_19937_),
    .Y(_19938_));
 sky130_fd_sc_hd__inv_2 _24129_ (.A(pcpi_rs2[20]),
    .Y(_02375_));
 sky130_fd_sc_hd__inv_2 _24130_ (.A(pcpi_rs1[20]),
    .Y(_19939_));
 sky130_fd_sc_hd__nor2_2 _24131_ (.A(_02375_),
    .B(_19939_),
    .Y(_19940_));
 sky130_fd_sc_hd__nand2_2 _24132_ (.A(_02375_),
    .B(_19939_),
    .Y(_19941_));
 sky130_fd_sc_hd__or2b_2 _24133_ (.A(_19940_),
    .B_N(_19941_),
    .X(_19942_));
 sky130_fd_sc_hd__and3_2 _24134_ (.A(_19933_),
    .B(_19938_),
    .C(_19942_),
    .X(_19943_));
 sky130_fd_sc_hd__nor2_2 _24135_ (.A(_19137_),
    .B(_19509_),
    .Y(_19944_));
 sky130_fd_sc_hd__inv_2 _24136_ (.A(pcpi_rs2[25]),
    .Y(_02390_));
 sky130_fd_sc_hd__inv_2 _24137_ (.A(pcpi_rs1[25]),
    .Y(_19945_));
 sky130_fd_sc_hd__nor2_2 _24138_ (.A(_02390_),
    .B(_19945_),
    .Y(_19946_));
 sky130_fd_sc_hd__nor2_2 _24139_ (.A(_19944_),
    .B(_19946_),
    .Y(_19947_));
 sky130_fd_sc_hd__nor2_2 _24140_ (.A(pcpi_rs2[28]),
    .B(_19507_),
    .Y(_19948_));
 sky130_fd_sc_hd__inv_2 _24141_ (.A(pcpi_rs2[28]),
    .Y(_02399_));
 sky130_fd_sc_hd__inv_2 _24142_ (.A(pcpi_rs1[28]),
    .Y(_19949_));
 sky130_fd_sc_hd__nor2_2 _24143_ (.A(_02399_),
    .B(_19949_),
    .Y(_19950_));
 sky130_fd_sc_hd__nor2_2 _24144_ (.A(_19948_),
    .B(_19950_),
    .Y(_19951_));
 sky130_fd_sc_hd__inv_2 _24145_ (.A(pcpi_rs2[26]),
    .Y(_02393_));
 sky130_fd_sc_hd__inv_2 _24146_ (.A(pcpi_rs1[26]),
    .Y(_19952_));
 sky130_fd_sc_hd__nand2_2 _24147_ (.A(_02393_),
    .B(_19952_),
    .Y(_19953_));
 sky130_fd_sc_hd__nand2_2 _24148_ (.A(pcpi_rs2[26]),
    .B(pcpi_rs1[26]),
    .Y(_19954_));
 sky130_fd_sc_hd__nand2_2 _24149_ (.A(_19953_),
    .B(_19954_),
    .Y(_19955_));
 sky130_fd_sc_hd__inv_2 _24150_ (.A(_19955_),
    .Y(_19956_));
 sky130_fd_sc_hd__inv_2 _24151_ (.A(pcpi_rs2[24]),
    .Y(_02387_));
 sky130_fd_sc_hd__inv_2 _24152_ (.A(pcpi_rs1[24]),
    .Y(_19957_));
 sky130_fd_sc_hd__nor2_2 _24153_ (.A(_02387_),
    .B(_19957_),
    .Y(_19958_));
 sky130_fd_sc_hd__nand2_2 _24154_ (.A(_02387_),
    .B(_19957_),
    .Y(_19959_));
 sky130_fd_sc_hd__or2b_2 _24155_ (.A(_19958_),
    .B_N(_19959_),
    .X(_19960_));
 sky130_fd_sc_hd__or4b_2 _24156_ (.A(_19947_),
    .B(_19951_),
    .C(_19956_),
    .D_N(_19960_),
    .X(_19961_));
 sky130_fd_sc_hd__nor2_2 _24157_ (.A(_19134_),
    .B(pcpi_rs1[29]),
    .Y(_19962_));
 sky130_fd_sc_hd__inv_2 _24158_ (.A(pcpi_rs2[29]),
    .Y(_02402_));
 sky130_fd_sc_hd__inv_2 _24159_ (.A(pcpi_rs1[29]),
    .Y(_19963_));
 sky130_fd_sc_hd__nor2_2 _24160_ (.A(_02402_),
    .B(_19963_),
    .Y(_19964_));
 sky130_fd_sc_hd__nor2_2 _24161_ (.A(_19962_),
    .B(_19964_),
    .Y(_19965_));
 sky130_fd_sc_hd__nor2_2 _24162_ (.A(_19135_),
    .B(pcpi_rs1[27]),
    .Y(_19966_));
 sky130_fd_sc_hd__inv_2 _24163_ (.A(pcpi_rs2[27]),
    .Y(_02396_));
 sky130_fd_sc_hd__inv_2 _24164_ (.A(pcpi_rs1[27]),
    .Y(_19967_));
 sky130_fd_sc_hd__nor2_2 _24165_ (.A(_02396_),
    .B(_19967_),
    .Y(_19968_));
 sky130_fd_sc_hd__nor2_2 _24166_ (.A(_19966_),
    .B(_19968_),
    .Y(_19969_));
 sky130_fd_sc_hd__nor2_2 _24167_ (.A(pcpi_rs1[31]),
    .B(pcpi_rs2[31]),
    .Y(_19970_));
 sky130_fd_sc_hd__inv_2 _24168_ (.A(pcpi_rs2[31]),
    .Y(_19971_));
 sky130_fd_sc_hd__nor2_2 _24169_ (.A(_18173_),
    .B(_19971_),
    .Y(_19972_));
 sky130_fd_sc_hd__nor2_2 _24170_ (.A(_19970_),
    .B(_19972_),
    .Y(_19973_));
 sky130_fd_sc_hd__nor2_2 _24171_ (.A(pcpi_rs2[30]),
    .B(pcpi_rs1[30]),
    .Y(_19974_));
 sky130_fd_sc_hd__inv_2 _24172_ (.A(pcpi_rs2[30]),
    .Y(_02405_));
 sky130_fd_sc_hd__inv_2 _24173_ (.A(pcpi_rs1[30]),
    .Y(_19975_));
 sky130_fd_sc_hd__nor2_2 _24174_ (.A(_02405_),
    .B(_19975_),
    .Y(_19976_));
 sky130_fd_sc_hd__nor2_2 _24175_ (.A(_19974_),
    .B(_19976_),
    .Y(_19977_));
 sky130_fd_sc_hd__nor2_2 _24176_ (.A(_19973_),
    .B(_19977_),
    .Y(_19978_));
 sky130_fd_sc_hd__inv_2 _24177_ (.A(_19978_),
    .Y(_19979_));
 sky130_fd_sc_hd__or3_2 _24178_ (.A(_19965_),
    .B(_19969_),
    .C(_19979_),
    .X(_19980_));
 sky130_fd_sc_hd__nor2_2 _24179_ (.A(_19961_),
    .B(_19980_),
    .Y(_19981_));
 sky130_fd_sc_hd__nor2_2 _24180_ (.A(pcpi_rs2[17]),
    .B(_19518_),
    .Y(_19982_));
 sky130_fd_sc_hd__inv_2 _24181_ (.A(pcpi_rs2[17]),
    .Y(_02366_));
 sky130_fd_sc_hd__inv_2 _24182_ (.A(pcpi_rs1[17]),
    .Y(_19983_));
 sky130_fd_sc_hd__nor2_2 _24183_ (.A(_02366_),
    .B(_19983_),
    .Y(_19984_));
 sky130_fd_sc_hd__nor2_2 _24184_ (.A(_19982_),
    .B(_19984_),
    .Y(_19985_));
 sky130_fd_sc_hd__inv_2 _24185_ (.A(_19985_),
    .Y(_19986_));
 sky130_fd_sc_hd__nor2_2 _24186_ (.A(pcpi_rs2[19]),
    .B(_19515_),
    .Y(_19987_));
 sky130_fd_sc_hd__inv_2 _24187_ (.A(pcpi_rs2[19]),
    .Y(_02372_));
 sky130_fd_sc_hd__inv_2 _24188_ (.A(pcpi_rs1[19]),
    .Y(_19988_));
 sky130_fd_sc_hd__nor2_2 _24189_ (.A(_02372_),
    .B(_19988_),
    .Y(_19989_));
 sky130_fd_sc_hd__nor2_2 _24190_ (.A(_19987_),
    .B(_19989_),
    .Y(_19990_));
 sky130_fd_sc_hd__inv_2 _24191_ (.A(_19990_),
    .Y(_19991_));
 sky130_fd_sc_hd__nor2_2 _24192_ (.A(_19141_),
    .B(_19517_),
    .Y(_19992_));
 sky130_fd_sc_hd__inv_2 _24193_ (.A(_19141_),
    .Y(_02369_));
 sky130_fd_sc_hd__inv_2 _24194_ (.A(pcpi_rs1[18]),
    .Y(_19993_));
 sky130_fd_sc_hd__nor2_2 _24195_ (.A(_02369_),
    .B(_19993_),
    .Y(_19994_));
 sky130_fd_sc_hd__nor2_2 _24196_ (.A(_19992_),
    .B(_19994_),
    .Y(_19995_));
 sky130_fd_sc_hd__inv_2 _24197_ (.A(_19995_),
    .Y(_19996_));
 sky130_fd_sc_hd__xnor2_2 _24198_ (.A(pcpi_rs2[16]),
    .B(_19519_),
    .Y(_19997_));
 sky130_fd_sc_hd__and4_2 _24199_ (.A(_19986_),
    .B(_19991_),
    .C(_19996_),
    .D(_19997_),
    .X(_19998_));
 sky130_fd_sc_hd__and4b_2 _24200_ (.A_N(_19924_),
    .B(_19943_),
    .C(_19981_),
    .D(_19998_),
    .X(_19999_));
 sky130_fd_sc_hd__buf_1 _24201_ (.A(_19999_),
    .X(_00000_));
 sky130_fd_sc_hd__o211a_2 _24202_ (.A1(pcpi_insn[13]),
    .A2(pcpi_insn[12]),
    .B1(_18161_),
    .C1(_18169_),
    .X(\pcpi_mul.instr_any_mulh ));
 sky130_fd_sc_hd__or3_2 _24203_ (.A(instr_slt),
    .B(instr_slti),
    .C(instr_blt),
    .X(_00006_));
 sky130_fd_sc_hd__or3_2 _24204_ (.A(instr_sltu),
    .B(instr_sltiu),
    .C(instr_bltu),
    .X(_00007_));
 sky130_fd_sc_hd__nand2_2 _24205_ (.A(_18008_),
    .B(_18053_),
    .Y(_00299_));
 sky130_fd_sc_hd__or3_2 _24206_ (.A(_18048_),
    .B(_00319_),
    .C(_00317_),
    .X(_20000_));
 sky130_fd_sc_hd__and3_2 _24207_ (.A(_18014_),
    .B(_18015_),
    .C(_18255_),
    .X(_20001_));
 sky130_fd_sc_hd__a211oi_2 _24208_ (.A1(_18204_),
    .A2(_00297_),
    .B1(_20000_),
    .C1(_20001_),
    .Y(_20002_));
 sky130_fd_sc_hd__nor2_2 _24209_ (.A(mem_do_wdata),
    .B(_18051_),
    .Y(_20003_));
 sky130_fd_sc_hd__or2_2 _24210_ (.A(instr_lhu),
    .B(instr_lh),
    .X(_20004_));
 sky130_fd_sc_hd__a32o_2 _24211_ (.A1(instr_sh),
    .A2(\cpu_state[5] ),
    .A3(_20003_),
    .B1(_18449_),
    .B2(_20004_),
    .X(_20005_));
 sky130_fd_sc_hd__a2bb2o_2 _24212_ (.A1_N(_19796_),
    .A2_N(_20002_),
    .B1(_18448_),
    .B2(_20005_),
    .X(_00047_));
 sky130_fd_sc_hd__buf_1 _24213_ (.A(_18444_),
    .X(_20006_));
 sky130_fd_sc_hd__and3_2 _24214_ (.A(_18188_),
    .B(_20006_),
    .C(_19500_),
    .X(_00336_));
 sky130_fd_sc_hd__o21ai_2 _24215_ (.A1(mem_do_rinst),
    .A2(_18447_),
    .B1(_18056_),
    .Y(_00338_));
 sky130_fd_sc_hd__inv_2 _24216_ (.A(alu_eq),
    .Y(_00340_));
 sky130_fd_sc_hd__nor2_2 _24217_ (.A(instr_bne),
    .B(is_slti_blt_slt),
    .Y(_20007_));
 sky130_fd_sc_hd__and3b_2 _24218_ (.A_N(is_sltiu_bltu_sltu),
    .B(_18210_),
    .C(_20007_),
    .X(_00341_));
 sky130_fd_sc_hd__nand2_2 _24219_ (.A(is_slti_blt_slt),
    .B(alu_lts),
    .Y(_20008_));
 sky130_fd_sc_hd__o221a_2 _24220_ (.A1(alu_eq),
    .A2(_18432_),
    .B1(_18424_),
    .B2(alu_ltu),
    .C1(_20008_),
    .X(_20009_));
 sky130_fd_sc_hd__or2b_2 _24221_ (.A(alu_lts),
    .B_N(instr_bge),
    .X(_20010_));
 sky130_fd_sc_hd__nand2_2 _24222_ (.A(is_sltiu_bltu_sltu),
    .B(alu_ltu),
    .Y(_20011_));
 sky130_fd_sc_hd__and3_2 _24223_ (.A(_20009_),
    .B(_20010_),
    .C(_20011_),
    .X(_00342_));
 sky130_fd_sc_hd__nand2_2 _24224_ (.A(_20587_),
    .B(_00343_),
    .Y(_00344_));
 sky130_fd_sc_hd__o22ai_2 _24225_ (.A1(_00346_),
    .A2(_18188_),
    .B1(_00339_),
    .B2(_00297_),
    .Y(_00347_));
 sky130_fd_sc_hd__nor2_2 _24226_ (.A(_18243_),
    .B(_18149_),
    .Y(_00349_));
 sky130_fd_sc_hd__and2_2 _24227_ (.A(_02410_),
    .B(_00349_),
    .X(_00351_));
 sky130_fd_sc_hd__o21a_2 _24228_ (.A1(_18188_),
    .A2(_18447_),
    .B1(_18443_),
    .X(_00355_));
 sky130_fd_sc_hd__inv_2 _24229_ (.A(\decoded_imm_uj[4] ),
    .Y(_00367_));
 sky130_fd_sc_hd__inv_2 _24230_ (.A(\cpuregs[0][1] ),
    .Y(_00371_));
 sky130_fd_sc_hd__inv_2 _24231_ (.A(\cpuregs[1][1] ),
    .Y(_00372_));
 sky130_fd_sc_hd__inv_2 _24232_ (.A(\cpuregs[2][1] ),
    .Y(_00373_));
 sky130_fd_sc_hd__inv_2 _24233_ (.A(\cpuregs[3][1] ),
    .Y(_00374_));
 sky130_fd_sc_hd__inv_2 _24234_ (.A(\cpuregs[4][1] ),
    .Y(_00376_));
 sky130_fd_sc_hd__inv_2 _24235_ (.A(\cpuregs[5][1] ),
    .Y(_00377_));
 sky130_fd_sc_hd__inv_2 _24236_ (.A(\cpuregs[6][1] ),
    .Y(_00378_));
 sky130_fd_sc_hd__inv_2 _24237_ (.A(\cpuregs[7][1] ),
    .Y(_00379_));
 sky130_fd_sc_hd__inv_2 _24238_ (.A(\cpuregs[8][1] ),
    .Y(_00381_));
 sky130_fd_sc_hd__inv_2 _24239_ (.A(\cpuregs[9][1] ),
    .Y(_00382_));
 sky130_fd_sc_hd__inv_2 _24240_ (.A(\cpuregs[10][1] ),
    .Y(_00383_));
 sky130_fd_sc_hd__inv_2 _24241_ (.A(\cpuregs[11][1] ),
    .Y(_00384_));
 sky130_fd_sc_hd__inv_2 _24242_ (.A(\cpuregs[12][1] ),
    .Y(_00386_));
 sky130_fd_sc_hd__inv_2 _24243_ (.A(\cpuregs[13][1] ),
    .Y(_00387_));
 sky130_fd_sc_hd__inv_2 _24244_ (.A(\cpuregs[14][1] ),
    .Y(_00388_));
 sky130_fd_sc_hd__inv_2 _24245_ (.A(\cpuregs[15][1] ),
    .Y(_00389_));
 sky130_fd_sc_hd__inv_2 _24246_ (.A(\cpuregs[16][1] ),
    .Y(_00392_));
 sky130_fd_sc_hd__inv_2 _24247_ (.A(\cpuregs[17][1] ),
    .Y(_00393_));
 sky130_fd_sc_hd__inv_2 _24248_ (.A(\cpuregs[18][1] ),
    .Y(_00394_));
 sky130_fd_sc_hd__inv_2 _24249_ (.A(\cpuregs[19][1] ),
    .Y(_00395_));
 sky130_fd_sc_hd__inv_2 _24250_ (.A(\cpuregs[0][2] ),
    .Y(_00398_));
 sky130_fd_sc_hd__inv_2 _24251_ (.A(\cpuregs[1][2] ),
    .Y(_00399_));
 sky130_fd_sc_hd__inv_2 _24252_ (.A(\cpuregs[2][2] ),
    .Y(_00400_));
 sky130_fd_sc_hd__inv_2 _24253_ (.A(\cpuregs[3][2] ),
    .Y(_00401_));
 sky130_fd_sc_hd__inv_2 _24254_ (.A(\cpuregs[4][2] ),
    .Y(_00403_));
 sky130_fd_sc_hd__inv_2 _24255_ (.A(\cpuregs[5][2] ),
    .Y(_00404_));
 sky130_fd_sc_hd__inv_2 _24256_ (.A(\cpuregs[6][2] ),
    .Y(_00405_));
 sky130_fd_sc_hd__inv_2 _24257_ (.A(\cpuregs[7][2] ),
    .Y(_00406_));
 sky130_fd_sc_hd__inv_2 _24258_ (.A(\cpuregs[8][2] ),
    .Y(_00408_));
 sky130_fd_sc_hd__inv_2 _24259_ (.A(\cpuregs[9][2] ),
    .Y(_00409_));
 sky130_fd_sc_hd__inv_2 _24260_ (.A(\cpuregs[10][2] ),
    .Y(_00410_));
 sky130_fd_sc_hd__inv_2 _24261_ (.A(\cpuregs[11][2] ),
    .Y(_00411_));
 sky130_fd_sc_hd__inv_2 _24262_ (.A(\cpuregs[12][2] ),
    .Y(_00413_));
 sky130_fd_sc_hd__inv_2 _24263_ (.A(\cpuregs[13][2] ),
    .Y(_00414_));
 sky130_fd_sc_hd__inv_2 _24264_ (.A(\cpuregs[14][2] ),
    .Y(_00415_));
 sky130_fd_sc_hd__inv_2 _24265_ (.A(\cpuregs[15][2] ),
    .Y(_00416_));
 sky130_fd_sc_hd__inv_2 _24266_ (.A(\cpuregs[16][2] ),
    .Y(_00419_));
 sky130_fd_sc_hd__inv_2 _24267_ (.A(\cpuregs[17][2] ),
    .Y(_00420_));
 sky130_fd_sc_hd__inv_2 _24268_ (.A(\cpuregs[18][2] ),
    .Y(_00421_));
 sky130_fd_sc_hd__inv_2 _24269_ (.A(\cpuregs[19][2] ),
    .Y(_00422_));
 sky130_fd_sc_hd__inv_2 _24270_ (.A(\cpuregs[0][3] ),
    .Y(_00425_));
 sky130_fd_sc_hd__inv_2 _24271_ (.A(\cpuregs[1][3] ),
    .Y(_00426_));
 sky130_fd_sc_hd__inv_2 _24272_ (.A(\cpuregs[2][3] ),
    .Y(_00427_));
 sky130_fd_sc_hd__inv_2 _24273_ (.A(\cpuregs[3][3] ),
    .Y(_00428_));
 sky130_fd_sc_hd__inv_2 _24274_ (.A(\cpuregs[4][3] ),
    .Y(_00430_));
 sky130_fd_sc_hd__inv_2 _24275_ (.A(\cpuregs[5][3] ),
    .Y(_00431_));
 sky130_fd_sc_hd__inv_2 _24276_ (.A(\cpuregs[6][3] ),
    .Y(_00432_));
 sky130_fd_sc_hd__inv_2 _24277_ (.A(\cpuregs[7][3] ),
    .Y(_00433_));
 sky130_fd_sc_hd__inv_2 _24278_ (.A(\cpuregs[8][3] ),
    .Y(_00435_));
 sky130_fd_sc_hd__inv_2 _24279_ (.A(\cpuregs[9][3] ),
    .Y(_00436_));
 sky130_fd_sc_hd__inv_2 _24280_ (.A(\cpuregs[10][3] ),
    .Y(_00437_));
 sky130_fd_sc_hd__inv_2 _24281_ (.A(\cpuregs[11][3] ),
    .Y(_00438_));
 sky130_fd_sc_hd__inv_2 _24282_ (.A(\cpuregs[12][3] ),
    .Y(_00440_));
 sky130_fd_sc_hd__inv_2 _24283_ (.A(\cpuregs[13][3] ),
    .Y(_00441_));
 sky130_fd_sc_hd__inv_2 _24284_ (.A(\cpuregs[14][3] ),
    .Y(_00442_));
 sky130_fd_sc_hd__inv_2 _24285_ (.A(\cpuregs[15][3] ),
    .Y(_00443_));
 sky130_fd_sc_hd__inv_2 _24286_ (.A(\cpuregs[16][3] ),
    .Y(_00446_));
 sky130_fd_sc_hd__inv_2 _24287_ (.A(\cpuregs[17][3] ),
    .Y(_00447_));
 sky130_fd_sc_hd__inv_2 _24288_ (.A(\cpuregs[18][3] ),
    .Y(_00448_));
 sky130_fd_sc_hd__inv_2 _24289_ (.A(\cpuregs[19][3] ),
    .Y(_00449_));
 sky130_fd_sc_hd__inv_2 _24290_ (.A(\cpuregs[0][4] ),
    .Y(_00452_));
 sky130_fd_sc_hd__inv_2 _24291_ (.A(\cpuregs[1][4] ),
    .Y(_00453_));
 sky130_fd_sc_hd__inv_2 _24292_ (.A(\cpuregs[2][4] ),
    .Y(_00454_));
 sky130_fd_sc_hd__inv_2 _24293_ (.A(\cpuregs[3][4] ),
    .Y(_00455_));
 sky130_fd_sc_hd__inv_2 _24294_ (.A(\cpuregs[4][4] ),
    .Y(_00457_));
 sky130_fd_sc_hd__inv_2 _24295_ (.A(\cpuregs[5][4] ),
    .Y(_00458_));
 sky130_fd_sc_hd__inv_2 _24296_ (.A(\cpuregs[6][4] ),
    .Y(_00459_));
 sky130_fd_sc_hd__inv_2 _24297_ (.A(\cpuregs[7][4] ),
    .Y(_00460_));
 sky130_fd_sc_hd__inv_2 _24298_ (.A(\cpuregs[8][4] ),
    .Y(_00462_));
 sky130_fd_sc_hd__inv_2 _24299_ (.A(\cpuregs[9][4] ),
    .Y(_00463_));
 sky130_fd_sc_hd__inv_2 _24300_ (.A(\cpuregs[10][4] ),
    .Y(_00464_));
 sky130_fd_sc_hd__inv_2 _24301_ (.A(\cpuregs[11][4] ),
    .Y(_00465_));
 sky130_fd_sc_hd__inv_2 _24302_ (.A(\cpuregs[12][4] ),
    .Y(_00467_));
 sky130_fd_sc_hd__inv_2 _24303_ (.A(\cpuregs[13][4] ),
    .Y(_00468_));
 sky130_fd_sc_hd__inv_2 _24304_ (.A(\cpuregs[14][4] ),
    .Y(_00469_));
 sky130_fd_sc_hd__inv_2 _24305_ (.A(\cpuregs[15][4] ),
    .Y(_00470_));
 sky130_fd_sc_hd__inv_2 _24306_ (.A(\cpuregs[16][4] ),
    .Y(_00473_));
 sky130_fd_sc_hd__inv_2 _24307_ (.A(\cpuregs[17][4] ),
    .Y(_00474_));
 sky130_fd_sc_hd__inv_2 _24308_ (.A(\cpuregs[18][4] ),
    .Y(_00475_));
 sky130_fd_sc_hd__inv_2 _24309_ (.A(\cpuregs[19][4] ),
    .Y(_00476_));
 sky130_fd_sc_hd__inv_2 _24310_ (.A(\cpuregs[0][5] ),
    .Y(_00479_));
 sky130_fd_sc_hd__inv_2 _24311_ (.A(\cpuregs[1][5] ),
    .Y(_00480_));
 sky130_fd_sc_hd__inv_2 _24312_ (.A(\cpuregs[2][5] ),
    .Y(_00481_));
 sky130_fd_sc_hd__inv_2 _24313_ (.A(\cpuregs[3][5] ),
    .Y(_00482_));
 sky130_fd_sc_hd__inv_2 _24314_ (.A(\cpuregs[4][5] ),
    .Y(_00484_));
 sky130_fd_sc_hd__inv_2 _24315_ (.A(\cpuregs[5][5] ),
    .Y(_00485_));
 sky130_fd_sc_hd__inv_2 _24316_ (.A(\cpuregs[6][5] ),
    .Y(_00486_));
 sky130_fd_sc_hd__inv_2 _24317_ (.A(\cpuregs[7][5] ),
    .Y(_00487_));
 sky130_fd_sc_hd__inv_2 _24318_ (.A(\cpuregs[8][5] ),
    .Y(_00489_));
 sky130_fd_sc_hd__inv_2 _24319_ (.A(\cpuregs[9][5] ),
    .Y(_00490_));
 sky130_fd_sc_hd__inv_2 _24320_ (.A(\cpuregs[10][5] ),
    .Y(_00491_));
 sky130_fd_sc_hd__inv_2 _24321_ (.A(\cpuregs[11][5] ),
    .Y(_00492_));
 sky130_fd_sc_hd__inv_2 _24322_ (.A(\cpuregs[12][5] ),
    .Y(_00494_));
 sky130_fd_sc_hd__inv_2 _24323_ (.A(\cpuregs[13][5] ),
    .Y(_00495_));
 sky130_fd_sc_hd__inv_2 _24324_ (.A(\cpuregs[14][5] ),
    .Y(_00496_));
 sky130_fd_sc_hd__inv_2 _24325_ (.A(\cpuregs[15][5] ),
    .Y(_00497_));
 sky130_fd_sc_hd__inv_2 _24326_ (.A(\cpuregs[16][5] ),
    .Y(_00500_));
 sky130_fd_sc_hd__inv_2 _24327_ (.A(\cpuregs[17][5] ),
    .Y(_00501_));
 sky130_fd_sc_hd__inv_2 _24328_ (.A(\cpuregs[18][5] ),
    .Y(_00502_));
 sky130_fd_sc_hd__inv_2 _24329_ (.A(\cpuregs[19][5] ),
    .Y(_00503_));
 sky130_fd_sc_hd__inv_2 _24330_ (.A(\cpuregs[0][6] ),
    .Y(_00506_));
 sky130_fd_sc_hd__inv_2 _24331_ (.A(\cpuregs[1][6] ),
    .Y(_00507_));
 sky130_fd_sc_hd__inv_2 _24332_ (.A(\cpuregs[2][6] ),
    .Y(_00508_));
 sky130_fd_sc_hd__inv_2 _24333_ (.A(\cpuregs[3][6] ),
    .Y(_00509_));
 sky130_fd_sc_hd__inv_2 _24334_ (.A(\cpuregs[4][6] ),
    .Y(_00511_));
 sky130_fd_sc_hd__inv_2 _24335_ (.A(\cpuregs[5][6] ),
    .Y(_00512_));
 sky130_fd_sc_hd__inv_2 _24336_ (.A(\cpuregs[6][6] ),
    .Y(_00513_));
 sky130_fd_sc_hd__inv_2 _24337_ (.A(\cpuregs[7][6] ),
    .Y(_00514_));
 sky130_fd_sc_hd__inv_2 _24338_ (.A(\cpuregs[8][6] ),
    .Y(_00516_));
 sky130_fd_sc_hd__inv_2 _24339_ (.A(\cpuregs[9][6] ),
    .Y(_00517_));
 sky130_fd_sc_hd__inv_2 _24340_ (.A(\cpuregs[10][6] ),
    .Y(_00518_));
 sky130_fd_sc_hd__inv_2 _24341_ (.A(\cpuregs[11][6] ),
    .Y(_00519_));
 sky130_fd_sc_hd__inv_2 _24342_ (.A(\cpuregs[12][6] ),
    .Y(_00521_));
 sky130_fd_sc_hd__inv_2 _24343_ (.A(\cpuregs[13][6] ),
    .Y(_00522_));
 sky130_fd_sc_hd__inv_2 _24344_ (.A(\cpuregs[14][6] ),
    .Y(_00523_));
 sky130_fd_sc_hd__inv_2 _24345_ (.A(\cpuregs[15][6] ),
    .Y(_00524_));
 sky130_fd_sc_hd__inv_2 _24346_ (.A(\cpuregs[16][6] ),
    .Y(_00527_));
 sky130_fd_sc_hd__inv_2 _24347_ (.A(\cpuregs[17][6] ),
    .Y(_00528_));
 sky130_fd_sc_hd__inv_2 _24348_ (.A(\cpuregs[18][6] ),
    .Y(_00529_));
 sky130_fd_sc_hd__inv_2 _24349_ (.A(\cpuregs[19][6] ),
    .Y(_00530_));
 sky130_fd_sc_hd__inv_2 _24350_ (.A(\cpuregs[0][7] ),
    .Y(_00533_));
 sky130_fd_sc_hd__inv_2 _24351_ (.A(\cpuregs[1][7] ),
    .Y(_00534_));
 sky130_fd_sc_hd__inv_2 _24352_ (.A(\cpuregs[2][7] ),
    .Y(_00535_));
 sky130_fd_sc_hd__inv_2 _24353_ (.A(\cpuregs[3][7] ),
    .Y(_00536_));
 sky130_fd_sc_hd__inv_2 _24354_ (.A(\cpuregs[4][7] ),
    .Y(_00538_));
 sky130_fd_sc_hd__inv_2 _24355_ (.A(\cpuregs[5][7] ),
    .Y(_00539_));
 sky130_fd_sc_hd__inv_2 _24356_ (.A(\cpuregs[6][7] ),
    .Y(_00540_));
 sky130_fd_sc_hd__inv_2 _24357_ (.A(\cpuregs[7][7] ),
    .Y(_00541_));
 sky130_fd_sc_hd__inv_2 _24358_ (.A(\cpuregs[8][7] ),
    .Y(_00543_));
 sky130_fd_sc_hd__inv_2 _24359_ (.A(\cpuregs[9][7] ),
    .Y(_00544_));
 sky130_fd_sc_hd__inv_2 _24360_ (.A(\cpuregs[10][7] ),
    .Y(_00545_));
 sky130_fd_sc_hd__inv_2 _24361_ (.A(\cpuregs[11][7] ),
    .Y(_00546_));
 sky130_fd_sc_hd__inv_2 _24362_ (.A(\cpuregs[12][7] ),
    .Y(_00548_));
 sky130_fd_sc_hd__inv_2 _24363_ (.A(\cpuregs[13][7] ),
    .Y(_00549_));
 sky130_fd_sc_hd__inv_2 _24364_ (.A(\cpuregs[14][7] ),
    .Y(_00550_));
 sky130_fd_sc_hd__inv_2 _24365_ (.A(\cpuregs[15][7] ),
    .Y(_00551_));
 sky130_fd_sc_hd__inv_2 _24366_ (.A(\cpuregs[16][7] ),
    .Y(_00554_));
 sky130_fd_sc_hd__inv_2 _24367_ (.A(\cpuregs[17][7] ),
    .Y(_00555_));
 sky130_fd_sc_hd__inv_2 _24368_ (.A(\cpuregs[18][7] ),
    .Y(_00556_));
 sky130_fd_sc_hd__inv_2 _24369_ (.A(\cpuregs[19][7] ),
    .Y(_00557_));
 sky130_fd_sc_hd__inv_2 _24370_ (.A(\cpuregs[0][8] ),
    .Y(_00560_));
 sky130_fd_sc_hd__inv_2 _24371_ (.A(\cpuregs[1][8] ),
    .Y(_00561_));
 sky130_fd_sc_hd__inv_2 _24372_ (.A(\cpuregs[2][8] ),
    .Y(_00562_));
 sky130_fd_sc_hd__inv_2 _24373_ (.A(\cpuregs[3][8] ),
    .Y(_00563_));
 sky130_fd_sc_hd__inv_2 _24374_ (.A(\cpuregs[4][8] ),
    .Y(_00565_));
 sky130_fd_sc_hd__inv_2 _24375_ (.A(\cpuregs[5][8] ),
    .Y(_00566_));
 sky130_fd_sc_hd__inv_2 _24376_ (.A(\cpuregs[6][8] ),
    .Y(_00567_));
 sky130_fd_sc_hd__inv_2 _24377_ (.A(\cpuregs[7][8] ),
    .Y(_00568_));
 sky130_fd_sc_hd__inv_2 _24378_ (.A(\cpuregs[8][8] ),
    .Y(_00570_));
 sky130_fd_sc_hd__inv_2 _24379_ (.A(\cpuregs[9][8] ),
    .Y(_00571_));
 sky130_fd_sc_hd__inv_2 _24380_ (.A(\cpuregs[10][8] ),
    .Y(_00572_));
 sky130_fd_sc_hd__inv_2 _24381_ (.A(\cpuregs[11][8] ),
    .Y(_00573_));
 sky130_fd_sc_hd__inv_2 _24382_ (.A(\cpuregs[12][8] ),
    .Y(_00575_));
 sky130_fd_sc_hd__inv_2 _24383_ (.A(\cpuregs[13][8] ),
    .Y(_00576_));
 sky130_fd_sc_hd__inv_2 _24384_ (.A(\cpuregs[14][8] ),
    .Y(_00577_));
 sky130_fd_sc_hd__inv_2 _24385_ (.A(\cpuregs[15][8] ),
    .Y(_00578_));
 sky130_fd_sc_hd__inv_2 _24386_ (.A(\cpuregs[16][8] ),
    .Y(_00581_));
 sky130_fd_sc_hd__inv_2 _24387_ (.A(\cpuregs[17][8] ),
    .Y(_00582_));
 sky130_fd_sc_hd__inv_2 _24388_ (.A(\cpuregs[18][8] ),
    .Y(_00583_));
 sky130_fd_sc_hd__inv_2 _24389_ (.A(\cpuregs[19][8] ),
    .Y(_00584_));
 sky130_fd_sc_hd__inv_2 _24390_ (.A(\cpuregs[0][9] ),
    .Y(_00587_));
 sky130_fd_sc_hd__inv_2 _24391_ (.A(\cpuregs[1][9] ),
    .Y(_00588_));
 sky130_fd_sc_hd__inv_2 _24392_ (.A(\cpuregs[2][9] ),
    .Y(_00589_));
 sky130_fd_sc_hd__inv_2 _24393_ (.A(\cpuregs[3][9] ),
    .Y(_00590_));
 sky130_fd_sc_hd__inv_2 _24394_ (.A(\cpuregs[4][9] ),
    .Y(_00592_));
 sky130_fd_sc_hd__inv_2 _24395_ (.A(\cpuregs[5][9] ),
    .Y(_00593_));
 sky130_fd_sc_hd__inv_2 _24396_ (.A(\cpuregs[6][9] ),
    .Y(_00594_));
 sky130_fd_sc_hd__inv_2 _24397_ (.A(\cpuregs[7][9] ),
    .Y(_00595_));
 sky130_fd_sc_hd__inv_2 _24398_ (.A(\cpuregs[8][9] ),
    .Y(_00597_));
 sky130_fd_sc_hd__inv_2 _24399_ (.A(\cpuregs[9][9] ),
    .Y(_00598_));
 sky130_fd_sc_hd__inv_2 _24400_ (.A(\cpuregs[10][9] ),
    .Y(_00599_));
 sky130_fd_sc_hd__inv_2 _24401_ (.A(\cpuregs[11][9] ),
    .Y(_00600_));
 sky130_fd_sc_hd__inv_2 _24402_ (.A(\cpuregs[12][9] ),
    .Y(_00602_));
 sky130_fd_sc_hd__inv_2 _24403_ (.A(\cpuregs[13][9] ),
    .Y(_00603_));
 sky130_fd_sc_hd__inv_2 _24404_ (.A(\cpuregs[14][9] ),
    .Y(_00604_));
 sky130_fd_sc_hd__inv_2 _24405_ (.A(\cpuregs[15][9] ),
    .Y(_00605_));
 sky130_fd_sc_hd__inv_2 _24406_ (.A(\cpuregs[16][9] ),
    .Y(_00608_));
 sky130_fd_sc_hd__inv_2 _24407_ (.A(\cpuregs[17][9] ),
    .Y(_00609_));
 sky130_fd_sc_hd__inv_2 _24408_ (.A(\cpuregs[18][9] ),
    .Y(_00610_));
 sky130_fd_sc_hd__inv_2 _24409_ (.A(\cpuregs[19][9] ),
    .Y(_00611_));
 sky130_fd_sc_hd__inv_2 _24410_ (.A(\cpuregs[0][10] ),
    .Y(_00614_));
 sky130_fd_sc_hd__inv_2 _24411_ (.A(\cpuregs[1][10] ),
    .Y(_00615_));
 sky130_fd_sc_hd__inv_2 _24412_ (.A(\cpuregs[2][10] ),
    .Y(_00616_));
 sky130_fd_sc_hd__inv_2 _24413_ (.A(\cpuregs[3][10] ),
    .Y(_00617_));
 sky130_fd_sc_hd__inv_2 _24414_ (.A(\cpuregs[4][10] ),
    .Y(_00619_));
 sky130_fd_sc_hd__inv_2 _24415_ (.A(\cpuregs[5][10] ),
    .Y(_00620_));
 sky130_fd_sc_hd__inv_2 _24416_ (.A(\cpuregs[6][10] ),
    .Y(_00621_));
 sky130_fd_sc_hd__inv_2 _24417_ (.A(\cpuregs[7][10] ),
    .Y(_00622_));
 sky130_fd_sc_hd__inv_2 _24418_ (.A(\cpuregs[8][10] ),
    .Y(_00624_));
 sky130_fd_sc_hd__inv_2 _24419_ (.A(\cpuregs[9][10] ),
    .Y(_00625_));
 sky130_fd_sc_hd__inv_2 _24420_ (.A(\cpuregs[10][10] ),
    .Y(_00626_));
 sky130_fd_sc_hd__inv_2 _24421_ (.A(\cpuregs[11][10] ),
    .Y(_00627_));
 sky130_fd_sc_hd__inv_2 _24422_ (.A(\cpuregs[12][10] ),
    .Y(_00629_));
 sky130_fd_sc_hd__inv_2 _24423_ (.A(\cpuregs[13][10] ),
    .Y(_00630_));
 sky130_fd_sc_hd__inv_2 _24424_ (.A(\cpuregs[14][10] ),
    .Y(_00631_));
 sky130_fd_sc_hd__inv_2 _24425_ (.A(\cpuregs[15][10] ),
    .Y(_00632_));
 sky130_fd_sc_hd__inv_2 _24426_ (.A(\cpuregs[16][10] ),
    .Y(_00635_));
 sky130_fd_sc_hd__inv_2 _24427_ (.A(\cpuregs[17][10] ),
    .Y(_00636_));
 sky130_fd_sc_hd__inv_2 _24428_ (.A(\cpuregs[18][10] ),
    .Y(_00637_));
 sky130_fd_sc_hd__inv_2 _24429_ (.A(\cpuregs[19][10] ),
    .Y(_00638_));
 sky130_fd_sc_hd__inv_2 _24430_ (.A(\cpuregs[0][11] ),
    .Y(_00641_));
 sky130_fd_sc_hd__inv_2 _24431_ (.A(\cpuregs[1][11] ),
    .Y(_00642_));
 sky130_fd_sc_hd__inv_2 _24432_ (.A(\cpuregs[2][11] ),
    .Y(_00643_));
 sky130_fd_sc_hd__inv_2 _24433_ (.A(\cpuregs[3][11] ),
    .Y(_00644_));
 sky130_fd_sc_hd__inv_2 _24434_ (.A(\cpuregs[4][11] ),
    .Y(_00646_));
 sky130_fd_sc_hd__inv_2 _24435_ (.A(\cpuregs[5][11] ),
    .Y(_00647_));
 sky130_fd_sc_hd__inv_2 _24436_ (.A(\cpuregs[6][11] ),
    .Y(_00648_));
 sky130_fd_sc_hd__inv_2 _24437_ (.A(\cpuregs[7][11] ),
    .Y(_00649_));
 sky130_fd_sc_hd__inv_2 _24438_ (.A(\cpuregs[8][11] ),
    .Y(_00651_));
 sky130_fd_sc_hd__inv_2 _24439_ (.A(\cpuregs[9][11] ),
    .Y(_00652_));
 sky130_fd_sc_hd__inv_2 _24440_ (.A(\cpuregs[10][11] ),
    .Y(_00653_));
 sky130_fd_sc_hd__inv_2 _24441_ (.A(\cpuregs[11][11] ),
    .Y(_00654_));
 sky130_fd_sc_hd__inv_2 _24442_ (.A(\cpuregs[12][11] ),
    .Y(_00656_));
 sky130_fd_sc_hd__inv_2 _24443_ (.A(\cpuregs[13][11] ),
    .Y(_00657_));
 sky130_fd_sc_hd__inv_2 _24444_ (.A(\cpuregs[14][11] ),
    .Y(_00658_));
 sky130_fd_sc_hd__inv_2 _24445_ (.A(\cpuregs[15][11] ),
    .Y(_00659_));
 sky130_fd_sc_hd__inv_2 _24446_ (.A(\cpuregs[16][11] ),
    .Y(_00662_));
 sky130_fd_sc_hd__inv_2 _24447_ (.A(\cpuregs[17][11] ),
    .Y(_00663_));
 sky130_fd_sc_hd__inv_2 _24448_ (.A(\cpuregs[18][11] ),
    .Y(_00664_));
 sky130_fd_sc_hd__inv_2 _24449_ (.A(\cpuregs[19][11] ),
    .Y(_00665_));
 sky130_fd_sc_hd__inv_2 _24450_ (.A(\cpuregs[0][12] ),
    .Y(_00668_));
 sky130_fd_sc_hd__inv_2 _24451_ (.A(\cpuregs[1][12] ),
    .Y(_00669_));
 sky130_fd_sc_hd__inv_2 _24452_ (.A(\cpuregs[2][12] ),
    .Y(_00670_));
 sky130_fd_sc_hd__inv_2 _24453_ (.A(\cpuregs[3][12] ),
    .Y(_00671_));
 sky130_fd_sc_hd__inv_2 _24454_ (.A(\cpuregs[4][12] ),
    .Y(_00673_));
 sky130_fd_sc_hd__inv_2 _24455_ (.A(\cpuregs[5][12] ),
    .Y(_00674_));
 sky130_fd_sc_hd__inv_2 _24456_ (.A(\cpuregs[6][12] ),
    .Y(_00675_));
 sky130_fd_sc_hd__inv_2 _24457_ (.A(\cpuregs[7][12] ),
    .Y(_00676_));
 sky130_fd_sc_hd__inv_2 _24458_ (.A(\cpuregs[8][12] ),
    .Y(_00678_));
 sky130_fd_sc_hd__inv_2 _24459_ (.A(\cpuregs[9][12] ),
    .Y(_00679_));
 sky130_fd_sc_hd__inv_2 _24460_ (.A(\cpuregs[10][12] ),
    .Y(_00680_));
 sky130_fd_sc_hd__inv_2 _24461_ (.A(\cpuregs[11][12] ),
    .Y(_00681_));
 sky130_fd_sc_hd__inv_2 _24462_ (.A(\cpuregs[12][12] ),
    .Y(_00683_));
 sky130_fd_sc_hd__inv_2 _24463_ (.A(\cpuregs[13][12] ),
    .Y(_00684_));
 sky130_fd_sc_hd__inv_2 _24464_ (.A(\cpuregs[14][12] ),
    .Y(_00685_));
 sky130_fd_sc_hd__inv_2 _24465_ (.A(\cpuregs[15][12] ),
    .Y(_00686_));
 sky130_fd_sc_hd__inv_2 _24466_ (.A(\cpuregs[16][12] ),
    .Y(_00689_));
 sky130_fd_sc_hd__inv_2 _24467_ (.A(\cpuregs[17][12] ),
    .Y(_00690_));
 sky130_fd_sc_hd__inv_2 _24468_ (.A(\cpuregs[18][12] ),
    .Y(_00691_));
 sky130_fd_sc_hd__inv_2 _24469_ (.A(\cpuregs[19][12] ),
    .Y(_00692_));
 sky130_fd_sc_hd__inv_2 _24470_ (.A(\cpuregs[0][13] ),
    .Y(_00695_));
 sky130_fd_sc_hd__inv_2 _24471_ (.A(\cpuregs[1][13] ),
    .Y(_00696_));
 sky130_fd_sc_hd__inv_2 _24472_ (.A(\cpuregs[2][13] ),
    .Y(_00697_));
 sky130_fd_sc_hd__inv_2 _24473_ (.A(\cpuregs[3][13] ),
    .Y(_00698_));
 sky130_fd_sc_hd__inv_2 _24474_ (.A(\cpuregs[4][13] ),
    .Y(_00700_));
 sky130_fd_sc_hd__inv_2 _24475_ (.A(\cpuregs[5][13] ),
    .Y(_00701_));
 sky130_fd_sc_hd__inv_2 _24476_ (.A(\cpuregs[6][13] ),
    .Y(_00702_));
 sky130_fd_sc_hd__inv_2 _24477_ (.A(\cpuregs[7][13] ),
    .Y(_00703_));
 sky130_fd_sc_hd__inv_2 _24478_ (.A(\cpuregs[8][13] ),
    .Y(_00705_));
 sky130_fd_sc_hd__inv_2 _24479_ (.A(\cpuregs[9][13] ),
    .Y(_00706_));
 sky130_fd_sc_hd__inv_2 _24480_ (.A(\cpuregs[10][13] ),
    .Y(_00707_));
 sky130_fd_sc_hd__inv_2 _24481_ (.A(\cpuregs[11][13] ),
    .Y(_00708_));
 sky130_fd_sc_hd__inv_2 _24482_ (.A(\cpuregs[12][13] ),
    .Y(_00710_));
 sky130_fd_sc_hd__inv_2 _24483_ (.A(\cpuregs[13][13] ),
    .Y(_00711_));
 sky130_fd_sc_hd__inv_2 _24484_ (.A(\cpuregs[14][13] ),
    .Y(_00712_));
 sky130_fd_sc_hd__inv_2 _24485_ (.A(\cpuregs[15][13] ),
    .Y(_00713_));
 sky130_fd_sc_hd__inv_2 _24486_ (.A(\cpuregs[16][13] ),
    .Y(_00716_));
 sky130_fd_sc_hd__inv_2 _24487_ (.A(\cpuregs[17][13] ),
    .Y(_00717_));
 sky130_fd_sc_hd__inv_2 _24488_ (.A(\cpuregs[18][13] ),
    .Y(_00718_));
 sky130_fd_sc_hd__inv_2 _24489_ (.A(\cpuregs[19][13] ),
    .Y(_00719_));
 sky130_fd_sc_hd__inv_2 _24490_ (.A(\cpuregs[0][14] ),
    .Y(_00722_));
 sky130_fd_sc_hd__inv_2 _24491_ (.A(\cpuregs[1][14] ),
    .Y(_00723_));
 sky130_fd_sc_hd__inv_2 _24492_ (.A(\cpuregs[2][14] ),
    .Y(_00724_));
 sky130_fd_sc_hd__inv_2 _24493_ (.A(\cpuregs[3][14] ),
    .Y(_00725_));
 sky130_fd_sc_hd__inv_2 _24494_ (.A(\cpuregs[4][14] ),
    .Y(_00727_));
 sky130_fd_sc_hd__inv_2 _24495_ (.A(\cpuregs[5][14] ),
    .Y(_00728_));
 sky130_fd_sc_hd__inv_2 _24496_ (.A(\cpuregs[6][14] ),
    .Y(_00729_));
 sky130_fd_sc_hd__inv_2 _24497_ (.A(\cpuregs[7][14] ),
    .Y(_00730_));
 sky130_fd_sc_hd__inv_2 _24498_ (.A(\cpuregs[8][14] ),
    .Y(_00732_));
 sky130_fd_sc_hd__inv_2 _24499_ (.A(\cpuregs[9][14] ),
    .Y(_00733_));
 sky130_fd_sc_hd__inv_2 _24500_ (.A(\cpuregs[10][14] ),
    .Y(_00734_));
 sky130_fd_sc_hd__inv_2 _24501_ (.A(\cpuregs[11][14] ),
    .Y(_00735_));
 sky130_fd_sc_hd__inv_2 _24502_ (.A(\cpuregs[12][14] ),
    .Y(_00737_));
 sky130_fd_sc_hd__inv_2 _24503_ (.A(\cpuregs[13][14] ),
    .Y(_00738_));
 sky130_fd_sc_hd__inv_2 _24504_ (.A(\cpuregs[14][14] ),
    .Y(_00739_));
 sky130_fd_sc_hd__inv_2 _24505_ (.A(\cpuregs[15][14] ),
    .Y(_00740_));
 sky130_fd_sc_hd__inv_2 _24506_ (.A(\cpuregs[16][14] ),
    .Y(_00743_));
 sky130_fd_sc_hd__inv_2 _24507_ (.A(\cpuregs[17][14] ),
    .Y(_00744_));
 sky130_fd_sc_hd__inv_2 _24508_ (.A(\cpuregs[18][14] ),
    .Y(_00745_));
 sky130_fd_sc_hd__inv_2 _24509_ (.A(\cpuregs[19][14] ),
    .Y(_00746_));
 sky130_fd_sc_hd__inv_2 _24510_ (.A(\cpuregs[0][15] ),
    .Y(_00749_));
 sky130_fd_sc_hd__inv_2 _24511_ (.A(\cpuregs[1][15] ),
    .Y(_00750_));
 sky130_fd_sc_hd__inv_2 _24512_ (.A(\cpuregs[2][15] ),
    .Y(_00751_));
 sky130_fd_sc_hd__inv_2 _24513_ (.A(\cpuregs[3][15] ),
    .Y(_00752_));
 sky130_fd_sc_hd__inv_2 _24514_ (.A(\cpuregs[4][15] ),
    .Y(_00754_));
 sky130_fd_sc_hd__inv_2 _24515_ (.A(\cpuregs[5][15] ),
    .Y(_00755_));
 sky130_fd_sc_hd__inv_2 _24516_ (.A(\cpuregs[6][15] ),
    .Y(_00756_));
 sky130_fd_sc_hd__inv_2 _24517_ (.A(\cpuregs[7][15] ),
    .Y(_00757_));
 sky130_fd_sc_hd__inv_2 _24518_ (.A(\cpuregs[8][15] ),
    .Y(_00759_));
 sky130_fd_sc_hd__inv_2 _24519_ (.A(\cpuregs[9][15] ),
    .Y(_00760_));
 sky130_fd_sc_hd__inv_2 _24520_ (.A(\cpuregs[10][15] ),
    .Y(_00761_));
 sky130_fd_sc_hd__inv_2 _24521_ (.A(\cpuregs[11][15] ),
    .Y(_00762_));
 sky130_fd_sc_hd__inv_2 _24522_ (.A(\cpuregs[12][15] ),
    .Y(_00764_));
 sky130_fd_sc_hd__inv_2 _24523_ (.A(\cpuregs[13][15] ),
    .Y(_00765_));
 sky130_fd_sc_hd__inv_2 _24524_ (.A(\cpuregs[14][15] ),
    .Y(_00766_));
 sky130_fd_sc_hd__inv_2 _24525_ (.A(\cpuregs[15][15] ),
    .Y(_00767_));
 sky130_fd_sc_hd__inv_2 _24526_ (.A(\cpuregs[16][15] ),
    .Y(_00770_));
 sky130_fd_sc_hd__inv_2 _24527_ (.A(\cpuregs[17][15] ),
    .Y(_00771_));
 sky130_fd_sc_hd__inv_2 _24528_ (.A(\cpuregs[18][15] ),
    .Y(_00772_));
 sky130_fd_sc_hd__inv_2 _24529_ (.A(\cpuregs[19][15] ),
    .Y(_00773_));
 sky130_fd_sc_hd__inv_2 _24530_ (.A(\cpuregs[0][16] ),
    .Y(_00776_));
 sky130_fd_sc_hd__inv_2 _24531_ (.A(\cpuregs[1][16] ),
    .Y(_00777_));
 sky130_fd_sc_hd__inv_2 _24532_ (.A(\cpuregs[2][16] ),
    .Y(_00778_));
 sky130_fd_sc_hd__inv_2 _24533_ (.A(\cpuregs[3][16] ),
    .Y(_00779_));
 sky130_fd_sc_hd__inv_2 _24534_ (.A(\cpuregs[4][16] ),
    .Y(_00781_));
 sky130_fd_sc_hd__inv_2 _24535_ (.A(\cpuregs[5][16] ),
    .Y(_00782_));
 sky130_fd_sc_hd__inv_2 _24536_ (.A(\cpuregs[6][16] ),
    .Y(_00783_));
 sky130_fd_sc_hd__inv_2 _24537_ (.A(\cpuregs[7][16] ),
    .Y(_00784_));
 sky130_fd_sc_hd__inv_2 _24538_ (.A(\cpuregs[8][16] ),
    .Y(_00786_));
 sky130_fd_sc_hd__inv_2 _24539_ (.A(\cpuregs[9][16] ),
    .Y(_00787_));
 sky130_fd_sc_hd__inv_2 _24540_ (.A(\cpuregs[10][16] ),
    .Y(_00788_));
 sky130_fd_sc_hd__inv_2 _24541_ (.A(\cpuregs[11][16] ),
    .Y(_00789_));
 sky130_fd_sc_hd__inv_2 _24542_ (.A(\cpuregs[12][16] ),
    .Y(_00791_));
 sky130_fd_sc_hd__inv_2 _24543_ (.A(\cpuregs[13][16] ),
    .Y(_00792_));
 sky130_fd_sc_hd__inv_2 _24544_ (.A(\cpuregs[14][16] ),
    .Y(_00793_));
 sky130_fd_sc_hd__inv_2 _24545_ (.A(\cpuregs[15][16] ),
    .Y(_00794_));
 sky130_fd_sc_hd__inv_2 _24546_ (.A(\cpuregs[16][16] ),
    .Y(_00797_));
 sky130_fd_sc_hd__inv_2 _24547_ (.A(\cpuregs[17][16] ),
    .Y(_00798_));
 sky130_fd_sc_hd__inv_2 _24548_ (.A(\cpuregs[18][16] ),
    .Y(_00799_));
 sky130_fd_sc_hd__inv_2 _24549_ (.A(\cpuregs[19][16] ),
    .Y(_00800_));
 sky130_fd_sc_hd__inv_2 _24550_ (.A(\cpuregs[0][17] ),
    .Y(_00803_));
 sky130_fd_sc_hd__inv_2 _24551_ (.A(\cpuregs[1][17] ),
    .Y(_00804_));
 sky130_fd_sc_hd__inv_2 _24552_ (.A(\cpuregs[2][17] ),
    .Y(_00805_));
 sky130_fd_sc_hd__inv_2 _24553_ (.A(\cpuregs[3][17] ),
    .Y(_00806_));
 sky130_fd_sc_hd__inv_2 _24554_ (.A(\cpuregs[4][17] ),
    .Y(_00808_));
 sky130_fd_sc_hd__inv_2 _24555_ (.A(\cpuregs[5][17] ),
    .Y(_00809_));
 sky130_fd_sc_hd__inv_2 _24556_ (.A(\cpuregs[6][17] ),
    .Y(_00810_));
 sky130_fd_sc_hd__inv_2 _24557_ (.A(\cpuregs[7][17] ),
    .Y(_00811_));
 sky130_fd_sc_hd__inv_2 _24558_ (.A(\cpuregs[8][17] ),
    .Y(_00813_));
 sky130_fd_sc_hd__inv_2 _24559_ (.A(\cpuregs[9][17] ),
    .Y(_00814_));
 sky130_fd_sc_hd__inv_2 _24560_ (.A(\cpuregs[10][17] ),
    .Y(_00815_));
 sky130_fd_sc_hd__inv_2 _24561_ (.A(\cpuregs[11][17] ),
    .Y(_00816_));
 sky130_fd_sc_hd__inv_2 _24562_ (.A(\cpuregs[12][17] ),
    .Y(_00818_));
 sky130_fd_sc_hd__inv_2 _24563_ (.A(\cpuregs[13][17] ),
    .Y(_00819_));
 sky130_fd_sc_hd__inv_2 _24564_ (.A(\cpuregs[14][17] ),
    .Y(_00820_));
 sky130_fd_sc_hd__inv_2 _24565_ (.A(\cpuregs[15][17] ),
    .Y(_00821_));
 sky130_fd_sc_hd__inv_2 _24566_ (.A(\cpuregs[16][17] ),
    .Y(_00824_));
 sky130_fd_sc_hd__inv_2 _24567_ (.A(\cpuregs[17][17] ),
    .Y(_00825_));
 sky130_fd_sc_hd__inv_2 _24568_ (.A(\cpuregs[18][17] ),
    .Y(_00826_));
 sky130_fd_sc_hd__inv_2 _24569_ (.A(\cpuregs[19][17] ),
    .Y(_00827_));
 sky130_fd_sc_hd__inv_2 _24570_ (.A(\cpuregs[0][18] ),
    .Y(_00830_));
 sky130_fd_sc_hd__inv_2 _24571_ (.A(\cpuregs[1][18] ),
    .Y(_00831_));
 sky130_fd_sc_hd__inv_2 _24572_ (.A(\cpuregs[2][18] ),
    .Y(_00832_));
 sky130_fd_sc_hd__inv_2 _24573_ (.A(\cpuregs[3][18] ),
    .Y(_00833_));
 sky130_fd_sc_hd__inv_2 _24574_ (.A(\cpuregs[4][18] ),
    .Y(_00835_));
 sky130_fd_sc_hd__inv_2 _24575_ (.A(\cpuregs[5][18] ),
    .Y(_00836_));
 sky130_fd_sc_hd__inv_2 _24576_ (.A(\cpuregs[6][18] ),
    .Y(_00837_));
 sky130_fd_sc_hd__inv_2 _24577_ (.A(\cpuregs[7][18] ),
    .Y(_00838_));
 sky130_fd_sc_hd__inv_2 _24578_ (.A(\cpuregs[8][18] ),
    .Y(_00840_));
 sky130_fd_sc_hd__inv_2 _24579_ (.A(\cpuregs[9][18] ),
    .Y(_00841_));
 sky130_fd_sc_hd__inv_2 _24580_ (.A(\cpuregs[10][18] ),
    .Y(_00842_));
 sky130_fd_sc_hd__inv_2 _24581_ (.A(\cpuregs[11][18] ),
    .Y(_00843_));
 sky130_fd_sc_hd__inv_2 _24582_ (.A(\cpuregs[12][18] ),
    .Y(_00845_));
 sky130_fd_sc_hd__inv_2 _24583_ (.A(\cpuregs[13][18] ),
    .Y(_00846_));
 sky130_fd_sc_hd__inv_2 _24584_ (.A(\cpuregs[14][18] ),
    .Y(_00847_));
 sky130_fd_sc_hd__inv_2 _24585_ (.A(\cpuregs[15][18] ),
    .Y(_00848_));
 sky130_fd_sc_hd__inv_2 _24586_ (.A(\cpuregs[16][18] ),
    .Y(_00851_));
 sky130_fd_sc_hd__inv_2 _24587_ (.A(\cpuregs[17][18] ),
    .Y(_00852_));
 sky130_fd_sc_hd__inv_2 _24588_ (.A(\cpuregs[18][18] ),
    .Y(_00853_));
 sky130_fd_sc_hd__inv_2 _24589_ (.A(\cpuregs[19][18] ),
    .Y(_00854_));
 sky130_fd_sc_hd__inv_2 _24590_ (.A(\cpuregs[0][19] ),
    .Y(_00857_));
 sky130_fd_sc_hd__inv_2 _24591_ (.A(\cpuregs[1][19] ),
    .Y(_00858_));
 sky130_fd_sc_hd__inv_2 _24592_ (.A(\cpuregs[2][19] ),
    .Y(_00859_));
 sky130_fd_sc_hd__inv_2 _24593_ (.A(\cpuregs[3][19] ),
    .Y(_00860_));
 sky130_fd_sc_hd__inv_2 _24594_ (.A(\cpuregs[4][19] ),
    .Y(_00862_));
 sky130_fd_sc_hd__inv_2 _24595_ (.A(\cpuregs[5][19] ),
    .Y(_00863_));
 sky130_fd_sc_hd__inv_2 _24596_ (.A(\cpuregs[6][19] ),
    .Y(_00864_));
 sky130_fd_sc_hd__inv_2 _24597_ (.A(\cpuregs[7][19] ),
    .Y(_00865_));
 sky130_fd_sc_hd__inv_2 _24598_ (.A(\cpuregs[8][19] ),
    .Y(_00867_));
 sky130_fd_sc_hd__inv_2 _24599_ (.A(\cpuregs[9][19] ),
    .Y(_00868_));
 sky130_fd_sc_hd__inv_2 _24600_ (.A(\cpuregs[10][19] ),
    .Y(_00869_));
 sky130_fd_sc_hd__inv_2 _24601_ (.A(\cpuregs[11][19] ),
    .Y(_00870_));
 sky130_fd_sc_hd__inv_2 _24602_ (.A(\cpuregs[12][19] ),
    .Y(_00872_));
 sky130_fd_sc_hd__inv_2 _24603_ (.A(\cpuregs[13][19] ),
    .Y(_00873_));
 sky130_fd_sc_hd__inv_2 _24604_ (.A(\cpuregs[14][19] ),
    .Y(_00874_));
 sky130_fd_sc_hd__inv_2 _24605_ (.A(\cpuregs[15][19] ),
    .Y(_00875_));
 sky130_fd_sc_hd__inv_2 _24606_ (.A(\cpuregs[16][19] ),
    .Y(_00878_));
 sky130_fd_sc_hd__inv_2 _24607_ (.A(\cpuregs[17][19] ),
    .Y(_00879_));
 sky130_fd_sc_hd__inv_2 _24608_ (.A(\cpuregs[18][19] ),
    .Y(_00880_));
 sky130_fd_sc_hd__inv_2 _24609_ (.A(\cpuregs[19][19] ),
    .Y(_00881_));
 sky130_fd_sc_hd__inv_2 _24610_ (.A(\cpuregs[0][20] ),
    .Y(_00884_));
 sky130_fd_sc_hd__inv_2 _24611_ (.A(\cpuregs[1][20] ),
    .Y(_00885_));
 sky130_fd_sc_hd__inv_2 _24612_ (.A(\cpuregs[2][20] ),
    .Y(_00886_));
 sky130_fd_sc_hd__inv_2 _24613_ (.A(\cpuregs[3][20] ),
    .Y(_00887_));
 sky130_fd_sc_hd__inv_2 _24614_ (.A(\cpuregs[4][20] ),
    .Y(_00889_));
 sky130_fd_sc_hd__inv_2 _24615_ (.A(\cpuregs[5][20] ),
    .Y(_00890_));
 sky130_fd_sc_hd__inv_2 _24616_ (.A(\cpuregs[6][20] ),
    .Y(_00891_));
 sky130_fd_sc_hd__inv_2 _24617_ (.A(\cpuregs[7][20] ),
    .Y(_00892_));
 sky130_fd_sc_hd__inv_2 _24618_ (.A(\cpuregs[8][20] ),
    .Y(_00894_));
 sky130_fd_sc_hd__inv_2 _24619_ (.A(\cpuregs[9][20] ),
    .Y(_00895_));
 sky130_fd_sc_hd__inv_2 _24620_ (.A(\cpuregs[10][20] ),
    .Y(_00896_));
 sky130_fd_sc_hd__inv_2 _24621_ (.A(\cpuregs[11][20] ),
    .Y(_00897_));
 sky130_fd_sc_hd__inv_2 _24622_ (.A(\cpuregs[12][20] ),
    .Y(_00899_));
 sky130_fd_sc_hd__inv_2 _24623_ (.A(\cpuregs[13][20] ),
    .Y(_00900_));
 sky130_fd_sc_hd__inv_2 _24624_ (.A(\cpuregs[14][20] ),
    .Y(_00901_));
 sky130_fd_sc_hd__inv_2 _24625_ (.A(\cpuregs[15][20] ),
    .Y(_00902_));
 sky130_fd_sc_hd__inv_2 _24626_ (.A(\cpuregs[16][20] ),
    .Y(_00905_));
 sky130_fd_sc_hd__inv_2 _24627_ (.A(\cpuregs[17][20] ),
    .Y(_00906_));
 sky130_fd_sc_hd__inv_2 _24628_ (.A(\cpuregs[18][20] ),
    .Y(_00907_));
 sky130_fd_sc_hd__inv_2 _24629_ (.A(\cpuregs[19][20] ),
    .Y(_00908_));
 sky130_fd_sc_hd__inv_2 _24630_ (.A(\cpuregs[0][21] ),
    .Y(_00911_));
 sky130_fd_sc_hd__inv_2 _24631_ (.A(\cpuregs[1][21] ),
    .Y(_00912_));
 sky130_fd_sc_hd__inv_2 _24632_ (.A(\cpuregs[2][21] ),
    .Y(_00913_));
 sky130_fd_sc_hd__inv_2 _24633_ (.A(\cpuregs[3][21] ),
    .Y(_00914_));
 sky130_fd_sc_hd__inv_2 _24634_ (.A(\cpuregs[4][21] ),
    .Y(_00916_));
 sky130_fd_sc_hd__inv_2 _24635_ (.A(\cpuregs[5][21] ),
    .Y(_00917_));
 sky130_fd_sc_hd__inv_2 _24636_ (.A(\cpuregs[6][21] ),
    .Y(_00918_));
 sky130_fd_sc_hd__inv_2 _24637_ (.A(\cpuregs[7][21] ),
    .Y(_00919_));
 sky130_fd_sc_hd__inv_2 _24638_ (.A(\cpuregs[8][21] ),
    .Y(_00921_));
 sky130_fd_sc_hd__inv_2 _24639_ (.A(\cpuregs[9][21] ),
    .Y(_00922_));
 sky130_fd_sc_hd__inv_2 _24640_ (.A(\cpuregs[10][21] ),
    .Y(_00923_));
 sky130_fd_sc_hd__inv_2 _24641_ (.A(\cpuregs[11][21] ),
    .Y(_00924_));
 sky130_fd_sc_hd__inv_2 _24642_ (.A(\cpuregs[12][21] ),
    .Y(_00926_));
 sky130_fd_sc_hd__inv_2 _24643_ (.A(\cpuregs[13][21] ),
    .Y(_00927_));
 sky130_fd_sc_hd__inv_2 _24644_ (.A(\cpuregs[14][21] ),
    .Y(_00928_));
 sky130_fd_sc_hd__inv_2 _24645_ (.A(\cpuregs[15][21] ),
    .Y(_00929_));
 sky130_fd_sc_hd__inv_2 _24646_ (.A(\cpuregs[16][21] ),
    .Y(_00932_));
 sky130_fd_sc_hd__inv_2 _24647_ (.A(\cpuregs[17][21] ),
    .Y(_00933_));
 sky130_fd_sc_hd__inv_2 _24648_ (.A(\cpuregs[18][21] ),
    .Y(_00934_));
 sky130_fd_sc_hd__inv_2 _24649_ (.A(\cpuregs[19][21] ),
    .Y(_00935_));
 sky130_fd_sc_hd__inv_2 _24650_ (.A(\cpuregs[0][22] ),
    .Y(_00938_));
 sky130_fd_sc_hd__inv_2 _24651_ (.A(\cpuregs[1][22] ),
    .Y(_00939_));
 sky130_fd_sc_hd__inv_2 _24652_ (.A(\cpuregs[2][22] ),
    .Y(_00940_));
 sky130_fd_sc_hd__inv_2 _24653_ (.A(\cpuregs[3][22] ),
    .Y(_00941_));
 sky130_fd_sc_hd__inv_2 _24654_ (.A(\cpuregs[4][22] ),
    .Y(_00943_));
 sky130_fd_sc_hd__inv_2 _24655_ (.A(\cpuregs[5][22] ),
    .Y(_00944_));
 sky130_fd_sc_hd__inv_2 _24656_ (.A(\cpuregs[6][22] ),
    .Y(_00945_));
 sky130_fd_sc_hd__inv_2 _24657_ (.A(\cpuregs[7][22] ),
    .Y(_00946_));
 sky130_fd_sc_hd__a32o_2 _24658_ (.A1(instr_sw),
    .A2(\cpu_state[5] ),
    .A3(_20003_),
    .B1(_18449_),
    .B2(instr_lw),
    .X(_20012_));
 sky130_fd_sc_hd__nor2_2 _24659_ (.A(_19803_),
    .B(_20002_),
    .Y(_20013_));
 sky130_fd_sc_hd__a211o_2 _24660_ (.A1(_18448_),
    .A2(_20012_),
    .B1(_19076_),
    .C1(_20013_),
    .X(_00045_));
 sky130_fd_sc_hd__inv_2 _24661_ (.A(\cpuregs[8][22] ),
    .Y(_00948_));
 sky130_fd_sc_hd__inv_2 _24662_ (.A(\cpuregs[9][22] ),
    .Y(_00949_));
 sky130_fd_sc_hd__inv_2 _24663_ (.A(\cpuregs[10][22] ),
    .Y(_00950_));
 sky130_fd_sc_hd__inv_2 _24664_ (.A(\cpuregs[11][22] ),
    .Y(_00951_));
 sky130_fd_sc_hd__inv_2 _24665_ (.A(\cpuregs[12][22] ),
    .Y(_00953_));
 sky130_fd_sc_hd__inv_2 _24666_ (.A(\cpuregs[13][22] ),
    .Y(_00954_));
 sky130_fd_sc_hd__inv_2 _24667_ (.A(\cpuregs[14][22] ),
    .Y(_00955_));
 sky130_fd_sc_hd__inv_2 _24668_ (.A(\cpuregs[15][22] ),
    .Y(_00956_));
 sky130_fd_sc_hd__inv_2 _24669_ (.A(\cpuregs[16][22] ),
    .Y(_00959_));
 sky130_fd_sc_hd__inv_2 _24670_ (.A(\cpuregs[17][22] ),
    .Y(_00960_));
 sky130_fd_sc_hd__inv_2 _24671_ (.A(\cpuregs[18][22] ),
    .Y(_00961_));
 sky130_fd_sc_hd__inv_2 _24672_ (.A(\cpuregs[19][22] ),
    .Y(_00962_));
 sky130_fd_sc_hd__inv_2 _24673_ (.A(\cpuregs[0][23] ),
    .Y(_00965_));
 sky130_fd_sc_hd__inv_2 _24674_ (.A(\cpuregs[1][23] ),
    .Y(_00966_));
 sky130_fd_sc_hd__inv_2 _24675_ (.A(\cpuregs[2][23] ),
    .Y(_00967_));
 sky130_fd_sc_hd__inv_2 _24676_ (.A(\cpuregs[3][23] ),
    .Y(_00968_));
 sky130_fd_sc_hd__inv_2 _24677_ (.A(\cpuregs[4][23] ),
    .Y(_00970_));
 sky130_fd_sc_hd__inv_2 _24678_ (.A(\cpuregs[5][23] ),
    .Y(_00971_));
 sky130_fd_sc_hd__inv_2 _24679_ (.A(\cpuregs[6][23] ),
    .Y(_00972_));
 sky130_fd_sc_hd__inv_2 _24680_ (.A(\cpuregs[7][23] ),
    .Y(_00973_));
 sky130_fd_sc_hd__inv_2 _24681_ (.A(\cpuregs[8][23] ),
    .Y(_00975_));
 sky130_fd_sc_hd__inv_2 _24682_ (.A(\cpuregs[9][23] ),
    .Y(_00976_));
 sky130_fd_sc_hd__inv_2 _24683_ (.A(\cpuregs[10][23] ),
    .Y(_00977_));
 sky130_fd_sc_hd__inv_2 _24684_ (.A(\cpuregs[11][23] ),
    .Y(_00978_));
 sky130_fd_sc_hd__inv_2 _24685_ (.A(\cpuregs[12][23] ),
    .Y(_00980_));
 sky130_fd_sc_hd__inv_2 _24686_ (.A(\cpuregs[13][23] ),
    .Y(_00981_));
 sky130_fd_sc_hd__inv_2 _24687_ (.A(\cpuregs[14][23] ),
    .Y(_00982_));
 sky130_fd_sc_hd__inv_2 _24688_ (.A(\cpuregs[15][23] ),
    .Y(_00983_));
 sky130_fd_sc_hd__inv_2 _24689_ (.A(\cpuregs[16][23] ),
    .Y(_00986_));
 sky130_fd_sc_hd__inv_2 _24690_ (.A(\cpuregs[17][23] ),
    .Y(_00987_));
 sky130_fd_sc_hd__inv_2 _24691_ (.A(\cpuregs[18][23] ),
    .Y(_00988_));
 sky130_fd_sc_hd__inv_2 _24692_ (.A(\cpuregs[19][23] ),
    .Y(_00989_));
 sky130_fd_sc_hd__inv_2 _24693_ (.A(\cpuregs[0][24] ),
    .Y(_00992_));
 sky130_fd_sc_hd__inv_2 _24694_ (.A(\cpuregs[1][24] ),
    .Y(_00993_));
 sky130_fd_sc_hd__inv_2 _24695_ (.A(\cpuregs[2][24] ),
    .Y(_00994_));
 sky130_fd_sc_hd__inv_2 _24696_ (.A(\cpuregs[3][24] ),
    .Y(_00995_));
 sky130_fd_sc_hd__inv_2 _24697_ (.A(\cpuregs[4][24] ),
    .Y(_00997_));
 sky130_fd_sc_hd__inv_2 _24698_ (.A(\cpuregs[5][24] ),
    .Y(_00998_));
 sky130_fd_sc_hd__inv_2 _24699_ (.A(\cpuregs[6][24] ),
    .Y(_00999_));
 sky130_fd_sc_hd__inv_2 _24700_ (.A(\cpuregs[7][24] ),
    .Y(_01000_));
 sky130_fd_sc_hd__inv_2 _24701_ (.A(\cpuregs[8][24] ),
    .Y(_01002_));
 sky130_fd_sc_hd__inv_2 _24702_ (.A(\cpuregs[9][24] ),
    .Y(_01003_));
 sky130_fd_sc_hd__inv_2 _24703_ (.A(\cpuregs[10][24] ),
    .Y(_01004_));
 sky130_fd_sc_hd__inv_2 _24704_ (.A(\cpuregs[11][24] ),
    .Y(_01005_));
 sky130_fd_sc_hd__inv_2 _24705_ (.A(\cpuregs[12][24] ),
    .Y(_01007_));
 sky130_fd_sc_hd__inv_2 _24706_ (.A(\cpuregs[13][24] ),
    .Y(_01008_));
 sky130_fd_sc_hd__inv_2 _24707_ (.A(\cpuregs[14][24] ),
    .Y(_01009_));
 sky130_fd_sc_hd__inv_2 _24708_ (.A(\cpuregs[15][24] ),
    .Y(_01010_));
 sky130_fd_sc_hd__inv_2 _24709_ (.A(\cpuregs[16][24] ),
    .Y(_01013_));
 sky130_fd_sc_hd__inv_2 _24710_ (.A(\cpuregs[17][24] ),
    .Y(_01014_));
 sky130_fd_sc_hd__inv_2 _24711_ (.A(\cpuregs[18][24] ),
    .Y(_01015_));
 sky130_fd_sc_hd__inv_2 _24712_ (.A(\cpuregs[19][24] ),
    .Y(_01016_));
 sky130_fd_sc_hd__inv_2 _24713_ (.A(\cpuregs[0][25] ),
    .Y(_01019_));
 sky130_fd_sc_hd__inv_2 _24714_ (.A(\cpuregs[1][25] ),
    .Y(_01020_));
 sky130_fd_sc_hd__inv_2 _24715_ (.A(\cpuregs[2][25] ),
    .Y(_01021_));
 sky130_fd_sc_hd__inv_2 _24716_ (.A(\cpuregs[3][25] ),
    .Y(_01022_));
 sky130_fd_sc_hd__inv_2 _24717_ (.A(\cpuregs[4][25] ),
    .Y(_01024_));
 sky130_fd_sc_hd__inv_2 _24718_ (.A(\cpuregs[5][25] ),
    .Y(_01025_));
 sky130_fd_sc_hd__inv_2 _24719_ (.A(\cpuregs[6][25] ),
    .Y(_01026_));
 sky130_fd_sc_hd__inv_2 _24720_ (.A(\cpuregs[7][25] ),
    .Y(_01027_));
 sky130_fd_sc_hd__nor2_2 _24721_ (.A(\mem_state[1] ),
    .B(_18039_),
    .Y(_00289_));
 sky130_fd_sc_hd__nand2_2 _24722_ (.A(_18053_),
    .B(_00289_),
    .Y(_00298_));
 sky130_fd_sc_hd__inv_2 _24723_ (.A(\cpuregs[8][25] ),
    .Y(_01029_));
 sky130_fd_sc_hd__inv_2 _24724_ (.A(\cpuregs[9][25] ),
    .Y(_01030_));
 sky130_fd_sc_hd__inv_2 _24725_ (.A(\cpuregs[10][25] ),
    .Y(_01031_));
 sky130_fd_sc_hd__inv_2 _24726_ (.A(\cpuregs[11][25] ),
    .Y(_01032_));
 sky130_fd_sc_hd__inv_2 _24727_ (.A(\cpuregs[12][25] ),
    .Y(_01034_));
 sky130_fd_sc_hd__inv_2 _24728_ (.A(\cpuregs[13][25] ),
    .Y(_01035_));
 sky130_fd_sc_hd__inv_2 _24729_ (.A(\cpuregs[14][25] ),
    .Y(_01036_));
 sky130_fd_sc_hd__inv_2 _24730_ (.A(\cpuregs[15][25] ),
    .Y(_01037_));
 sky130_fd_sc_hd__inv_2 _24731_ (.A(\cpuregs[16][25] ),
    .Y(_01040_));
 sky130_fd_sc_hd__inv_2 _24732_ (.A(\cpuregs[17][25] ),
    .Y(_01041_));
 sky130_fd_sc_hd__inv_2 _24733_ (.A(\cpuregs[18][25] ),
    .Y(_01042_));
 sky130_fd_sc_hd__inv_2 _24734_ (.A(\cpuregs[19][25] ),
    .Y(_01043_));
 sky130_fd_sc_hd__inv_2 _24735_ (.A(\cpuregs[0][26] ),
    .Y(_01046_));
 sky130_fd_sc_hd__inv_2 _24736_ (.A(\cpuregs[1][26] ),
    .Y(_01047_));
 sky130_fd_sc_hd__inv_2 _24737_ (.A(\cpuregs[2][26] ),
    .Y(_01048_));
 sky130_fd_sc_hd__inv_2 _24738_ (.A(\cpuregs[3][26] ),
    .Y(_01049_));
 sky130_fd_sc_hd__inv_2 _24739_ (.A(\cpuregs[4][26] ),
    .Y(_01051_));
 sky130_fd_sc_hd__inv_2 _24740_ (.A(\cpuregs[5][26] ),
    .Y(_01052_));
 sky130_fd_sc_hd__inv_2 _24741_ (.A(\cpuregs[6][26] ),
    .Y(_01053_));
 sky130_fd_sc_hd__inv_2 _24742_ (.A(\cpuregs[7][26] ),
    .Y(_01054_));
 sky130_fd_sc_hd__inv_2 _24743_ (.A(\cpuregs[8][26] ),
    .Y(_01056_));
 sky130_fd_sc_hd__inv_2 _24744_ (.A(\cpuregs[9][26] ),
    .Y(_01057_));
 sky130_fd_sc_hd__inv_2 _24745_ (.A(\cpuregs[10][26] ),
    .Y(_01058_));
 sky130_fd_sc_hd__inv_2 _24746_ (.A(\cpuregs[11][26] ),
    .Y(_01059_));
 sky130_fd_sc_hd__inv_2 _24747_ (.A(\cpuregs[12][26] ),
    .Y(_01061_));
 sky130_fd_sc_hd__inv_2 _24748_ (.A(\cpuregs[13][26] ),
    .Y(_01062_));
 sky130_fd_sc_hd__inv_2 _24749_ (.A(\cpuregs[14][26] ),
    .Y(_01063_));
 sky130_fd_sc_hd__inv_2 _24750_ (.A(\cpuregs[15][26] ),
    .Y(_01064_));
 sky130_fd_sc_hd__inv_2 _24751_ (.A(\cpuregs[16][26] ),
    .Y(_01067_));
 sky130_fd_sc_hd__inv_2 _24752_ (.A(\cpuregs[17][26] ),
    .Y(_01068_));
 sky130_fd_sc_hd__inv_2 _24753_ (.A(\cpuregs[18][26] ),
    .Y(_01069_));
 sky130_fd_sc_hd__inv_2 _24754_ (.A(\cpuregs[19][26] ),
    .Y(_01070_));
 sky130_fd_sc_hd__inv_2 _24755_ (.A(\mem_wordsize[1] ),
    .Y(_20014_));
 sky130_fd_sc_hd__buf_1 _24756_ (.A(_20014_),
    .X(_20015_));
 sky130_fd_sc_hd__buf_1 _24757_ (.A(_18019_),
    .X(_20016_));
 sky130_fd_sc_hd__o211a_2 _24758_ (.A1(instr_lbu),
    .A2(instr_lb),
    .B1(_18029_),
    .C1(_20016_),
    .X(_20017_));
 sky130_fd_sc_hd__a31o_2 _24759_ (.A1(_00291_),
    .A2(instr_sb),
    .A3(\cpu_state[5] ),
    .B1(_20017_),
    .X(_20018_));
 sky130_fd_sc_hd__a2bb2o_2 _24760_ (.A1_N(_20015_),
    .A2_N(_20002_),
    .B1(_18018_),
    .B2(_20018_),
    .X(_00046_));
 sky130_fd_sc_hd__inv_2 _24761_ (.A(\cpuregs[0][27] ),
    .Y(_01073_));
 sky130_fd_sc_hd__inv_2 _24762_ (.A(\cpuregs[1][27] ),
    .Y(_01074_));
 sky130_fd_sc_hd__inv_2 _24763_ (.A(\cpuregs[2][27] ),
    .Y(_01075_));
 sky130_fd_sc_hd__inv_2 _24764_ (.A(\cpuregs[3][27] ),
    .Y(_01076_));
 sky130_fd_sc_hd__inv_2 _24765_ (.A(\cpuregs[4][27] ),
    .Y(_01078_));
 sky130_fd_sc_hd__inv_2 _24766_ (.A(\cpuregs[5][27] ),
    .Y(_01079_));
 sky130_fd_sc_hd__inv_2 _24767_ (.A(\cpuregs[6][27] ),
    .Y(_01080_));
 sky130_fd_sc_hd__inv_2 _24768_ (.A(\cpuregs[7][27] ),
    .Y(_01081_));
 sky130_fd_sc_hd__inv_2 _24769_ (.A(\cpuregs[8][27] ),
    .Y(_01083_));
 sky130_fd_sc_hd__inv_2 _24770_ (.A(\cpuregs[9][27] ),
    .Y(_01084_));
 sky130_fd_sc_hd__inv_2 _24771_ (.A(\cpuregs[10][27] ),
    .Y(_01085_));
 sky130_fd_sc_hd__inv_2 _24772_ (.A(\cpuregs[11][27] ),
    .Y(_01086_));
 sky130_fd_sc_hd__inv_2 _24773_ (.A(\cpuregs[12][27] ),
    .Y(_01088_));
 sky130_fd_sc_hd__inv_2 _24774_ (.A(\cpuregs[13][27] ),
    .Y(_01089_));
 sky130_fd_sc_hd__inv_2 _24775_ (.A(\cpuregs[14][27] ),
    .Y(_01090_));
 sky130_fd_sc_hd__inv_2 _24776_ (.A(\cpuregs[15][27] ),
    .Y(_01091_));
 sky130_fd_sc_hd__inv_2 _24777_ (.A(\cpuregs[16][27] ),
    .Y(_01094_));
 sky130_fd_sc_hd__inv_2 _24778_ (.A(\cpuregs[17][27] ),
    .Y(_01095_));
 sky130_fd_sc_hd__inv_2 _24779_ (.A(\cpuregs[18][27] ),
    .Y(_01096_));
 sky130_fd_sc_hd__inv_2 _24780_ (.A(\cpuregs[19][27] ),
    .Y(_01097_));
 sky130_fd_sc_hd__inv_2 _24781_ (.A(\cpuregs[0][28] ),
    .Y(_01100_));
 sky130_fd_sc_hd__inv_2 _24782_ (.A(\cpuregs[1][28] ),
    .Y(_01101_));
 sky130_fd_sc_hd__inv_2 _24783_ (.A(\cpuregs[2][28] ),
    .Y(_01102_));
 sky130_fd_sc_hd__inv_2 _24784_ (.A(\cpuregs[3][28] ),
    .Y(_01103_));
 sky130_fd_sc_hd__inv_2 _24785_ (.A(\cpuregs[4][28] ),
    .Y(_01105_));
 sky130_fd_sc_hd__inv_2 _24786_ (.A(\cpuregs[5][28] ),
    .Y(_01106_));
 sky130_fd_sc_hd__inv_2 _24787_ (.A(\cpuregs[6][28] ),
    .Y(_01107_));
 sky130_fd_sc_hd__inv_2 _24788_ (.A(\cpuregs[7][28] ),
    .Y(_01108_));
 sky130_fd_sc_hd__inv_2 _24789_ (.A(\cpuregs[8][28] ),
    .Y(_01110_));
 sky130_fd_sc_hd__inv_2 _24790_ (.A(\cpuregs[9][28] ),
    .Y(_01111_));
 sky130_fd_sc_hd__inv_2 _24791_ (.A(\cpuregs[10][28] ),
    .Y(_01112_));
 sky130_fd_sc_hd__inv_2 _24792_ (.A(\cpuregs[11][28] ),
    .Y(_01113_));
 sky130_fd_sc_hd__inv_2 _24793_ (.A(\cpuregs[12][28] ),
    .Y(_01115_));
 sky130_fd_sc_hd__inv_2 _24794_ (.A(\cpuregs[13][28] ),
    .Y(_01116_));
 sky130_fd_sc_hd__inv_2 _24795_ (.A(\cpuregs[14][28] ),
    .Y(_01117_));
 sky130_fd_sc_hd__inv_2 _24796_ (.A(\cpuregs[15][28] ),
    .Y(_01118_));
 sky130_fd_sc_hd__inv_2 _24797_ (.A(\cpuregs[16][28] ),
    .Y(_01121_));
 sky130_fd_sc_hd__inv_2 _24798_ (.A(\cpuregs[17][28] ),
    .Y(_01122_));
 sky130_fd_sc_hd__inv_2 _24799_ (.A(\cpuregs[18][28] ),
    .Y(_01123_));
 sky130_fd_sc_hd__inv_2 _24800_ (.A(\cpuregs[19][28] ),
    .Y(_01124_));
 sky130_fd_sc_hd__inv_2 _24801_ (.A(\cpuregs[0][29] ),
    .Y(_01127_));
 sky130_fd_sc_hd__inv_2 _24802_ (.A(\cpuregs[1][29] ),
    .Y(_01128_));
 sky130_fd_sc_hd__inv_2 _24803_ (.A(\cpuregs[2][29] ),
    .Y(_01129_));
 sky130_fd_sc_hd__inv_2 _24804_ (.A(\cpuregs[3][29] ),
    .Y(_01130_));
 sky130_fd_sc_hd__inv_2 _24805_ (.A(\cpuregs[4][29] ),
    .Y(_01132_));
 sky130_fd_sc_hd__inv_2 _24806_ (.A(\cpuregs[5][29] ),
    .Y(_01133_));
 sky130_fd_sc_hd__inv_2 _24807_ (.A(\cpuregs[6][29] ),
    .Y(_01134_));
 sky130_fd_sc_hd__inv_2 _24808_ (.A(\cpuregs[7][29] ),
    .Y(_01135_));
 sky130_fd_sc_hd__inv_2 _24809_ (.A(\cpuregs[8][29] ),
    .Y(_01137_));
 sky130_fd_sc_hd__inv_2 _24810_ (.A(\cpuregs[9][29] ),
    .Y(_01138_));
 sky130_fd_sc_hd__inv_2 _24811_ (.A(\cpuregs[10][29] ),
    .Y(_01139_));
 sky130_fd_sc_hd__inv_2 _24812_ (.A(\cpuregs[11][29] ),
    .Y(_01140_));
 sky130_fd_sc_hd__inv_2 _24813_ (.A(\cpuregs[12][29] ),
    .Y(_01142_));
 sky130_fd_sc_hd__inv_2 _24814_ (.A(\cpuregs[13][29] ),
    .Y(_01143_));
 sky130_fd_sc_hd__buf_1 _24815_ (.A(latched_branch),
    .X(_20019_));
 sky130_fd_sc_hd__buf_1 _24816_ (.A(_20019_),
    .X(_20020_));
 sky130_fd_sc_hd__and2_2 _24817_ (.A(_20020_),
    .B(_00294_),
    .X(_00295_));
 sky130_fd_sc_hd__inv_2 _24818_ (.A(\cpuregs[14][29] ),
    .Y(_01144_));
 sky130_fd_sc_hd__inv_2 _24819_ (.A(\cpuregs[15][29] ),
    .Y(_01145_));
 sky130_fd_sc_hd__inv_2 _24820_ (.A(\cpuregs[16][29] ),
    .Y(_01148_));
 sky130_fd_sc_hd__inv_2 _24821_ (.A(\cpuregs[17][29] ),
    .Y(_01149_));
 sky130_fd_sc_hd__inv_2 _24822_ (.A(\cpuregs[18][29] ),
    .Y(_01150_));
 sky130_fd_sc_hd__inv_2 _24823_ (.A(\cpuregs[19][29] ),
    .Y(_01151_));
 sky130_fd_sc_hd__inv_2 _24824_ (.A(\cpuregs[0][30] ),
    .Y(_01154_));
 sky130_fd_sc_hd__inv_2 _24825_ (.A(\cpuregs[1][30] ),
    .Y(_01155_));
 sky130_fd_sc_hd__inv_2 _24826_ (.A(\cpuregs[2][30] ),
    .Y(_01156_));
 sky130_fd_sc_hd__inv_2 _24827_ (.A(\cpuregs[3][30] ),
    .Y(_01157_));
 sky130_fd_sc_hd__inv_2 _24828_ (.A(\cpuregs[4][30] ),
    .Y(_01159_));
 sky130_fd_sc_hd__inv_2 _24829_ (.A(\cpuregs[5][30] ),
    .Y(_01160_));
 sky130_fd_sc_hd__inv_2 _24830_ (.A(\cpuregs[6][30] ),
    .Y(_01161_));
 sky130_fd_sc_hd__inv_2 _24831_ (.A(\cpuregs[7][30] ),
    .Y(_01162_));
 sky130_fd_sc_hd__inv_2 _24832_ (.A(\cpuregs[8][30] ),
    .Y(_01164_));
 sky130_fd_sc_hd__inv_2 _24833_ (.A(\cpuregs[9][30] ),
    .Y(_01165_));
 sky130_fd_sc_hd__inv_2 _24834_ (.A(\cpuregs[10][30] ),
    .Y(_01166_));
 sky130_fd_sc_hd__inv_2 _24835_ (.A(\cpuregs[11][30] ),
    .Y(_01167_));
 sky130_fd_sc_hd__inv_2 _24836_ (.A(\cpuregs[12][30] ),
    .Y(_01169_));
 sky130_fd_sc_hd__inv_2 _24837_ (.A(\cpuregs[13][30] ),
    .Y(_01170_));
 sky130_fd_sc_hd__inv_2 _24838_ (.A(\cpuregs[14][30] ),
    .Y(_01171_));
 sky130_fd_sc_hd__inv_2 _24839_ (.A(\cpuregs[15][30] ),
    .Y(_01172_));
 sky130_fd_sc_hd__inv_2 _24840_ (.A(\cpuregs[16][30] ),
    .Y(_01175_));
 sky130_fd_sc_hd__inv_2 _24841_ (.A(\cpuregs[17][30] ),
    .Y(_01176_));
 sky130_fd_sc_hd__inv_2 _24842_ (.A(\cpuregs[18][30] ),
    .Y(_01177_));
 sky130_fd_sc_hd__inv_2 _24843_ (.A(\cpuregs[19][30] ),
    .Y(_01178_));
 sky130_fd_sc_hd__inv_2 _24844_ (.A(\cpuregs[0][31] ),
    .Y(_01181_));
 sky130_fd_sc_hd__inv_2 _24845_ (.A(\cpuregs[1][31] ),
    .Y(_01182_));
 sky130_fd_sc_hd__inv_2 _24846_ (.A(\cpuregs[2][31] ),
    .Y(_01183_));
 sky130_fd_sc_hd__inv_2 _24847_ (.A(\cpuregs[3][31] ),
    .Y(_01184_));
 sky130_fd_sc_hd__inv_2 _24848_ (.A(\cpuregs[4][31] ),
    .Y(_01186_));
 sky130_fd_sc_hd__inv_2 _24849_ (.A(\cpuregs[5][31] ),
    .Y(_01187_));
 sky130_fd_sc_hd__inv_2 _24850_ (.A(\cpuregs[6][31] ),
    .Y(_01188_));
 sky130_fd_sc_hd__inv_2 _24851_ (.A(\cpuregs[7][31] ),
    .Y(_01189_));
 sky130_fd_sc_hd__inv_2 _24852_ (.A(\cpuregs[8][31] ),
    .Y(_01191_));
 sky130_fd_sc_hd__inv_2 _24853_ (.A(\cpuregs[9][31] ),
    .Y(_01192_));
 sky130_fd_sc_hd__inv_2 _24854_ (.A(\cpuregs[10][31] ),
    .Y(_01193_));
 sky130_fd_sc_hd__inv_2 _24855_ (.A(\cpuregs[11][31] ),
    .Y(_01194_));
 sky130_fd_sc_hd__inv_2 _24856_ (.A(\cpuregs[12][31] ),
    .Y(_01196_));
 sky130_fd_sc_hd__inv_2 _24857_ (.A(\cpuregs[13][31] ),
    .Y(_01197_));
 sky130_fd_sc_hd__inv_2 _24858_ (.A(\cpuregs[14][31] ),
    .Y(_01198_));
 sky130_fd_sc_hd__inv_2 _24859_ (.A(\cpuregs[15][31] ),
    .Y(_01199_));
 sky130_fd_sc_hd__inv_2 _24860_ (.A(\cpuregs[16][31] ),
    .Y(_01202_));
 sky130_fd_sc_hd__inv_2 _24861_ (.A(\cpuregs[17][31] ),
    .Y(_01203_));
 sky130_fd_sc_hd__inv_2 _24862_ (.A(\cpuregs[18][31] ),
    .Y(_01204_));
 sky130_fd_sc_hd__inv_2 _24863_ (.A(\cpuregs[19][31] ),
    .Y(_01205_));
 sky130_fd_sc_hd__or4_2 _24864_ (.A(\timer[21] ),
    .B(\timer[20] ),
    .C(\timer[23] ),
    .D(\timer[22] ),
    .X(_20021_));
 sky130_fd_sc_hd__nor2_2 _24865_ (.A(\timer[5] ),
    .B(\timer[4] ),
    .Y(_20022_));
 sky130_fd_sc_hd__inv_2 _24866_ (.A(_20022_),
    .Y(_20023_));
 sky130_fd_sc_hd__or2_2 _24867_ (.A(\timer[1] ),
    .B(\timer[0] ),
    .X(_20024_));
 sky130_fd_sc_hd__nor2_2 _24868_ (.A(\timer[2] ),
    .B(_20024_),
    .Y(_20025_));
 sky130_fd_sc_hd__inv_2 _24869_ (.A(\timer[3] ),
    .Y(_20026_));
 sky130_fd_sc_hd__nand2_2 _24870_ (.A(_20025_),
    .B(_20026_),
    .Y(_20027_));
 sky130_fd_sc_hd__nor2_2 _24871_ (.A(_20023_),
    .B(_20027_),
    .Y(_20028_));
 sky130_fd_sc_hd__inv_2 _24872_ (.A(_20028_),
    .Y(_20029_));
 sky130_fd_sc_hd__nor2_2 _24873_ (.A(\timer[6] ),
    .B(_20029_),
    .Y(_20030_));
 sky130_fd_sc_hd__inv_2 _24874_ (.A(_20030_),
    .Y(_20031_));
 sky130_fd_sc_hd__nor2_2 _24875_ (.A(\timer[7] ),
    .B(_20031_),
    .Y(_20032_));
 sky130_fd_sc_hd__nor2_2 _24876_ (.A(\timer[9] ),
    .B(\timer[8] ),
    .Y(_20033_));
 sky130_fd_sc_hd__nand2_2 _24877_ (.A(_20032_),
    .B(_20033_),
    .Y(_20034_));
 sky130_fd_sc_hd__or2_2 _24878_ (.A(\timer[10] ),
    .B(_20034_),
    .X(_20035_));
 sky130_fd_sc_hd__or2_2 _24879_ (.A(\timer[11] ),
    .B(_20035_),
    .X(_20036_));
 sky130_fd_sc_hd__or2_2 _24880_ (.A(\timer[12] ),
    .B(_20036_),
    .X(_20037_));
 sky130_fd_sc_hd__nor2_2 _24881_ (.A(\timer[13] ),
    .B(_20037_),
    .Y(_20038_));
 sky130_fd_sc_hd__inv_2 _24882_ (.A(\timer[14] ),
    .Y(_20039_));
 sky130_fd_sc_hd__nand2_2 _24883_ (.A(_20038_),
    .B(_20039_),
    .Y(_20040_));
 sky130_fd_sc_hd__nor2_2 _24884_ (.A(\timer[15] ),
    .B(_20040_),
    .Y(_20041_));
 sky130_fd_sc_hd__nor2_2 _24885_ (.A(\timer[17] ),
    .B(\timer[16] ),
    .Y(_20042_));
 sky130_fd_sc_hd__inv_2 _24886_ (.A(\timer[19] ),
    .Y(_20043_));
 sky130_fd_sc_hd__inv_2 _24887_ (.A(\timer[18] ),
    .Y(_20044_));
 sky130_fd_sc_hd__and3_2 _24888_ (.A(_20042_),
    .B(_20043_),
    .C(_20044_),
    .X(_20045_));
 sky130_fd_sc_hd__nand2_2 _24889_ (.A(_20041_),
    .B(_20045_),
    .Y(_20046_));
 sky130_fd_sc_hd__nor2_2 _24890_ (.A(_20021_),
    .B(_20046_),
    .Y(_20047_));
 sky130_fd_sc_hd__nor2_2 _24891_ (.A(\timer[25] ),
    .B(\timer[24] ),
    .Y(_20048_));
 sky130_fd_sc_hd__nand2_2 _24892_ (.A(_20047_),
    .B(_20048_),
    .Y(_20049_));
 sky130_fd_sc_hd__or2_2 _24893_ (.A(\timer[26] ),
    .B(_20049_),
    .X(_20050_));
 sky130_fd_sc_hd__nor2_2 _24894_ (.A(\timer[27] ),
    .B(_20050_),
    .Y(_20051_));
 sky130_fd_sc_hd__nor2_2 _24895_ (.A(\timer[29] ),
    .B(\timer[28] ),
    .Y(_20052_));
 sky130_fd_sc_hd__nand2_2 _24896_ (.A(_20051_),
    .B(_20052_),
    .Y(_20053_));
 sky130_fd_sc_hd__or2_2 _24897_ (.A(\timer[30] ),
    .B(_20053_),
    .X(_20054_));
 sky130_fd_sc_hd__nor2_2 _24898_ (.A(\timer[31] ),
    .B(_20054_),
    .Y(_01208_));
 sky130_fd_sc_hd__nor2_2 _24899_ (.A(\timer[0] ),
    .B(_01208_),
    .Y(_01209_));
 sky130_fd_sc_hd__nand2_2 _24900_ (.A(\timer[1] ),
    .B(\timer[0] ),
    .Y(_20055_));
 sky130_fd_sc_hd__nand2_2 _24901_ (.A(_20024_),
    .B(_20055_),
    .Y(_01211_));
 sky130_fd_sc_hd__and2_2 _24902_ (.A(_20024_),
    .B(\timer[2] ),
    .X(_20056_));
 sky130_fd_sc_hd__or2_2 _24903_ (.A(_20025_),
    .B(_20056_),
    .X(_01214_));
 sky130_fd_sc_hd__or2_2 _24904_ (.A(_20026_),
    .B(_20025_),
    .X(_20057_));
 sky130_fd_sc_hd__nand2_2 _24905_ (.A(_20057_),
    .B(_20027_),
    .Y(_01217_));
 sky130_fd_sc_hd__or2_2 _24906_ (.A(\timer[4] ),
    .B(_20027_),
    .X(_20058_));
 sky130_fd_sc_hd__nand2_2 _24907_ (.A(_20027_),
    .B(\timer[4] ),
    .Y(_20059_));
 sky130_fd_sc_hd__nand2_2 _24908_ (.A(_20058_),
    .B(_20059_),
    .Y(_01220_));
 sky130_fd_sc_hd__a21o_2 _24909_ (.A1(_20058_),
    .A2(\timer[5] ),
    .B1(_20028_),
    .X(_01223_));
 sky130_fd_sc_hd__nand2_2 _24910_ (.A(_20029_),
    .B(\timer[6] ),
    .Y(_20060_));
 sky130_fd_sc_hd__nand2_2 _24911_ (.A(_20031_),
    .B(_20060_),
    .Y(_01226_));
 sky130_fd_sc_hd__inv_2 _24912_ (.A(\timer[7] ),
    .Y(_20061_));
 sky130_fd_sc_hd__nor2_2 _24913_ (.A(_20061_),
    .B(_20030_),
    .Y(_20062_));
 sky130_fd_sc_hd__or2_2 _24914_ (.A(_20062_),
    .B(_20032_),
    .X(_01229_));
 sky130_fd_sc_hd__inv_2 _24915_ (.A(\timer[8] ),
    .Y(_20063_));
 sky130_fd_sc_hd__or2_2 _24916_ (.A(_20063_),
    .B(_20032_),
    .X(_20064_));
 sky130_fd_sc_hd__nand2_2 _24917_ (.A(_20032_),
    .B(_20063_),
    .Y(_20065_));
 sky130_fd_sc_hd__nand2_2 _24918_ (.A(_20064_),
    .B(_20065_),
    .Y(_01232_));
 sky130_fd_sc_hd__nand2_2 _24919_ (.A(_20065_),
    .B(\timer[9] ),
    .Y(_20066_));
 sky130_fd_sc_hd__nand2_2 _24920_ (.A(_20066_),
    .B(_20034_),
    .Y(_01235_));
 sky130_fd_sc_hd__nand2_2 _24921_ (.A(_20034_),
    .B(\timer[10] ),
    .Y(_20067_));
 sky130_fd_sc_hd__nand2_2 _24922_ (.A(_20035_),
    .B(_20067_),
    .Y(_01238_));
 sky130_fd_sc_hd__nand2_2 _24923_ (.A(_20035_),
    .B(\timer[11] ),
    .Y(_20068_));
 sky130_fd_sc_hd__nand2_2 _24924_ (.A(_20036_),
    .B(_20068_),
    .Y(_01241_));
 sky130_fd_sc_hd__nand2_2 _24925_ (.A(_20036_),
    .B(\timer[12] ),
    .Y(_20069_));
 sky130_fd_sc_hd__nand2_2 _24926_ (.A(_20037_),
    .B(_20069_),
    .Y(_01244_));
 sky130_fd_sc_hd__and2_2 _24927_ (.A(_20037_),
    .B(\timer[13] ),
    .X(_20070_));
 sky130_fd_sc_hd__or2_2 _24928_ (.A(_20038_),
    .B(_20070_),
    .X(_01247_));
 sky130_fd_sc_hd__or2_2 _24929_ (.A(_20039_),
    .B(_20038_),
    .X(_20071_));
 sky130_fd_sc_hd__nand2_2 _24930_ (.A(_20071_),
    .B(_20040_),
    .Y(_01250_));
 sky130_fd_sc_hd__inv_2 _24931_ (.A(_20041_),
    .Y(_20072_));
 sky130_fd_sc_hd__nand2_2 _24932_ (.A(_20040_),
    .B(\timer[15] ),
    .Y(_20073_));
 sky130_fd_sc_hd__nand2_2 _24933_ (.A(_20072_),
    .B(_20073_),
    .Y(_01253_));
 sky130_fd_sc_hd__nand2_2 _24934_ (.A(_20072_),
    .B(\timer[16] ),
    .Y(_20074_));
 sky130_fd_sc_hd__inv_2 _24935_ (.A(\timer[16] ),
    .Y(_20075_));
 sky130_fd_sc_hd__nand2_2 _24936_ (.A(_20041_),
    .B(_20075_),
    .Y(_20076_));
 sky130_fd_sc_hd__nand2_2 _24937_ (.A(_20074_),
    .B(_20076_),
    .Y(_01256_));
 sky130_fd_sc_hd__nand2_2 _24938_ (.A(_20076_),
    .B(\timer[17] ),
    .Y(_20077_));
 sky130_fd_sc_hd__nand2_2 _24939_ (.A(_20041_),
    .B(_20042_),
    .Y(_20078_));
 sky130_fd_sc_hd__nand2_2 _24940_ (.A(_20077_),
    .B(_20078_),
    .Y(_01259_));
 sky130_fd_sc_hd__or2_2 _24941_ (.A(\timer[18] ),
    .B(_20078_),
    .X(_20079_));
 sky130_fd_sc_hd__nand2_2 _24942_ (.A(_20078_),
    .B(\timer[18] ),
    .Y(_20080_));
 sky130_fd_sc_hd__nand2_2 _24943_ (.A(_20079_),
    .B(_20080_),
    .Y(_01262_));
 sky130_fd_sc_hd__nand2_2 _24944_ (.A(_20079_),
    .B(\timer[19] ),
    .Y(_20081_));
 sky130_fd_sc_hd__nand2_2 _24945_ (.A(_20081_),
    .B(_20046_),
    .Y(_01265_));
 sky130_fd_sc_hd__or2_2 _24946_ (.A(\timer[20] ),
    .B(_20046_),
    .X(_20082_));
 sky130_fd_sc_hd__nand2_2 _24947_ (.A(_20046_),
    .B(\timer[20] ),
    .Y(_20083_));
 sky130_fd_sc_hd__nand2_2 _24948_ (.A(_20082_),
    .B(_20083_),
    .Y(_01268_));
 sky130_fd_sc_hd__or2_2 _24949_ (.A(\timer[21] ),
    .B(_20082_),
    .X(_20084_));
 sky130_fd_sc_hd__nand2_2 _24950_ (.A(_20082_),
    .B(\timer[21] ),
    .Y(_20085_));
 sky130_fd_sc_hd__nand2_2 _24951_ (.A(_20084_),
    .B(_20085_),
    .Y(_01271_));
 sky130_fd_sc_hd__or2_2 _24952_ (.A(\timer[22] ),
    .B(_20084_),
    .X(_20086_));
 sky130_fd_sc_hd__nand2_2 _24953_ (.A(_20084_),
    .B(\timer[22] ),
    .Y(_20087_));
 sky130_fd_sc_hd__nand2_2 _24954_ (.A(_20086_),
    .B(_20087_),
    .Y(_01274_));
 sky130_fd_sc_hd__nand2_2 _24955_ (.A(_20086_),
    .B(\timer[23] ),
    .Y(_20088_));
 sky130_fd_sc_hd__inv_2 _24956_ (.A(_20047_),
    .Y(_20089_));
 sky130_fd_sc_hd__nand2_2 _24957_ (.A(_20088_),
    .B(_20089_),
    .Y(_01277_));
 sky130_fd_sc_hd__nand2_2 _24958_ (.A(_20089_),
    .B(\timer[24] ),
    .Y(_20090_));
 sky130_fd_sc_hd__inv_2 _24959_ (.A(\timer[24] ),
    .Y(_20091_));
 sky130_fd_sc_hd__nand2_2 _24960_ (.A(_20047_),
    .B(_20091_),
    .Y(_20092_));
 sky130_fd_sc_hd__nand2_2 _24961_ (.A(_20090_),
    .B(_20092_),
    .Y(_01280_));
 sky130_fd_sc_hd__nand2_2 _24962_ (.A(_20092_),
    .B(\timer[25] ),
    .Y(_20093_));
 sky130_fd_sc_hd__nand2_2 _24963_ (.A(_20093_),
    .B(_20049_),
    .Y(_01283_));
 sky130_fd_sc_hd__nand2_2 _24964_ (.A(_20049_),
    .B(\timer[26] ),
    .Y(_20094_));
 sky130_fd_sc_hd__nand2_2 _24965_ (.A(_20050_),
    .B(_20094_),
    .Y(_01286_));
 sky130_fd_sc_hd__inv_2 _24966_ (.A(_20051_),
    .Y(_20095_));
 sky130_fd_sc_hd__nand2_2 _24967_ (.A(_20050_),
    .B(\timer[27] ),
    .Y(_20096_));
 sky130_fd_sc_hd__nand2_2 _24968_ (.A(_20095_),
    .B(_20096_),
    .Y(_01289_));
 sky130_fd_sc_hd__nand2_2 _24969_ (.A(_20095_),
    .B(\timer[28] ),
    .Y(_20097_));
 sky130_fd_sc_hd__inv_2 _24970_ (.A(\timer[28] ),
    .Y(_20098_));
 sky130_fd_sc_hd__nand2_2 _24971_ (.A(_20051_),
    .B(_20098_),
    .Y(_20099_));
 sky130_fd_sc_hd__nand2_2 _24972_ (.A(_20097_),
    .B(_20099_),
    .Y(_01292_));
 sky130_fd_sc_hd__nand2_2 _24973_ (.A(_20099_),
    .B(\timer[29] ),
    .Y(_20100_));
 sky130_fd_sc_hd__nand2_2 _24974_ (.A(_20100_),
    .B(_20053_),
    .Y(_01295_));
 sky130_fd_sc_hd__nand2_2 _24975_ (.A(_20053_),
    .B(\timer[30] ),
    .Y(_20101_));
 sky130_fd_sc_hd__nand2_2 _24976_ (.A(_20054_),
    .B(_20101_),
    .Y(_01298_));
 sky130_fd_sc_hd__and2_2 _24977_ (.A(_20054_),
    .B(\timer[31] ),
    .X(_20102_));
 sky130_fd_sc_hd__or2_2 _24978_ (.A(_01208_),
    .B(_20102_),
    .X(_01301_));
 sky130_fd_sc_hd__buf_1 _24979_ (.A(_19422_),
    .X(_20103_));
 sky130_fd_sc_hd__inv_2 _24980_ (.A(\decoded_imm[5] ),
    .Y(_20104_));
 sky130_fd_sc_hd__nor2_2 _24981_ (.A(_20103_),
    .B(_20104_),
    .Y(_01315_));
 sky130_fd_sc_hd__inv_2 _24982_ (.A(\decoded_imm[6] ),
    .Y(_20105_));
 sky130_fd_sc_hd__nor2_2 _24983_ (.A(_20103_),
    .B(_20105_),
    .Y(_01317_));
 sky130_fd_sc_hd__inv_2 _24984_ (.A(\decoded_imm[7] ),
    .Y(_20106_));
 sky130_fd_sc_hd__nor2_2 _24985_ (.A(_20103_),
    .B(_20106_),
    .Y(_01319_));
 sky130_fd_sc_hd__inv_2 _24986_ (.A(\decoded_imm[8] ),
    .Y(_20107_));
 sky130_fd_sc_hd__nor2_2 _24987_ (.A(_20103_),
    .B(_20107_),
    .Y(_01321_));
 sky130_fd_sc_hd__inv_2 _24988_ (.A(\decoded_imm[9] ),
    .Y(_20108_));
 sky130_fd_sc_hd__nor2_2 _24989_ (.A(_20103_),
    .B(_20108_),
    .Y(_01323_));
 sky130_fd_sc_hd__inv_2 _24990_ (.A(\decoded_imm[10] ),
    .Y(_20109_));
 sky130_fd_sc_hd__nor2_2 _24991_ (.A(_20103_),
    .B(_20109_),
    .Y(_01325_));
 sky130_fd_sc_hd__buf_1 _24992_ (.A(_19422_),
    .X(_20110_));
 sky130_fd_sc_hd__inv_2 _24993_ (.A(\decoded_imm[11] ),
    .Y(_20111_));
 sky130_fd_sc_hd__nor2_2 _24994_ (.A(_20110_),
    .B(_20111_),
    .Y(_01327_));
 sky130_fd_sc_hd__inv_2 _24995_ (.A(\decoded_imm[12] ),
    .Y(_20112_));
 sky130_fd_sc_hd__nor2_2 _24996_ (.A(_20110_),
    .B(_20112_),
    .Y(_01329_));
 sky130_fd_sc_hd__inv_2 _24997_ (.A(\decoded_imm[13] ),
    .Y(_20113_));
 sky130_fd_sc_hd__nor2_2 _24998_ (.A(_20110_),
    .B(_20113_),
    .Y(_01331_));
 sky130_fd_sc_hd__inv_2 _24999_ (.A(\decoded_imm[14] ),
    .Y(_20114_));
 sky130_fd_sc_hd__nor2_2 _25000_ (.A(_20110_),
    .B(_20114_),
    .Y(_01333_));
 sky130_fd_sc_hd__inv_2 _25001_ (.A(\decoded_imm[15] ),
    .Y(_20115_));
 sky130_fd_sc_hd__nor2_2 _25002_ (.A(_20110_),
    .B(_20115_),
    .Y(_01335_));
 sky130_fd_sc_hd__inv_2 _25003_ (.A(\decoded_imm[16] ),
    .Y(_20116_));
 sky130_fd_sc_hd__nor2_2 _25004_ (.A(_20110_),
    .B(_20116_),
    .Y(_01337_));
 sky130_fd_sc_hd__buf_1 _25005_ (.A(is_slli_srli_srai),
    .X(_20117_));
 sky130_fd_sc_hd__inv_2 _25006_ (.A(\decoded_imm[17] ),
    .Y(_20118_));
 sky130_fd_sc_hd__nor2_2 _25007_ (.A(_20117_),
    .B(_20118_),
    .Y(_01339_));
 sky130_fd_sc_hd__inv_2 _25008_ (.A(\decoded_imm[18] ),
    .Y(_20119_));
 sky130_fd_sc_hd__nor2_2 _25009_ (.A(_20117_),
    .B(_20119_),
    .Y(_01341_));
 sky130_fd_sc_hd__inv_2 _25010_ (.A(\decoded_imm[19] ),
    .Y(_20120_));
 sky130_fd_sc_hd__nor2_2 _25011_ (.A(_20117_),
    .B(_20120_),
    .Y(_01343_));
 sky130_fd_sc_hd__inv_2 _25012_ (.A(\decoded_imm[20] ),
    .Y(_20121_));
 sky130_fd_sc_hd__nor2_2 _25013_ (.A(_20117_),
    .B(_20121_),
    .Y(_01345_));
 sky130_fd_sc_hd__inv_2 _25014_ (.A(\decoded_imm[21] ),
    .Y(_20122_));
 sky130_fd_sc_hd__nor2_2 _25015_ (.A(_20117_),
    .B(_20122_),
    .Y(_01347_));
 sky130_fd_sc_hd__inv_2 _25016_ (.A(\decoded_imm[22] ),
    .Y(_20123_));
 sky130_fd_sc_hd__nor2_2 _25017_ (.A(_20117_),
    .B(_20123_),
    .Y(_01349_));
 sky130_fd_sc_hd__buf_1 _25018_ (.A(is_slli_srli_srai),
    .X(_20124_));
 sky130_fd_sc_hd__inv_2 _25019_ (.A(\decoded_imm[23] ),
    .Y(_20125_));
 sky130_fd_sc_hd__nor2_2 _25020_ (.A(_20124_),
    .B(_20125_),
    .Y(_01351_));
 sky130_fd_sc_hd__inv_2 _25021_ (.A(\decoded_imm[24] ),
    .Y(_20126_));
 sky130_fd_sc_hd__nor2_2 _25022_ (.A(_20124_),
    .B(_20126_),
    .Y(_01353_));
 sky130_fd_sc_hd__inv_2 _25023_ (.A(\decoded_imm[25] ),
    .Y(_20127_));
 sky130_fd_sc_hd__nor2_2 _25024_ (.A(_20124_),
    .B(_20127_),
    .Y(_01355_));
 sky130_fd_sc_hd__inv_2 _25025_ (.A(\decoded_imm[26] ),
    .Y(_20128_));
 sky130_fd_sc_hd__nor2_2 _25026_ (.A(_20124_),
    .B(_20128_),
    .Y(_01357_));
 sky130_fd_sc_hd__inv_2 _25027_ (.A(\decoded_imm[27] ),
    .Y(_20129_));
 sky130_fd_sc_hd__nor2_2 _25028_ (.A(_20124_),
    .B(_20129_),
    .Y(_01359_));
 sky130_fd_sc_hd__inv_2 _25029_ (.A(\decoded_imm[28] ),
    .Y(_20130_));
 sky130_fd_sc_hd__nor2_2 _25030_ (.A(_20124_),
    .B(_20130_),
    .Y(_01361_));
 sky130_fd_sc_hd__inv_2 _25031_ (.A(\decoded_imm[29] ),
    .Y(_20131_));
 sky130_fd_sc_hd__nor2_2 _25032_ (.A(_19422_),
    .B(_20131_),
    .Y(_01363_));
 sky130_fd_sc_hd__inv_2 _25033_ (.A(\decoded_imm[30] ),
    .Y(_20132_));
 sky130_fd_sc_hd__nor2_2 _25034_ (.A(_19422_),
    .B(_20132_),
    .Y(_01365_));
 sky130_fd_sc_hd__inv_2 _25035_ (.A(\decoded_imm[31] ),
    .Y(_20133_));
 sky130_fd_sc_hd__nor2_2 _25036_ (.A(_19422_),
    .B(_20133_),
    .Y(_01367_));
 sky130_fd_sc_hd__buf_1 _25037_ (.A(_19492_),
    .X(_20134_));
 sky130_fd_sc_hd__inv_2 _25038_ (.A(\reg_next_pc[0] ),
    .Y(_20135_));
 sky130_fd_sc_hd__nor2_2 _25039_ (.A(_20134_),
    .B(_20135_),
    .Y(_01369_));
 sky130_fd_sc_hd__inv_2 _25040_ (.A(\decoded_imm[0] ),
    .Y(_20136_));
 sky130_fd_sc_hd__nand2_2 _25041_ (.A(_20136_),
    .B(_19790_),
    .Y(_20137_));
 sky130_fd_sc_hd__nand2_2 _25042_ (.A(\decoded_imm[0] ),
    .B(pcpi_rs1[0]),
    .Y(_20138_));
 sky130_fd_sc_hd__and2_2 _25043_ (.A(_20137_),
    .B(_20138_),
    .X(_01371_));
 sky130_fd_sc_hd__nor2_2 _25044_ (.A(_20134_),
    .B(_18573_),
    .Y(_01372_));
 sky130_fd_sc_hd__nor2_2 _25045_ (.A(pcpi_rs1[1]),
    .B(\decoded_imm[1] ),
    .Y(_20139_));
 sky130_fd_sc_hd__nand2_2 _25046_ (.A(_19533_),
    .B(\decoded_imm[1] ),
    .Y(_20140_));
 sky130_fd_sc_hd__or2b_2 _25047_ (.A(_20139_),
    .B_N(_20140_),
    .X(_20141_));
 sky130_fd_sc_hd__xor2_2 _25048_ (.A(_20138_),
    .B(_20141_),
    .X(_01374_));
 sky130_fd_sc_hd__inv_2 _25049_ (.A(\reg_pc[2] ),
    .Y(_02073_));
 sky130_fd_sc_hd__nor2_2 _25050_ (.A(_20134_),
    .B(_02073_),
    .Y(_01375_));
 sky130_fd_sc_hd__nand2_2 _25051_ (.A(_19532_),
    .B(\decoded_imm[2] ),
    .Y(_20142_));
 sky130_fd_sc_hd__nand2_2 _25052_ (.A(_19915_),
    .B(_19702_),
    .Y(_20143_));
 sky130_fd_sc_hd__o21ai_2 _25053_ (.A1(_20138_),
    .A2(_20139_),
    .B1(_20140_),
    .Y(_20144_));
 sky130_fd_sc_hd__a21oi_2 _25054_ (.A1(_20142_),
    .A2(_20143_),
    .B1(_20144_),
    .Y(_20145_));
 sky130_fd_sc_hd__and3_2 _25055_ (.A(_20144_),
    .B(_20142_),
    .C(_20143_),
    .X(_20146_));
 sky130_fd_sc_hd__nor2_2 _25056_ (.A(_20145_),
    .B(_20146_),
    .Y(_01377_));
 sky130_fd_sc_hd__inv_2 _25057_ (.A(\reg_pc[3] ),
    .Y(_20147_));
 sky130_fd_sc_hd__nor2_2 _25058_ (.A(_20134_),
    .B(_20147_),
    .Y(_01378_));
 sky130_fd_sc_hd__nor2_2 _25059_ (.A(_19531_),
    .B(\decoded_imm[3] ),
    .Y(_20148_));
 sky130_fd_sc_hd__nor2_2 _25060_ (.A(_19911_),
    .B(_19708_),
    .Y(_20149_));
 sky130_fd_sc_hd__nor2_2 _25061_ (.A(_20148_),
    .B(_20149_),
    .Y(_20150_));
 sky130_fd_sc_hd__nand2_2 _25062_ (.A(_20144_),
    .B(_20143_),
    .Y(_20151_));
 sky130_fd_sc_hd__nand2_2 _25063_ (.A(_20151_),
    .B(_20142_),
    .Y(_20152_));
 sky130_fd_sc_hd__xor2_2 _25064_ (.A(_20150_),
    .B(_20152_),
    .X(_01380_));
 sky130_fd_sc_hd__inv_2 _25065_ (.A(\reg_pc[4] ),
    .Y(_20153_));
 sky130_fd_sc_hd__nor2_2 _25066_ (.A(_20134_),
    .B(_20153_),
    .Y(_01381_));
 sky130_fd_sc_hd__nor2_2 _25067_ (.A(pcpi_rs1[4]),
    .B(\decoded_imm[4] ),
    .Y(_20154_));
 sky130_fd_sc_hd__inv_2 _25068_ (.A(_20154_),
    .Y(_20155_));
 sky130_fd_sc_hd__nand2_2 _25069_ (.A(_19530_),
    .B(\decoded_imm[4] ),
    .Y(_20156_));
 sky130_fd_sc_hd__nand2_2 _25070_ (.A(_20155_),
    .B(_20156_),
    .Y(_20157_));
 sky130_fd_sc_hd__a21oi_2 _25071_ (.A1(_20151_),
    .A2(_20142_),
    .B1(_20148_),
    .Y(_20158_));
 sky130_fd_sc_hd__nor2_2 _25072_ (.A(_20149_),
    .B(_20158_),
    .Y(_20159_));
 sky130_fd_sc_hd__xor2_2 _25073_ (.A(_20157_),
    .B(_20159_),
    .X(_01383_));
 sky130_fd_sc_hd__buf_1 _25074_ (.A(_19492_),
    .X(_20160_));
 sky130_fd_sc_hd__inv_2 _25075_ (.A(\reg_pc[5] ),
    .Y(_20161_));
 sky130_fd_sc_hd__nor2_2 _25076_ (.A(_20160_),
    .B(_20161_),
    .Y(_01384_));
 sky130_fd_sc_hd__nor2_2 _25077_ (.A(_19529_),
    .B(\decoded_imm[5] ),
    .Y(_20162_));
 sky130_fd_sc_hd__nor2_2 _25078_ (.A(_19918_),
    .B(_20104_),
    .Y(_20163_));
 sky130_fd_sc_hd__nor2_2 _25079_ (.A(_20162_),
    .B(_20163_),
    .Y(_20164_));
 sky130_fd_sc_hd__o21ai_2 _25080_ (.A1(_20149_),
    .A2(_20158_),
    .B1(_20155_),
    .Y(_20165_));
 sky130_fd_sc_hd__nand2_2 _25081_ (.A(_20165_),
    .B(_20156_),
    .Y(_20166_));
 sky130_fd_sc_hd__xor2_2 _25082_ (.A(_20164_),
    .B(_20166_),
    .X(_01386_));
 sky130_fd_sc_hd__nor2_2 _25083_ (.A(_20160_),
    .B(_18564_),
    .Y(_01387_));
 sky130_fd_sc_hd__xor2_2 _25084_ (.A(pcpi_rs1[6]),
    .B(\decoded_imm[6] ),
    .X(_20167_));
 sky130_fd_sc_hd__a21oi_2 _25085_ (.A1(_20165_),
    .A2(_20156_),
    .B1(_20162_),
    .Y(_20168_));
 sky130_fd_sc_hd__or2_2 _25086_ (.A(_20163_),
    .B(_20168_),
    .X(_20169_));
 sky130_fd_sc_hd__or2_2 _25087_ (.A(_20167_),
    .B(_20169_),
    .X(_20170_));
 sky130_fd_sc_hd__nand2_2 _25088_ (.A(_20169_),
    .B(_20167_),
    .Y(_20171_));
 sky130_fd_sc_hd__and2_2 _25089_ (.A(_20170_),
    .B(_20171_),
    .X(_01389_));
 sky130_fd_sc_hd__inv_2 _25090_ (.A(\reg_pc[7] ),
    .Y(_20172_));
 sky130_fd_sc_hd__nor2_2 _25091_ (.A(_20160_),
    .B(_20172_),
    .Y(_01390_));
 sky130_fd_sc_hd__nor2_2 _25092_ (.A(pcpi_rs1[7]),
    .B(\decoded_imm[7] ),
    .Y(_20173_));
 sky130_fd_sc_hd__nor2_2 _25093_ (.A(_19862_),
    .B(_20106_),
    .Y(_20174_));
 sky130_fd_sc_hd__nor2_2 _25094_ (.A(_20173_),
    .B(_20174_),
    .Y(_20175_));
 sky130_fd_sc_hd__o21ai_2 _25095_ (.A1(_19858_),
    .A2(_20105_),
    .B1(_20171_),
    .Y(_20176_));
 sky130_fd_sc_hd__xor2_2 _25096_ (.A(_20175_),
    .B(_20176_),
    .X(_01392_));
 sky130_fd_sc_hd__inv_2 _25097_ (.A(\reg_pc[8] ),
    .Y(_20177_));
 sky130_fd_sc_hd__nor2_2 _25098_ (.A(_20160_),
    .B(_20177_),
    .Y(_01393_));
 sky130_fd_sc_hd__nor2_2 _25099_ (.A(_19526_),
    .B(\decoded_imm[8] ),
    .Y(_20178_));
 sky130_fd_sc_hd__nor2_2 _25100_ (.A(_19898_),
    .B(_20107_),
    .Y(_20179_));
 sky130_fd_sc_hd__nor2_2 _25101_ (.A(_20178_),
    .B(_20179_),
    .Y(_20180_));
 sky130_fd_sc_hd__o211ai_2 _25102_ (.A1(_20163_),
    .A2(_20168_),
    .B1(_20167_),
    .C1(_20175_),
    .Y(_20181_));
 sky130_fd_sc_hd__nor2_2 _25103_ (.A(_20105_),
    .B(_20173_),
    .Y(_20182_));
 sky130_fd_sc_hd__a21oi_2 _25104_ (.A1(_20182_),
    .A2(_19528_),
    .B1(_20174_),
    .Y(_20183_));
 sky130_fd_sc_hd__nand2_2 _25105_ (.A(_20181_),
    .B(_20183_),
    .Y(_20184_));
 sky130_fd_sc_hd__xor2_2 _25106_ (.A(_20180_),
    .B(_20184_),
    .X(_01395_));
 sky130_fd_sc_hd__inv_2 _25107_ (.A(\reg_pc[9] ),
    .Y(_20185_));
 sky130_fd_sc_hd__nor2_2 _25108_ (.A(_20160_),
    .B(_20185_),
    .Y(_01396_));
 sky130_fd_sc_hd__nor2_2 _25109_ (.A(_19525_),
    .B(\decoded_imm[9] ),
    .Y(_20186_));
 sky130_fd_sc_hd__nor2_2 _25110_ (.A(_19894_),
    .B(_20108_),
    .Y(_20187_));
 sky130_fd_sc_hd__nor2_2 _25111_ (.A(_20186_),
    .B(_20187_),
    .Y(_20188_));
 sky130_fd_sc_hd__inv_2 _25112_ (.A(_20178_),
    .Y(_20189_));
 sky130_fd_sc_hd__a21oi_2 _25113_ (.A1(_20184_),
    .A2(_20189_),
    .B1(_20179_),
    .Y(_20190_));
 sky130_fd_sc_hd__xnor2_2 _25114_ (.A(_20188_),
    .B(_20190_),
    .Y(_01398_));
 sky130_fd_sc_hd__inv_2 _25115_ (.A(\reg_pc[10] ),
    .Y(_20191_));
 sky130_fd_sc_hd__nor2_2 _25116_ (.A(_20160_),
    .B(_20191_),
    .Y(_01399_));
 sky130_fd_sc_hd__nor2_2 _25117_ (.A(pcpi_rs1[10]),
    .B(\decoded_imm[10] ),
    .Y(_20192_));
 sky130_fd_sc_hd__nor2_2 _25118_ (.A(_19902_),
    .B(_20109_),
    .Y(_20193_));
 sky130_fd_sc_hd__nor2_2 _25119_ (.A(_20192_),
    .B(_20193_),
    .Y(_20194_));
 sky130_fd_sc_hd__nor2_2 _25120_ (.A(_20107_),
    .B(_20186_),
    .Y(_20195_));
 sky130_fd_sc_hd__a21o_2 _25121_ (.A1(_20195_),
    .A2(_19526_),
    .B1(_20187_),
    .X(_20196_));
 sky130_fd_sc_hd__nand2_2 _25122_ (.A(_20180_),
    .B(_20188_),
    .Y(_20197_));
 sky130_fd_sc_hd__a21oi_2 _25123_ (.A1(_20181_),
    .A2(_20183_),
    .B1(_20197_),
    .Y(_20198_));
 sky130_fd_sc_hd__nor3_2 _25124_ (.A(_20194_),
    .B(_20196_),
    .C(_20198_),
    .Y(_20199_));
 sky130_fd_sc_hd__o21ai_2 _25125_ (.A1(_20196_),
    .A2(_20198_),
    .B1(_20194_),
    .Y(_20200_));
 sky130_fd_sc_hd__nor2b_2 _25126_ (.A(_20199_),
    .B_N(_20200_),
    .Y(_01401_));
 sky130_fd_sc_hd__buf_1 _25127_ (.A(_19492_),
    .X(_20201_));
 sky130_fd_sc_hd__nor2_2 _25128_ (.A(_20201_),
    .B(_18552_),
    .Y(_01402_));
 sky130_fd_sc_hd__inv_2 _25129_ (.A(_20193_),
    .Y(_20202_));
 sky130_fd_sc_hd__nor2_2 _25130_ (.A(_19524_),
    .B(\decoded_imm[11] ),
    .Y(_20203_));
 sky130_fd_sc_hd__nor2_2 _25131_ (.A(_19890_),
    .B(_20111_),
    .Y(_20204_));
 sky130_fd_sc_hd__or2_2 _25132_ (.A(_20203_),
    .B(_20204_),
    .X(_20205_));
 sky130_fd_sc_hd__a21oi_2 _25133_ (.A1(_20200_),
    .A2(_20202_),
    .B1(_20205_),
    .Y(_20206_));
 sky130_fd_sc_hd__and3_2 _25134_ (.A(_20200_),
    .B(_20202_),
    .C(_20205_),
    .X(_20207_));
 sky130_fd_sc_hd__nor2_2 _25135_ (.A(_20206_),
    .B(_20207_),
    .Y(_01404_));
 sky130_fd_sc_hd__inv_2 _25136_ (.A(\reg_pc[12] ),
    .Y(_20208_));
 sky130_fd_sc_hd__nor2_2 _25137_ (.A(_20201_),
    .B(_20208_),
    .Y(_01405_));
 sky130_fd_sc_hd__nor2_2 _25138_ (.A(_20204_),
    .B(_20206_),
    .Y(_20209_));
 sky130_fd_sc_hd__nor2_2 _25139_ (.A(_19523_),
    .B(\decoded_imm[12] ),
    .Y(_20210_));
 sky130_fd_sc_hd__nor2_2 _25140_ (.A(_19881_),
    .B(_20112_),
    .Y(_20211_));
 sky130_fd_sc_hd__or2_2 _25141_ (.A(_20210_),
    .B(_20211_),
    .X(_20212_));
 sky130_fd_sc_hd__nand2_2 _25142_ (.A(_20209_),
    .B(_20212_),
    .Y(_20213_));
 sky130_fd_sc_hd__o21bai_2 _25143_ (.A1(_20204_),
    .A2(_20206_),
    .B1_N(_20212_),
    .Y(_20214_));
 sky130_fd_sc_hd__and2_2 _25144_ (.A(_20213_),
    .B(_20214_),
    .X(_01407_));
 sky130_fd_sc_hd__inv_2 _25145_ (.A(\reg_pc[13] ),
    .Y(_20215_));
 sky130_fd_sc_hd__nor2_2 _25146_ (.A(_20201_),
    .B(_20215_),
    .Y(_01408_));
 sky130_fd_sc_hd__inv_2 _25147_ (.A(_20211_),
    .Y(_20216_));
 sky130_fd_sc_hd__nor2_2 _25148_ (.A(_19521_),
    .B(\decoded_imm[13] ),
    .Y(_20217_));
 sky130_fd_sc_hd__nor2_2 _25149_ (.A(_19877_),
    .B(_20113_),
    .Y(_20218_));
 sky130_fd_sc_hd__or2_2 _25150_ (.A(_20217_),
    .B(_20218_),
    .X(_20219_));
 sky130_fd_sc_hd__a21oi_2 _25151_ (.A1(_20214_),
    .A2(_20216_),
    .B1(_20219_),
    .Y(_20220_));
 sky130_fd_sc_hd__and3_2 _25152_ (.A(_20214_),
    .B(_20216_),
    .C(_20219_),
    .X(_20221_));
 sky130_fd_sc_hd__nor2_2 _25153_ (.A(_20220_),
    .B(_20221_),
    .Y(_01410_));
 sky130_fd_sc_hd__inv_2 _25154_ (.A(\reg_pc[14] ),
    .Y(_20222_));
 sky130_fd_sc_hd__nor2_2 _25155_ (.A(_20201_),
    .B(_20222_),
    .Y(_01411_));
 sky130_fd_sc_hd__nor2_2 _25156_ (.A(pcpi_rs1[14]),
    .B(_20114_),
    .Y(_20223_));
 sky130_fd_sc_hd__nor2_2 _25157_ (.A(\decoded_imm[14] ),
    .B(_19885_),
    .Y(_20224_));
 sky130_fd_sc_hd__or4_2 _25158_ (.A(_20218_),
    .B(_20223_),
    .C(_20224_),
    .D(_20220_),
    .X(_20225_));
 sky130_fd_sc_hd__o22ai_2 _25159_ (.A1(_20223_),
    .A2(_20224_),
    .B1(_20218_),
    .B2(_20220_),
    .Y(_20226_));
 sky130_fd_sc_hd__and2_2 _25160_ (.A(_20225_),
    .B(_20226_),
    .X(_01413_));
 sky130_fd_sc_hd__inv_2 _25161_ (.A(\reg_pc[15] ),
    .Y(_20227_));
 sky130_fd_sc_hd__nor2_2 _25162_ (.A(_20201_),
    .B(_20227_),
    .Y(_01414_));
 sky130_fd_sc_hd__nor2_2 _25163_ (.A(_19885_),
    .B(_20114_),
    .Y(_20228_));
 sky130_fd_sc_hd__inv_2 _25164_ (.A(_20228_),
    .Y(_20229_));
 sky130_fd_sc_hd__nor2_2 _25165_ (.A(_19520_),
    .B(\decoded_imm[15] ),
    .Y(_20230_));
 sky130_fd_sc_hd__nor2_2 _25166_ (.A(_19873_),
    .B(_20115_),
    .Y(_20231_));
 sky130_fd_sc_hd__or2_2 _25167_ (.A(_20230_),
    .B(_20231_),
    .X(_20232_));
 sky130_fd_sc_hd__a21oi_2 _25168_ (.A1(_20226_),
    .A2(_20229_),
    .B1(_20232_),
    .Y(_20233_));
 sky130_fd_sc_hd__and3_2 _25169_ (.A(_20226_),
    .B(_20229_),
    .C(_20232_),
    .X(_20234_));
 sky130_fd_sc_hd__nor2_2 _25170_ (.A(_20233_),
    .B(_20234_),
    .Y(_01416_));
 sky130_fd_sc_hd__inv_2 _25171_ (.A(\reg_pc[16] ),
    .Y(_20235_));
 sky130_fd_sc_hd__nor2_2 _25172_ (.A(_20201_),
    .B(_20235_),
    .Y(_01417_));
 sky130_fd_sc_hd__nor2_2 _25173_ (.A(pcpi_rs1[16]),
    .B(\decoded_imm[16] ),
    .Y(_20236_));
 sky130_fd_sc_hd__inv_2 _25174_ (.A(pcpi_rs1[16]),
    .Y(_20237_));
 sky130_fd_sc_hd__nor2_2 _25175_ (.A(_20237_),
    .B(_20116_),
    .Y(_20238_));
 sky130_fd_sc_hd__or2_2 _25176_ (.A(_20236_),
    .B(_20238_),
    .X(_20239_));
 sky130_fd_sc_hd__nor2_2 _25177_ (.A(_20231_),
    .B(_20233_),
    .Y(_20240_));
 sky130_fd_sc_hd__xor2_2 _25178_ (.A(_20239_),
    .B(_20240_),
    .X(_01419_));
 sky130_fd_sc_hd__buf_1 _25179_ (.A(instr_lui),
    .X(_20241_));
 sky130_fd_sc_hd__inv_2 _25180_ (.A(\reg_pc[17] ),
    .Y(_20242_));
 sky130_fd_sc_hd__nor2_2 _25181_ (.A(_20241_),
    .B(_20242_),
    .Y(_01420_));
 sky130_fd_sc_hd__nor2_2 _25182_ (.A(_19518_),
    .B(\decoded_imm[17] ),
    .Y(_20243_));
 sky130_fd_sc_hd__nor2_2 _25183_ (.A(_19983_),
    .B(_20118_),
    .Y(_20244_));
 sky130_fd_sc_hd__nor2_2 _25184_ (.A(_20243_),
    .B(_20244_),
    .Y(_20245_));
 sky130_fd_sc_hd__inv_2 _25185_ (.A(_20245_),
    .Y(_20246_));
 sky130_fd_sc_hd__o21ba_2 _25186_ (.A1(_20236_),
    .A2(_20240_),
    .B1_N(_20238_),
    .X(_20247_));
 sky130_fd_sc_hd__xor2_2 _25187_ (.A(_20246_),
    .B(_20247_),
    .X(_01422_));
 sky130_fd_sc_hd__inv_2 _25188_ (.A(\reg_pc[18] ),
    .Y(_20248_));
 sky130_fd_sc_hd__nor2_2 _25189_ (.A(_20241_),
    .B(_20248_),
    .Y(_01423_));
 sky130_fd_sc_hd__nor2_2 _25190_ (.A(_19517_),
    .B(\decoded_imm[18] ),
    .Y(_20249_));
 sky130_fd_sc_hd__nor2_2 _25191_ (.A(_19993_),
    .B(_20119_),
    .Y(_20250_));
 sky130_fd_sc_hd__nor2_2 _25192_ (.A(_20249_),
    .B(_20250_),
    .Y(_20251_));
 sky130_fd_sc_hd__nor2_2 _25193_ (.A(_20239_),
    .B(_20246_),
    .Y(_20252_));
 sky130_fd_sc_hd__o21ai_2 _25194_ (.A1(_20231_),
    .A2(_20233_),
    .B1(_20252_),
    .Y(_20253_));
 sky130_fd_sc_hd__nor2_2 _25195_ (.A(_20116_),
    .B(_20243_),
    .Y(_20254_));
 sky130_fd_sc_hd__a21oi_2 _25196_ (.A1(_20254_),
    .A2(_19519_),
    .B1(_20244_),
    .Y(_20255_));
 sky130_fd_sc_hd__nand2_2 _25197_ (.A(_20253_),
    .B(_20255_),
    .Y(_20256_));
 sky130_fd_sc_hd__xor2_2 _25198_ (.A(_20251_),
    .B(_20256_),
    .X(_01425_));
 sky130_fd_sc_hd__inv_2 _25199_ (.A(\reg_pc[19] ),
    .Y(_20257_));
 sky130_fd_sc_hd__nor2_2 _25200_ (.A(_20241_),
    .B(_20257_),
    .Y(_01426_));
 sky130_fd_sc_hd__nor2_2 _25201_ (.A(_19515_),
    .B(_20120_),
    .Y(_20258_));
 sky130_fd_sc_hd__nor2_2 _25202_ (.A(\decoded_imm[19] ),
    .B(_19988_),
    .Y(_20259_));
 sky130_fd_sc_hd__a21oi_2 _25203_ (.A1(_20253_),
    .A2(_20255_),
    .B1(_20249_),
    .Y(_20260_));
 sky130_fd_sc_hd__or4_2 _25204_ (.A(_20250_),
    .B(_20258_),
    .C(_20259_),
    .D(_20260_),
    .X(_20261_));
 sky130_fd_sc_hd__o22ai_2 _25205_ (.A1(_20258_),
    .A2(_20259_),
    .B1(_20250_),
    .B2(_20260_),
    .Y(_20262_));
 sky130_fd_sc_hd__and2_2 _25206_ (.A(_20261_),
    .B(_20262_),
    .X(_01428_));
 sky130_fd_sc_hd__inv_2 _25207_ (.A(\reg_pc[20] ),
    .Y(_20263_));
 sky130_fd_sc_hd__nor2_2 _25208_ (.A(_20241_),
    .B(_20263_),
    .Y(_01429_));
 sky130_fd_sc_hd__nor2_2 _25209_ (.A(_19988_),
    .B(_20120_),
    .Y(_20264_));
 sky130_fd_sc_hd__inv_2 _25210_ (.A(_20264_),
    .Y(_20265_));
 sky130_fd_sc_hd__nor2_2 _25211_ (.A(pcpi_rs1[20]),
    .B(\decoded_imm[20] ),
    .Y(_20266_));
 sky130_fd_sc_hd__nor2_2 _25212_ (.A(_19939_),
    .B(_20121_),
    .Y(_20267_));
 sky130_fd_sc_hd__nor2_2 _25213_ (.A(_20266_),
    .B(_20267_),
    .Y(_20268_));
 sky130_fd_sc_hd__inv_2 _25214_ (.A(_20268_),
    .Y(_20269_));
 sky130_fd_sc_hd__a21oi_2 _25215_ (.A1(_20262_),
    .A2(_20265_),
    .B1(_20269_),
    .Y(_20270_));
 sky130_fd_sc_hd__and3_2 _25216_ (.A(_20262_),
    .B(_20265_),
    .C(_20269_),
    .X(_20271_));
 sky130_fd_sc_hd__nor2_2 _25217_ (.A(_20270_),
    .B(_20271_),
    .Y(_01431_));
 sky130_fd_sc_hd__inv_2 _25218_ (.A(\reg_pc[21] ),
    .Y(_20272_));
 sky130_fd_sc_hd__nor2_2 _25219_ (.A(_20241_),
    .B(_20272_),
    .Y(_01432_));
 sky130_fd_sc_hd__nor2_2 _25220_ (.A(_19514_),
    .B(_20122_),
    .Y(_20273_));
 sky130_fd_sc_hd__nor2_2 _25221_ (.A(\decoded_imm[21] ),
    .B(_19926_),
    .Y(_20274_));
 sky130_fd_sc_hd__or4_2 _25222_ (.A(_20267_),
    .B(_20273_),
    .C(_20274_),
    .D(_20270_),
    .X(_20275_));
 sky130_fd_sc_hd__o22ai_2 _25223_ (.A1(_20273_),
    .A2(_20274_),
    .B1(_20267_),
    .B2(_20270_),
    .Y(_20276_));
 sky130_fd_sc_hd__and2_2 _25224_ (.A(_20275_),
    .B(_20276_),
    .X(_01434_));
 sky130_fd_sc_hd__inv_2 _25225_ (.A(\reg_pc[22] ),
    .Y(_20277_));
 sky130_fd_sc_hd__nor2_2 _25226_ (.A(_20241_),
    .B(_20277_),
    .Y(_01435_));
 sky130_fd_sc_hd__nand2_2 _25227_ (.A(_19514_),
    .B(\decoded_imm[21] ),
    .Y(_20278_));
 sky130_fd_sc_hd__nor2_2 _25228_ (.A(pcpi_rs1[22]),
    .B(\decoded_imm[22] ),
    .Y(_20279_));
 sky130_fd_sc_hd__nor2_2 _25229_ (.A(_19935_),
    .B(_20123_),
    .Y(_20280_));
 sky130_fd_sc_hd__nor2_2 _25230_ (.A(_20279_),
    .B(_20280_),
    .Y(_20281_));
 sky130_fd_sc_hd__inv_2 _25231_ (.A(_20281_),
    .Y(_20282_));
 sky130_fd_sc_hd__a21oi_2 _25232_ (.A1(_20276_),
    .A2(_20278_),
    .B1(_20282_),
    .Y(_20283_));
 sky130_fd_sc_hd__and3_2 _25233_ (.A(_20276_),
    .B(_20278_),
    .C(_20282_),
    .X(_20284_));
 sky130_fd_sc_hd__nor2_2 _25234_ (.A(_20283_),
    .B(_20284_),
    .Y(_01437_));
 sky130_fd_sc_hd__buf_1 _25235_ (.A(instr_lui),
    .X(_20285_));
 sky130_fd_sc_hd__inv_2 _25236_ (.A(\reg_pc[23] ),
    .Y(_20286_));
 sky130_fd_sc_hd__nor2_2 _25237_ (.A(_20285_),
    .B(_20286_),
    .Y(_01438_));
 sky130_fd_sc_hd__nor2_2 _25238_ (.A(_19512_),
    .B(_20125_),
    .Y(_20287_));
 sky130_fd_sc_hd__nor2_2 _25239_ (.A(\decoded_imm[23] ),
    .B(_19930_),
    .Y(_20288_));
 sky130_fd_sc_hd__or4_2 _25240_ (.A(_20280_),
    .B(_20287_),
    .C(_20288_),
    .D(_20283_),
    .X(_20289_));
 sky130_fd_sc_hd__o22ai_2 _25241_ (.A1(_20287_),
    .A2(_20288_),
    .B1(_20280_),
    .B2(_20283_),
    .Y(_20290_));
 sky130_fd_sc_hd__and2_2 _25242_ (.A(_20289_),
    .B(_20290_),
    .X(_01440_));
 sky130_fd_sc_hd__inv_2 _25243_ (.A(\reg_pc[24] ),
    .Y(_20291_));
 sky130_fd_sc_hd__nor2_2 _25244_ (.A(_20285_),
    .B(_20291_),
    .Y(_01441_));
 sky130_fd_sc_hd__xor2_2 _25245_ (.A(_19511_),
    .B(\decoded_imm[24] ),
    .X(_20292_));
 sky130_fd_sc_hd__nand2_2 _25246_ (.A(_19512_),
    .B(\decoded_imm[23] ),
    .Y(_20293_));
 sky130_fd_sc_hd__nand2_2 _25247_ (.A(_20290_),
    .B(_20293_),
    .Y(_20294_));
 sky130_fd_sc_hd__or2_2 _25248_ (.A(_20292_),
    .B(_20294_),
    .X(_20295_));
 sky130_fd_sc_hd__nand2_2 _25249_ (.A(_20294_),
    .B(_20292_),
    .Y(_20296_));
 sky130_fd_sc_hd__and2_2 _25250_ (.A(_20295_),
    .B(_20296_),
    .X(_01443_));
 sky130_fd_sc_hd__inv_2 _25251_ (.A(\reg_pc[25] ),
    .Y(_20297_));
 sky130_fd_sc_hd__nor2_2 _25252_ (.A(_20285_),
    .B(_20297_),
    .Y(_01444_));
 sky130_fd_sc_hd__nor2_2 _25253_ (.A(_19509_),
    .B(\decoded_imm[25] ),
    .Y(_20298_));
 sky130_fd_sc_hd__nor2_2 _25254_ (.A(_19945_),
    .B(_20127_),
    .Y(_20299_));
 sky130_fd_sc_hd__or2_2 _25255_ (.A(_20298_),
    .B(_20299_),
    .X(_20300_));
 sky130_fd_sc_hd__inv_2 _25256_ (.A(_20300_),
    .Y(_20301_));
 sky130_fd_sc_hd__o21ai_2 _25257_ (.A1(_19957_),
    .A2(_20126_),
    .B1(_20296_),
    .Y(_20302_));
 sky130_fd_sc_hd__xor2_2 _25258_ (.A(_20301_),
    .B(_20302_),
    .X(_01446_));
 sky130_fd_sc_hd__inv_2 _25259_ (.A(\reg_pc[26] ),
    .Y(_20303_));
 sky130_fd_sc_hd__nor2_2 _25260_ (.A(_20285_),
    .B(_20303_),
    .Y(_01447_));
 sky130_fd_sc_hd__nor2_2 _25261_ (.A(_19508_),
    .B(\decoded_imm[26] ),
    .Y(_20304_));
 sky130_fd_sc_hd__nor2_2 _25262_ (.A(_19952_),
    .B(_20128_),
    .Y(_20305_));
 sky130_fd_sc_hd__nor2_2 _25263_ (.A(_20304_),
    .B(_20305_),
    .Y(_20306_));
 sky130_fd_sc_hd__nor2_2 _25264_ (.A(_20126_),
    .B(_20298_),
    .Y(_20307_));
 sky130_fd_sc_hd__a21o_2 _25265_ (.A1(_20307_),
    .A2(_19511_),
    .B1(_20299_),
    .X(_20308_));
 sky130_fd_sc_hd__nand2_2 _25266_ (.A(_20301_),
    .B(_20292_),
    .Y(_20309_));
 sky130_fd_sc_hd__a21oi_2 _25267_ (.A1(_20290_),
    .A2(_20293_),
    .B1(_20309_),
    .Y(_20310_));
 sky130_fd_sc_hd__or2_2 _25268_ (.A(_20308_),
    .B(_20310_),
    .X(_20311_));
 sky130_fd_sc_hd__xor2_2 _25269_ (.A(_20306_),
    .B(_20311_),
    .X(_01449_));
 sky130_fd_sc_hd__inv_2 _25270_ (.A(\reg_pc[27] ),
    .Y(_20312_));
 sky130_fd_sc_hd__nor2_2 _25271_ (.A(_20285_),
    .B(_20312_),
    .Y(_01450_));
 sky130_fd_sc_hd__nor2_2 _25272_ (.A(pcpi_rs1[27]),
    .B(\decoded_imm[27] ),
    .Y(_20313_));
 sky130_fd_sc_hd__nor2_2 _25273_ (.A(_19967_),
    .B(_20129_),
    .Y(_20314_));
 sky130_fd_sc_hd__nor2_2 _25274_ (.A(_20313_),
    .B(_20314_),
    .Y(_20315_));
 sky130_fd_sc_hd__a21oi_2 _25275_ (.A1(_20311_),
    .A2(_20306_),
    .B1(_20305_),
    .Y(_20316_));
 sky130_fd_sc_hd__xnor2_2 _25276_ (.A(_20315_),
    .B(_20316_),
    .Y(_01452_));
 sky130_fd_sc_hd__inv_2 _25277_ (.A(\reg_pc[28] ),
    .Y(_20317_));
 sky130_fd_sc_hd__nor2_2 _25278_ (.A(_20285_),
    .B(_20317_),
    .Y(_01453_));
 sky130_fd_sc_hd__nand2_2 _25279_ (.A(_20306_),
    .B(_20315_),
    .Y(_20318_));
 sky130_fd_sc_hd__o21bai_2 _25280_ (.A1(_20308_),
    .A2(_20310_),
    .B1_N(_20318_),
    .Y(_20319_));
 sky130_fd_sc_hd__nor2_2 _25281_ (.A(_20128_),
    .B(_20313_),
    .Y(_20320_));
 sky130_fd_sc_hd__a21oi_2 _25282_ (.A1(_20320_),
    .A2(_19508_),
    .B1(_20314_),
    .Y(_20321_));
 sky130_fd_sc_hd__nor2_2 _25283_ (.A(_19507_),
    .B(\decoded_imm[28] ),
    .Y(_20322_));
 sky130_fd_sc_hd__nor2_2 _25284_ (.A(_19949_),
    .B(_20130_),
    .Y(_20323_));
 sky130_fd_sc_hd__or2_2 _25285_ (.A(_20322_),
    .B(_20323_),
    .X(_20324_));
 sky130_fd_sc_hd__a21oi_2 _25286_ (.A1(_20319_),
    .A2(_20321_),
    .B1(_20324_),
    .Y(_20325_));
 sky130_fd_sc_hd__and3_2 _25287_ (.A(_20319_),
    .B(_20321_),
    .C(_20324_),
    .X(_20326_));
 sky130_fd_sc_hd__nor2_2 _25288_ (.A(_20325_),
    .B(_20326_),
    .Y(_01455_));
 sky130_fd_sc_hd__inv_2 _25289_ (.A(\reg_pc[29] ),
    .Y(_20327_));
 sky130_fd_sc_hd__nor2_2 _25290_ (.A(_19492_),
    .B(_20327_),
    .Y(_01456_));
 sky130_fd_sc_hd__nand2_2 _25291_ (.A(_19963_),
    .B(_20131_),
    .Y(_20328_));
 sky130_fd_sc_hd__nand2_2 _25292_ (.A(_19506_),
    .B(\decoded_imm[29] ),
    .Y(_20329_));
 sky130_fd_sc_hd__nand2_2 _25293_ (.A(_20328_),
    .B(_20329_),
    .Y(_20330_));
 sky130_fd_sc_hd__a22oi_2 _25294_ (.A1(_19949_),
    .A2(_20130_),
    .B1(_20319_),
    .B2(_20321_),
    .Y(_20331_));
 sky130_fd_sc_hd__or3_2 _25295_ (.A(_20323_),
    .B(_20330_),
    .C(_20331_),
    .X(_20332_));
 sky130_fd_sc_hd__o21ai_2 _25296_ (.A1(_20323_),
    .A2(_20331_),
    .B1(_20330_),
    .Y(_20333_));
 sky130_fd_sc_hd__nand2_2 _25297_ (.A(_20332_),
    .B(_20333_),
    .Y(_01458_));
 sky130_fd_sc_hd__nor2_2 _25298_ (.A(_19492_),
    .B(_18505_),
    .Y(_01459_));
 sky130_fd_sc_hd__o22ai_2 _25299_ (.A1(_19506_),
    .A2(\decoded_imm[29] ),
    .B1(_20323_),
    .B2(_20331_),
    .Y(_20334_));
 sky130_fd_sc_hd__nor2_2 _25300_ (.A(_19505_),
    .B(\decoded_imm[30] ),
    .Y(_20335_));
 sky130_fd_sc_hd__nor2_2 _25301_ (.A(_19975_),
    .B(_20132_),
    .Y(_20336_));
 sky130_fd_sc_hd__nor2_2 _25302_ (.A(_20335_),
    .B(_20336_),
    .Y(_20337_));
 sky130_fd_sc_hd__inv_2 _25303_ (.A(_20337_),
    .Y(_20338_));
 sky130_fd_sc_hd__a21oi_2 _25304_ (.A1(_20334_),
    .A2(_20329_),
    .B1(_20338_),
    .Y(_20339_));
 sky130_fd_sc_hd__nand2_2 _25305_ (.A(_20334_),
    .B(_20329_),
    .Y(_20340_));
 sky130_fd_sc_hd__nor2_2 _25306_ (.A(_20337_),
    .B(_20340_),
    .Y(_20341_));
 sky130_fd_sc_hd__nor2_2 _25307_ (.A(_20339_),
    .B(_20341_),
    .Y(_01461_));
 sky130_fd_sc_hd__nor2b_2 _25308_ (.A(_20134_),
    .B_N(\reg_pc[31] ),
    .Y(_01462_));
 sky130_fd_sc_hd__nor2_2 _25309_ (.A(pcpi_rs1[31]),
    .B(\decoded_imm[31] ),
    .Y(_20342_));
 sky130_fd_sc_hd__nor2_2 _25310_ (.A(_18173_),
    .B(_20133_),
    .Y(_20343_));
 sky130_fd_sc_hd__o22ai_2 _25311_ (.A1(_20342_),
    .A2(_20343_),
    .B1(_20336_),
    .B2(_20339_),
    .Y(_20344_));
 sky130_fd_sc_hd__or3_2 _25312_ (.A(_20342_),
    .B(_20336_),
    .C(_20343_),
    .X(_20345_));
 sky130_fd_sc_hd__a21o_2 _25313_ (.A1(_20340_),
    .A2(_20337_),
    .B1(_20345_),
    .X(_20346_));
 sky130_fd_sc_hd__nand2_2 _25314_ (.A(_20344_),
    .B(_20346_),
    .Y(_01464_));
 sky130_fd_sc_hd__and2_2 _25315_ (.A(_20020_),
    .B(_01466_),
    .X(_01467_));
 sky130_fd_sc_hd__and2_2 _25316_ (.A(_20020_),
    .B(_01469_),
    .X(_01470_));
 sky130_fd_sc_hd__buf_1 _25317_ (.A(_18243_),
    .X(_20347_));
 sky130_fd_sc_hd__a21oi_2 _25318_ (.A1(_20020_),
    .A2(_01473_),
    .B1(_20347_),
    .Y(_01474_));
 sky130_fd_sc_hd__and2_2 _25319_ (.A(_20020_),
    .B(_01477_),
    .X(_01478_));
 sky130_fd_sc_hd__buf_1 _25320_ (.A(_20019_),
    .X(_20348_));
 sky130_fd_sc_hd__and2_2 _25321_ (.A(_20348_),
    .B(_01480_),
    .X(_01481_));
 sky130_fd_sc_hd__and2_2 _25322_ (.A(_20348_),
    .B(_01483_),
    .X(_01484_));
 sky130_fd_sc_hd__and2_2 _25323_ (.A(_20348_),
    .B(_01486_),
    .X(_01487_));
 sky130_fd_sc_hd__and2_2 _25324_ (.A(_20348_),
    .B(_01489_),
    .X(_01490_));
 sky130_fd_sc_hd__and2_2 _25325_ (.A(_20348_),
    .B(_01492_),
    .X(_01493_));
 sky130_fd_sc_hd__and2_2 _25326_ (.A(_20348_),
    .B(_01495_),
    .X(_01496_));
 sky130_fd_sc_hd__buf_1 _25327_ (.A(_20019_),
    .X(_20349_));
 sky130_fd_sc_hd__and2_2 _25328_ (.A(_20349_),
    .B(_01498_),
    .X(_01499_));
 sky130_fd_sc_hd__and2_2 _25329_ (.A(_20349_),
    .B(_01501_),
    .X(_01502_));
 sky130_fd_sc_hd__and2_2 _25330_ (.A(_20349_),
    .B(_01504_),
    .X(_01505_));
 sky130_fd_sc_hd__and2_2 _25331_ (.A(_20349_),
    .B(_01507_),
    .X(_01508_));
 sky130_fd_sc_hd__and2_2 _25332_ (.A(_20349_),
    .B(_01510_),
    .X(_01511_));
 sky130_fd_sc_hd__and2_2 _25333_ (.A(_20349_),
    .B(_01513_),
    .X(_01514_));
 sky130_fd_sc_hd__buf_1 _25334_ (.A(_20019_),
    .X(_20350_));
 sky130_fd_sc_hd__and2_2 _25335_ (.A(_20350_),
    .B(_01516_),
    .X(_01517_));
 sky130_fd_sc_hd__and2_2 _25336_ (.A(_20350_),
    .B(_01519_),
    .X(_01520_));
 sky130_fd_sc_hd__and2_2 _25337_ (.A(_20350_),
    .B(_01522_),
    .X(_01523_));
 sky130_fd_sc_hd__and2_2 _25338_ (.A(_20350_),
    .B(_01525_),
    .X(_01526_));
 sky130_fd_sc_hd__and2_2 _25339_ (.A(_20350_),
    .B(_01528_),
    .X(_01529_));
 sky130_fd_sc_hd__and2_2 _25340_ (.A(_20350_),
    .B(_01531_),
    .X(_01532_));
 sky130_fd_sc_hd__buf_1 _25341_ (.A(latched_branch),
    .X(_20351_));
 sky130_fd_sc_hd__and2_2 _25342_ (.A(_20351_),
    .B(_01534_),
    .X(_01535_));
 sky130_fd_sc_hd__and2_2 _25343_ (.A(_20351_),
    .B(_01537_),
    .X(_01538_));
 sky130_fd_sc_hd__and2_2 _25344_ (.A(_20351_),
    .B(_01540_),
    .X(_01541_));
 sky130_fd_sc_hd__and2_2 _25345_ (.A(_20351_),
    .B(_01543_),
    .X(_01544_));
 sky130_fd_sc_hd__and2_2 _25346_ (.A(_20351_),
    .B(_01546_),
    .X(_01547_));
 sky130_fd_sc_hd__and2_2 _25347_ (.A(_20351_),
    .B(_01549_),
    .X(_01550_));
 sky130_fd_sc_hd__and2_2 _25348_ (.A(_20019_),
    .B(_01552_),
    .X(_01553_));
 sky130_fd_sc_hd__and2_2 _25349_ (.A(_20019_),
    .B(_01555_),
    .X(_01556_));
 sky130_fd_sc_hd__nor2_2 _25350_ (.A(_02590_),
    .B(\decoded_imm_uj[1] ),
    .Y(_20352_));
 sky130_fd_sc_hd__and2_2 _25351_ (.A(_02590_),
    .B(\decoded_imm_uj[1] ),
    .X(_20353_));
 sky130_fd_sc_hd__nor2_2 _25352_ (.A(_20352_),
    .B(_20353_),
    .Y(_01557_));
 sky130_fd_sc_hd__nor2_2 _25353_ (.A(_02560_),
    .B(\decoded_imm_uj[2] ),
    .Y(_20354_));
 sky130_fd_sc_hd__and2_2 _25354_ (.A(_02560_),
    .B(\decoded_imm_uj[2] ),
    .X(_20355_));
 sky130_fd_sc_hd__nor2_2 _25355_ (.A(_20354_),
    .B(_20355_),
    .Y(_20356_));
 sky130_fd_sc_hd__xor2_2 _25356_ (.A(_20353_),
    .B(_20356_),
    .X(_01562_));
 sky130_fd_sc_hd__xor2_2 _25357_ (.A(_01561_),
    .B(_02410_),
    .X(_01565_));
 sky130_fd_sc_hd__nor2_2 _25358_ (.A(_02571_),
    .B(_02560_),
    .Y(_20357_));
 sky130_fd_sc_hd__nand2_2 _25359_ (.A(_02571_),
    .B(_02560_),
    .Y(_20358_));
 sky130_fd_sc_hd__inv_2 _25360_ (.A(_20358_),
    .Y(_20359_));
 sky130_fd_sc_hd__nor2_2 _25361_ (.A(_20357_),
    .B(_20359_),
    .Y(_01567_));
 sky130_fd_sc_hd__or2_2 _25362_ (.A(_02571_),
    .B(\decoded_imm_uj[3] ),
    .X(_20360_));
 sky130_fd_sc_hd__nand2_2 _25363_ (.A(_02571_),
    .B(\decoded_imm_uj[3] ),
    .Y(_20361_));
 sky130_fd_sc_hd__nand2_2 _25364_ (.A(_20360_),
    .B(_20361_),
    .Y(_20362_));
 sky130_fd_sc_hd__a21o_2 _25365_ (.A1(_20356_),
    .A2(_20353_),
    .B1(_20355_),
    .X(_20363_));
 sky130_fd_sc_hd__xnor2_2 _25366_ (.A(_20362_),
    .B(_20363_),
    .Y(_01568_));
 sky130_fd_sc_hd__nor2_2 _25367_ (.A(_01475_),
    .B(_20358_),
    .Y(_20364_));
 sky130_fd_sc_hd__nor2_2 _25368_ (.A(_02582_),
    .B(_20359_),
    .Y(_20365_));
 sky130_fd_sc_hd__nor2_2 _25369_ (.A(_20364_),
    .B(_20365_),
    .Y(_01571_));
 sky130_fd_sc_hd__nor2_2 _25370_ (.A(_01475_),
    .B(_00367_),
    .Y(_20366_));
 sky130_fd_sc_hd__nor2_2 _25371_ (.A(\decoded_imm_uj[4] ),
    .B(_02582_),
    .Y(_20367_));
 sky130_fd_sc_hd__nor2_2 _25372_ (.A(_20366_),
    .B(_20367_),
    .Y(_20368_));
 sky130_fd_sc_hd__nand2_2 _25373_ (.A(_20363_),
    .B(_20360_),
    .Y(_20369_));
 sky130_fd_sc_hd__nand2_2 _25374_ (.A(_20369_),
    .B(_20361_),
    .Y(_20370_));
 sky130_fd_sc_hd__xor2_2 _25375_ (.A(_20368_),
    .B(_20370_),
    .X(_01572_));
 sky130_fd_sc_hd__nor2_2 _25376_ (.A(_02583_),
    .B(_20364_),
    .Y(_20371_));
 sky130_fd_sc_hd__and2_2 _25377_ (.A(_20364_),
    .B(_02583_),
    .X(_20372_));
 sky130_fd_sc_hd__nor2_2 _25378_ (.A(_20371_),
    .B(_20372_),
    .Y(_01575_));
 sky130_fd_sc_hd__a21oi_2 _25379_ (.A1(_20369_),
    .A2(_20361_),
    .B1(_20367_),
    .Y(_20373_));
 sky130_fd_sc_hd__and2_2 _25380_ (.A(_02583_),
    .B(\decoded_imm_uj[5] ),
    .X(_20374_));
 sky130_fd_sc_hd__inv_2 _25381_ (.A(_20374_),
    .Y(_20375_));
 sky130_fd_sc_hd__nor2_2 _25382_ (.A(_02583_),
    .B(\decoded_imm_uj[5] ),
    .Y(_20376_));
 sky130_fd_sc_hd__inv_2 _25383_ (.A(_20376_),
    .Y(_20377_));
 sky130_fd_sc_hd__nand2_2 _25384_ (.A(_20375_),
    .B(_20377_),
    .Y(_20378_));
 sky130_fd_sc_hd__o21ai_2 _25385_ (.A1(_20366_),
    .A2(_20373_),
    .B1(_20378_),
    .Y(_20379_));
 sky130_fd_sc_hd__or3_2 _25386_ (.A(_20366_),
    .B(_20378_),
    .C(_20373_),
    .X(_20380_));
 sky130_fd_sc_hd__nand2_2 _25387_ (.A(_20379_),
    .B(_20380_),
    .Y(_01576_));
 sky130_fd_sc_hd__nor2_2 _25388_ (.A(_02584_),
    .B(_20372_),
    .Y(_20381_));
 sky130_fd_sc_hd__nand2_2 _25389_ (.A(_20372_),
    .B(_02584_),
    .Y(_20382_));
 sky130_fd_sc_hd__inv_2 _25390_ (.A(_20382_),
    .Y(_20383_));
 sky130_fd_sc_hd__nor2_2 _25391_ (.A(_20381_),
    .B(_20383_),
    .Y(_01579_));
 sky130_fd_sc_hd__nor2_2 _25392_ (.A(_02584_),
    .B(\decoded_imm_uj[6] ),
    .Y(_20384_));
 sky130_fd_sc_hd__nand2_2 _25393_ (.A(_02584_),
    .B(\decoded_imm_uj[6] ),
    .Y(_20385_));
 sky130_fd_sc_hd__inv_2 _25394_ (.A(_20385_),
    .Y(_20386_));
 sky130_fd_sc_hd__nor2_2 _25395_ (.A(_20384_),
    .B(_20386_),
    .Y(_20387_));
 sky130_fd_sc_hd__o21ai_2 _25396_ (.A1(_20366_),
    .A2(_20373_),
    .B1(_20377_),
    .Y(_20388_));
 sky130_fd_sc_hd__nand2_2 _25397_ (.A(_20388_),
    .B(_20375_),
    .Y(_20389_));
 sky130_fd_sc_hd__xor2_2 _25398_ (.A(_20387_),
    .B(_20389_),
    .X(_01580_));
 sky130_fd_sc_hd__nor2_2 _25399_ (.A(_18562_),
    .B(_20382_),
    .Y(_20390_));
 sky130_fd_sc_hd__nor2_2 _25400_ (.A(_02585_),
    .B(_20383_),
    .Y(_20391_));
 sky130_fd_sc_hd__nor2_2 _25401_ (.A(_20390_),
    .B(_20391_),
    .Y(_01583_));
 sky130_fd_sc_hd__or2_2 _25402_ (.A(_02585_),
    .B(\decoded_imm_uj[7] ),
    .X(_20392_));
 sky130_fd_sc_hd__nand2_2 _25403_ (.A(_02585_),
    .B(\decoded_imm_uj[7] ),
    .Y(_20393_));
 sky130_fd_sc_hd__nand2_2 _25404_ (.A(_20392_),
    .B(_20393_),
    .Y(_20394_));
 sky130_fd_sc_hd__a21oi_2 _25405_ (.A1(_20388_),
    .A2(_20375_),
    .B1(_20384_),
    .Y(_20395_));
 sky130_fd_sc_hd__nor2_2 _25406_ (.A(_20386_),
    .B(_20395_),
    .Y(_20396_));
 sky130_fd_sc_hd__xor2_2 _25407_ (.A(_20394_),
    .B(_20396_),
    .X(_01584_));
 sky130_fd_sc_hd__or2_2 _25408_ (.A(_02586_),
    .B(_20390_),
    .X(_20397_));
 sky130_fd_sc_hd__nand2_2 _25409_ (.A(_20390_),
    .B(_02586_),
    .Y(_20398_));
 sky130_fd_sc_hd__and2_2 _25410_ (.A(_20397_),
    .B(_20398_),
    .X(_01587_));
 sky130_fd_sc_hd__nor2_2 _25411_ (.A(_02586_),
    .B(\decoded_imm_uj[8] ),
    .Y(_20399_));
 sky130_fd_sc_hd__and2_2 _25412_ (.A(_02586_),
    .B(\decoded_imm_uj[8] ),
    .X(_20400_));
 sky130_fd_sc_hd__nor2_2 _25413_ (.A(_20399_),
    .B(_20400_),
    .Y(_20401_));
 sky130_fd_sc_hd__o21ai_2 _25414_ (.A1(_20386_),
    .A2(_20395_),
    .B1(_20392_),
    .Y(_20402_));
 sky130_fd_sc_hd__nand2_2 _25415_ (.A(_20402_),
    .B(_20393_),
    .Y(_20403_));
 sky130_fd_sc_hd__xor2_2 _25416_ (.A(_20401_),
    .B(_20403_),
    .X(_01588_));
 sky130_fd_sc_hd__nor2_2 _25417_ (.A(_18558_),
    .B(_20398_),
    .Y(_20404_));
 sky130_fd_sc_hd__and2_2 _25418_ (.A(_20398_),
    .B(_18558_),
    .X(_20405_));
 sky130_fd_sc_hd__nor2_2 _25419_ (.A(_20404_),
    .B(_20405_),
    .Y(_01591_));
 sky130_fd_sc_hd__or2_2 _25420_ (.A(_02587_),
    .B(\decoded_imm_uj[9] ),
    .X(_20406_));
 sky130_fd_sc_hd__nand2_2 _25421_ (.A(_02587_),
    .B(\decoded_imm_uj[9] ),
    .Y(_20407_));
 sky130_fd_sc_hd__nand2_2 _25422_ (.A(_20406_),
    .B(_20407_),
    .Y(_20408_));
 sky130_fd_sc_hd__a21oi_2 _25423_ (.A1(_20402_),
    .A2(_20393_),
    .B1(_20399_),
    .Y(_20409_));
 sky130_fd_sc_hd__nor2_2 _25424_ (.A(_20400_),
    .B(_20409_),
    .Y(_20410_));
 sky130_fd_sc_hd__xor2_2 _25425_ (.A(_20408_),
    .B(_20410_),
    .X(_01592_));
 sky130_fd_sc_hd__nor2_2 _25426_ (.A(_02588_),
    .B(_20404_),
    .Y(_20411_));
 sky130_fd_sc_hd__and2_2 _25427_ (.A(_20404_),
    .B(_02588_),
    .X(_20412_));
 sky130_fd_sc_hd__nor2_2 _25428_ (.A(_20411_),
    .B(_20412_),
    .Y(_01595_));
 sky130_fd_sc_hd__nor2_2 _25429_ (.A(_02588_),
    .B(\decoded_imm_uj[10] ),
    .Y(_20413_));
 sky130_fd_sc_hd__and2_2 _25430_ (.A(_02588_),
    .B(\decoded_imm_uj[10] ),
    .X(_20414_));
 sky130_fd_sc_hd__nor2_2 _25431_ (.A(_20413_),
    .B(_20414_),
    .Y(_20415_));
 sky130_fd_sc_hd__o21ai_2 _25432_ (.A1(_20400_),
    .A2(_20409_),
    .B1(_20406_),
    .Y(_20416_));
 sky130_fd_sc_hd__nand2_2 _25433_ (.A(_20416_),
    .B(_20407_),
    .Y(_20417_));
 sky130_fd_sc_hd__xor2_2 _25434_ (.A(_20415_),
    .B(_20417_),
    .X(_01596_));
 sky130_fd_sc_hd__or2_2 _25435_ (.A(_02589_),
    .B(_20412_),
    .X(_20418_));
 sky130_fd_sc_hd__nand2_2 _25436_ (.A(_20412_),
    .B(_02589_),
    .Y(_20419_));
 sky130_fd_sc_hd__and2_2 _25437_ (.A(_20418_),
    .B(_20419_),
    .X(_01599_));
 sky130_fd_sc_hd__a21oi_2 _25438_ (.A1(_20416_),
    .A2(_20407_),
    .B1(_20413_),
    .Y(_20420_));
 sky130_fd_sc_hd__nor2_2 _25439_ (.A(_20414_),
    .B(_20420_),
    .Y(_20421_));
 sky130_fd_sc_hd__nor2_2 _25440_ (.A(_02589_),
    .B(\decoded_imm_uj[11] ),
    .Y(_20422_));
 sky130_fd_sc_hd__nand2_2 _25441_ (.A(_02589_),
    .B(\decoded_imm_uj[11] ),
    .Y(_20423_));
 sky130_fd_sc_hd__inv_2 _25442_ (.A(_20423_),
    .Y(_20424_));
 sky130_fd_sc_hd__or2_2 _25443_ (.A(_20422_),
    .B(_20424_),
    .X(_20425_));
 sky130_fd_sc_hd__nand2_2 _25444_ (.A(_20421_),
    .B(_20425_),
    .Y(_20426_));
 sky130_fd_sc_hd__o21bai_2 _25445_ (.A1(_20414_),
    .A2(_20420_),
    .B1_N(_20425_),
    .Y(_20427_));
 sky130_fd_sc_hd__and2_2 _25446_ (.A(_20426_),
    .B(_20427_),
    .X(_01600_));
 sky130_fd_sc_hd__nor2_2 _25447_ (.A(_18550_),
    .B(_20419_),
    .Y(_20428_));
 sky130_fd_sc_hd__and2_2 _25448_ (.A(_20419_),
    .B(_18550_),
    .X(_20429_));
 sky130_fd_sc_hd__nor2_2 _25449_ (.A(_20428_),
    .B(_20429_),
    .Y(_01603_));
 sky130_fd_sc_hd__nor2_2 _25450_ (.A(_02561_),
    .B(\decoded_imm_uj[12] ),
    .Y(_20430_));
 sky130_fd_sc_hd__and2_2 _25451_ (.A(_02561_),
    .B(\decoded_imm_uj[12] ),
    .X(_20431_));
 sky130_fd_sc_hd__or2_2 _25452_ (.A(_20430_),
    .B(_20431_),
    .X(_20432_));
 sky130_fd_sc_hd__a21oi_2 _25453_ (.A1(_20427_),
    .A2(_20423_),
    .B1(_20432_),
    .Y(_20433_));
 sky130_fd_sc_hd__and3_2 _25454_ (.A(_20427_),
    .B(_20423_),
    .C(_20432_),
    .X(_20434_));
 sky130_fd_sc_hd__nor2_2 _25455_ (.A(_20433_),
    .B(_20434_),
    .Y(_01604_));
 sky130_fd_sc_hd__or2_2 _25456_ (.A(_02562_),
    .B(_20428_),
    .X(_20435_));
 sky130_fd_sc_hd__nand2_2 _25457_ (.A(_20428_),
    .B(_02562_),
    .Y(_20436_));
 sky130_fd_sc_hd__and2_2 _25458_ (.A(_20435_),
    .B(_20436_),
    .X(_01607_));
 sky130_fd_sc_hd__inv_2 _25459_ (.A(\decoded_imm_uj[13] ),
    .Y(_20437_));
 sky130_fd_sc_hd__nor2_2 _25460_ (.A(_02562_),
    .B(_20437_),
    .Y(_20438_));
 sky130_fd_sc_hd__nor2_2 _25461_ (.A(\decoded_imm_uj[13] ),
    .B(_18548_),
    .Y(_20439_));
 sky130_fd_sc_hd__or4_2 _25462_ (.A(_20431_),
    .B(_20438_),
    .C(_20439_),
    .D(_20433_),
    .X(_20440_));
 sky130_fd_sc_hd__nor2_2 _25463_ (.A(_20438_),
    .B(_20439_),
    .Y(_20441_));
 sky130_fd_sc_hd__o21bai_2 _25464_ (.A1(_20431_),
    .A2(_20433_),
    .B1_N(_20441_),
    .Y(_20442_));
 sky130_fd_sc_hd__and2_2 _25465_ (.A(_20440_),
    .B(_20442_),
    .X(_01608_));
 sky130_fd_sc_hd__nor2_2 _25466_ (.A(_18545_),
    .B(_20436_),
    .Y(_20443_));
 sky130_fd_sc_hd__and2_2 _25467_ (.A(_20436_),
    .B(_18545_),
    .X(_20444_));
 sky130_fd_sc_hd__nor2_2 _25468_ (.A(_20443_),
    .B(_20444_),
    .Y(_01611_));
 sky130_fd_sc_hd__nor2_2 _25469_ (.A(_18548_),
    .B(_20437_),
    .Y(_20445_));
 sky130_fd_sc_hd__inv_2 _25470_ (.A(_20445_),
    .Y(_20446_));
 sky130_fd_sc_hd__nor2_2 _25471_ (.A(_02563_),
    .B(\decoded_imm_uj[14] ),
    .Y(_20447_));
 sky130_fd_sc_hd__and2_2 _25472_ (.A(_02563_),
    .B(\decoded_imm_uj[14] ),
    .X(_20448_));
 sky130_fd_sc_hd__or2_2 _25473_ (.A(_20447_),
    .B(_20448_),
    .X(_20449_));
 sky130_fd_sc_hd__a21oi_2 _25474_ (.A1(_20442_),
    .A2(_20446_),
    .B1(_20449_),
    .Y(_20450_));
 sky130_fd_sc_hd__and3_2 _25475_ (.A(_20442_),
    .B(_20446_),
    .C(_20449_),
    .X(_20451_));
 sky130_fd_sc_hd__nor2_2 _25476_ (.A(_20450_),
    .B(_20451_),
    .Y(_01612_));
 sky130_fd_sc_hd__nor2_2 _25477_ (.A(_02564_),
    .B(_20443_),
    .Y(_20452_));
 sky130_fd_sc_hd__nand2_2 _25478_ (.A(_20443_),
    .B(_02564_),
    .Y(_20453_));
 sky130_fd_sc_hd__inv_2 _25479_ (.A(_20453_),
    .Y(_20454_));
 sky130_fd_sc_hd__nor2_2 _25480_ (.A(_20452_),
    .B(_20454_),
    .Y(_01615_));
 sky130_fd_sc_hd__nor2_2 _25481_ (.A(_02564_),
    .B(_19430_),
    .Y(_20455_));
 sky130_fd_sc_hd__nor2_2 _25482_ (.A(\decoded_imm_uj[15] ),
    .B(_18543_),
    .Y(_20456_));
 sky130_fd_sc_hd__or4_2 _25483_ (.A(_20448_),
    .B(_20455_),
    .C(_20456_),
    .D(_20450_),
    .X(_20457_));
 sky130_fd_sc_hd__nor2_2 _25484_ (.A(_20455_),
    .B(_20456_),
    .Y(_20458_));
 sky130_fd_sc_hd__o21bai_2 _25485_ (.A1(_20448_),
    .A2(_20450_),
    .B1_N(_20458_),
    .Y(_20459_));
 sky130_fd_sc_hd__and2_2 _25486_ (.A(_20457_),
    .B(_20459_),
    .X(_01616_));
 sky130_fd_sc_hd__nor2_2 _25487_ (.A(_18540_),
    .B(_20453_),
    .Y(_20460_));
 sky130_fd_sc_hd__nor2_2 _25488_ (.A(_02565_),
    .B(_20454_),
    .Y(_20461_));
 sky130_fd_sc_hd__nor2_2 _25489_ (.A(_20460_),
    .B(_20461_),
    .Y(_01619_));
 sky130_fd_sc_hd__nor2_2 _25490_ (.A(_18543_),
    .B(_19430_),
    .Y(_20462_));
 sky130_fd_sc_hd__inv_2 _25491_ (.A(_20462_),
    .Y(_20463_));
 sky130_fd_sc_hd__nor2_2 _25492_ (.A(_02565_),
    .B(\decoded_imm_uj[16] ),
    .Y(_20464_));
 sky130_fd_sc_hd__nor2_2 _25493_ (.A(_18540_),
    .B(_19429_),
    .Y(_20465_));
 sky130_fd_sc_hd__nor2_2 _25494_ (.A(_20464_),
    .B(_20465_),
    .Y(_20466_));
 sky130_fd_sc_hd__inv_2 _25495_ (.A(_20466_),
    .Y(_20467_));
 sky130_fd_sc_hd__a21oi_2 _25496_ (.A1(_20459_),
    .A2(_20463_),
    .B1(_20467_),
    .Y(_20468_));
 sky130_fd_sc_hd__and3_2 _25497_ (.A(_20459_),
    .B(_20463_),
    .C(_20467_),
    .X(_20469_));
 sky130_fd_sc_hd__nor2_2 _25498_ (.A(_20468_),
    .B(_20469_),
    .Y(_01620_));
 sky130_fd_sc_hd__nor2_2 _25499_ (.A(_02566_),
    .B(_20460_),
    .Y(_20470_));
 sky130_fd_sc_hd__nand2_2 _25500_ (.A(_20460_),
    .B(_02566_),
    .Y(_20471_));
 sky130_fd_sc_hd__inv_2 _25501_ (.A(_20471_),
    .Y(_20472_));
 sky130_fd_sc_hd__nor2_2 _25502_ (.A(_20470_),
    .B(_20472_),
    .Y(_01623_));
 sky130_fd_sc_hd__nor2_2 _25503_ (.A(_02566_),
    .B(\decoded_imm_uj[17] ),
    .Y(_20473_));
 sky130_fd_sc_hd__nor2_2 _25504_ (.A(_18537_),
    .B(_19428_),
    .Y(_20474_));
 sky130_fd_sc_hd__or2_2 _25505_ (.A(_20473_),
    .B(_20474_),
    .X(_20475_));
 sky130_fd_sc_hd__or3b_2 _25506_ (.A(_20465_),
    .B(_20468_),
    .C_N(_20475_),
    .X(_20476_));
 sky130_fd_sc_hd__o21bai_2 _25507_ (.A1(_20465_),
    .A2(_20468_),
    .B1_N(_20475_),
    .Y(_20477_));
 sky130_fd_sc_hd__and2_2 _25508_ (.A(_20476_),
    .B(_20477_),
    .X(_01624_));
 sky130_fd_sc_hd__nor2_2 _25509_ (.A(_18535_),
    .B(_20471_),
    .Y(_20478_));
 sky130_fd_sc_hd__nor2_2 _25510_ (.A(_02567_),
    .B(_20472_),
    .Y(_20479_));
 sky130_fd_sc_hd__nor2_2 _25511_ (.A(_20478_),
    .B(_20479_),
    .Y(_01627_));
 sky130_fd_sc_hd__nor2_2 _25512_ (.A(_02567_),
    .B(\decoded_imm_uj[18] ),
    .Y(_20480_));
 sky130_fd_sc_hd__nor2_2 _25513_ (.A(_18535_),
    .B(_19427_),
    .Y(_20481_));
 sky130_fd_sc_hd__nor2_2 _25514_ (.A(_20480_),
    .B(_20481_),
    .Y(_20482_));
 sky130_fd_sc_hd__inv_2 _25515_ (.A(_20474_),
    .Y(_20483_));
 sky130_fd_sc_hd__nand2_2 _25516_ (.A(_20477_),
    .B(_20483_),
    .Y(_20484_));
 sky130_fd_sc_hd__xor2_2 _25517_ (.A(_20482_),
    .B(_20484_),
    .X(_01628_));
 sky130_fd_sc_hd__nor2_2 _25518_ (.A(_02568_),
    .B(_20478_),
    .Y(_20485_));
 sky130_fd_sc_hd__nand2_2 _25519_ (.A(_20478_),
    .B(_02568_),
    .Y(_20486_));
 sky130_fd_sc_hd__inv_2 _25520_ (.A(_20486_),
    .Y(_20487_));
 sky130_fd_sc_hd__nor2_2 _25521_ (.A(_20485_),
    .B(_20487_),
    .Y(_01631_));
 sky130_fd_sc_hd__a21oi_2 _25522_ (.A1(_20477_),
    .A2(_20483_),
    .B1(_20480_),
    .Y(_20488_));
 sky130_fd_sc_hd__nor2_2 _25523_ (.A(_02568_),
    .B(\decoded_imm_uj[19] ),
    .Y(_20489_));
 sky130_fd_sc_hd__inv_2 _25524_ (.A(\decoded_imm_uj[19] ),
    .Y(_20490_));
 sky130_fd_sc_hd__nor2_2 _25525_ (.A(_18533_),
    .B(_20490_),
    .Y(_20491_));
 sky130_fd_sc_hd__or2_2 _25526_ (.A(_20489_),
    .B(_20491_),
    .X(_20492_));
 sky130_fd_sc_hd__or3b_2 _25527_ (.A(_20481_),
    .B(_20488_),
    .C_N(_20492_),
    .X(_20493_));
 sky130_fd_sc_hd__o21bai_2 _25528_ (.A1(_20481_),
    .A2(_20488_),
    .B1_N(_20492_),
    .Y(_20494_));
 sky130_fd_sc_hd__and2_2 _25529_ (.A(_20493_),
    .B(_20494_),
    .X(_01632_));
 sky130_fd_sc_hd__nor2_2 _25530_ (.A(_18530_),
    .B(_20486_),
    .Y(_20495_));
 sky130_fd_sc_hd__nor2_2 _25531_ (.A(_02569_),
    .B(_20487_),
    .Y(_20496_));
 sky130_fd_sc_hd__nor2_2 _25532_ (.A(_20495_),
    .B(_20496_),
    .Y(_01635_));
 sky130_fd_sc_hd__inv_2 _25533_ (.A(_20491_),
    .Y(_20497_));
 sky130_fd_sc_hd__nor2_2 _25534_ (.A(_02569_),
    .B(_19424_),
    .Y(_20498_));
 sky130_fd_sc_hd__inv_2 _25535_ (.A(\decoded_imm_uj[20] ),
    .Y(_20499_));
 sky130_fd_sc_hd__nor2_2 _25536_ (.A(_18530_),
    .B(_20499_),
    .Y(_20500_));
 sky130_fd_sc_hd__or2_2 _25537_ (.A(_20498_),
    .B(_20500_),
    .X(_20501_));
 sky130_fd_sc_hd__a21oi_2 _25538_ (.A1(_20494_),
    .A2(_20497_),
    .B1(_20501_),
    .Y(_20502_));
 sky130_fd_sc_hd__and3_2 _25539_ (.A(_20494_),
    .B(_20497_),
    .C(_20501_),
    .X(_20503_));
 sky130_fd_sc_hd__nor2_2 _25540_ (.A(_20502_),
    .B(_20503_),
    .Y(_01636_));
 sky130_fd_sc_hd__nor2_2 _25541_ (.A(_02570_),
    .B(_20495_),
    .Y(_20504_));
 sky130_fd_sc_hd__and2_2 _25542_ (.A(_20495_),
    .B(_02570_),
    .X(_20505_));
 sky130_fd_sc_hd__nor2_2 _25543_ (.A(_20504_),
    .B(_20505_),
    .Y(_01639_));
 sky130_fd_sc_hd__nor2_2 _25544_ (.A(_02570_),
    .B(\decoded_imm_uj[20] ),
    .Y(_20506_));
 sky130_fd_sc_hd__nor2_2 _25545_ (.A(_18528_),
    .B(_20499_),
    .Y(_20507_));
 sky130_fd_sc_hd__or2_2 _25546_ (.A(_20506_),
    .B(_20507_),
    .X(_20508_));
 sky130_fd_sc_hd__inv_2 _25547_ (.A(_20508_),
    .Y(_20509_));
 sky130_fd_sc_hd__a21oi_2 _25548_ (.A1(_20494_),
    .A2(_20497_),
    .B1(_20498_),
    .Y(_20510_));
 sky130_fd_sc_hd__or2_2 _25549_ (.A(_20500_),
    .B(_20510_),
    .X(_20511_));
 sky130_fd_sc_hd__or2_2 _25550_ (.A(_20509_),
    .B(_20511_),
    .X(_20512_));
 sky130_fd_sc_hd__nand2_2 _25551_ (.A(_20511_),
    .B(_20509_),
    .Y(_20513_));
 sky130_fd_sc_hd__and2_2 _25552_ (.A(_20512_),
    .B(_20513_),
    .X(_01640_));
 sky130_fd_sc_hd__nor2_2 _25553_ (.A(_02572_),
    .B(_20505_),
    .Y(_20514_));
 sky130_fd_sc_hd__nand2_2 _25554_ (.A(_20505_),
    .B(_02572_),
    .Y(_20515_));
 sky130_fd_sc_hd__inv_2 _25555_ (.A(_20515_),
    .Y(_20516_));
 sky130_fd_sc_hd__nor2_2 _25556_ (.A(_20514_),
    .B(_20516_),
    .Y(_01643_));
 sky130_fd_sc_hd__xnor2_2 _25557_ (.A(_02572_),
    .B(\decoded_imm_uj[20] ),
    .Y(_20517_));
 sky130_fd_sc_hd__a21oi_2 _25558_ (.A1(_20511_),
    .A2(_20509_),
    .B1(_20507_),
    .Y(_20518_));
 sky130_fd_sc_hd__xor2_2 _25559_ (.A(_20517_),
    .B(_20518_),
    .X(_01644_));
 sky130_fd_sc_hd__nor2_2 _25560_ (.A(_18522_),
    .B(_20515_),
    .Y(_20519_));
 sky130_fd_sc_hd__nor2_2 _25561_ (.A(_02573_),
    .B(_20516_),
    .Y(_20520_));
 sky130_fd_sc_hd__nor2_2 _25562_ (.A(_20519_),
    .B(_20520_),
    .Y(_01647_));
 sky130_fd_sc_hd__nor2_2 _25563_ (.A(_20517_),
    .B(_20513_),
    .Y(_20521_));
 sky130_fd_sc_hd__nor2_2 _25564_ (.A(_18522_),
    .B(_20499_),
    .Y(_20522_));
 sky130_fd_sc_hd__inv_2 _25565_ (.A(_20522_),
    .Y(_20523_));
 sky130_fd_sc_hd__nand2_2 _25566_ (.A(_18522_),
    .B(_20499_),
    .Y(_20524_));
 sky130_fd_sc_hd__o21a_2 _25567_ (.A1(_02572_),
    .A2(_02570_),
    .B1(_19425_),
    .X(_20525_));
 sky130_fd_sc_hd__a21o_2 _25568_ (.A1(_20523_),
    .A2(_20524_),
    .B1(_20525_),
    .X(_20526_));
 sky130_fd_sc_hd__nand2_2 _25569_ (.A(_20523_),
    .B(_20524_),
    .Y(_20527_));
 sky130_fd_sc_hd__o21bai_2 _25570_ (.A1(_20525_),
    .A2(_20521_),
    .B1_N(_20527_),
    .Y(_20528_));
 sky130_fd_sc_hd__o21a_2 _25571_ (.A1(_20521_),
    .A2(_20526_),
    .B1(_20528_),
    .X(_01648_));
 sky130_fd_sc_hd__nor2_2 _25572_ (.A(_02574_),
    .B(_20519_),
    .Y(_20529_));
 sky130_fd_sc_hd__and2_2 _25573_ (.A(_20519_),
    .B(_02574_),
    .X(_20530_));
 sky130_fd_sc_hd__nor2_2 _25574_ (.A(_20529_),
    .B(_20530_),
    .Y(_01651_));
 sky130_fd_sc_hd__xnor2_2 _25575_ (.A(_02574_),
    .B(\decoded_imm_uj[20] ),
    .Y(_20531_));
 sky130_fd_sc_hd__a21oi_2 _25576_ (.A1(_20528_),
    .A2(_20523_),
    .B1(_20531_),
    .Y(_20532_));
 sky130_fd_sc_hd__and3_2 _25577_ (.A(_20528_),
    .B(_20523_),
    .C(_20531_),
    .X(_20533_));
 sky130_fd_sc_hd__nor2_2 _25578_ (.A(_20532_),
    .B(_20533_),
    .Y(_01652_));
 sky130_fd_sc_hd__or2_2 _25579_ (.A(_02575_),
    .B(_20530_),
    .X(_20534_));
 sky130_fd_sc_hd__nand2_2 _25580_ (.A(_20530_),
    .B(_02575_),
    .Y(_20535_));
 sky130_fd_sc_hd__and2_2 _25581_ (.A(_20534_),
    .B(_20535_),
    .X(_01655_));
 sky130_fd_sc_hd__buf_1 _25582_ (.A(_20499_),
    .X(_20536_));
 sky130_fd_sc_hd__nor2_2 _25583_ (.A(_02575_),
    .B(_20536_),
    .Y(_20537_));
 sky130_fd_sc_hd__nor2_2 _25584_ (.A(_19425_),
    .B(_18518_),
    .Y(_20538_));
 sky130_fd_sc_hd__or2_2 _25585_ (.A(_20537_),
    .B(_20538_),
    .X(_20539_));
 sky130_fd_sc_hd__inv_2 _25586_ (.A(_20517_),
    .Y(_20540_));
 sky130_fd_sc_hd__nor2_2 _25587_ (.A(_20531_),
    .B(_20527_),
    .Y(_20541_));
 sky130_fd_sc_hd__o2111ai_2 _25588_ (.A1(_20500_),
    .A2(_20510_),
    .B1(_20509_),
    .C1(_20540_),
    .D1(_20541_),
    .Y(_20542_));
 sky130_fd_sc_hd__a41o_2 _25589_ (.A1(_18520_),
    .A2(_18522_),
    .A3(_18525_),
    .A4(_18528_),
    .B1(_20536_),
    .X(_20543_));
 sky130_fd_sc_hd__nand2_2 _25590_ (.A(_20542_),
    .B(_20543_),
    .Y(_20544_));
 sky130_fd_sc_hd__or2_2 _25591_ (.A(_20539_),
    .B(_20544_),
    .X(_20545_));
 sky130_fd_sc_hd__nand2_2 _25592_ (.A(_20544_),
    .B(_20539_),
    .Y(_20546_));
 sky130_fd_sc_hd__and2_2 _25593_ (.A(_20545_),
    .B(_20546_),
    .X(_01656_));
 sky130_fd_sc_hd__nor2_2 _25594_ (.A(_18515_),
    .B(_20535_),
    .Y(_20547_));
 sky130_fd_sc_hd__and2_2 _25595_ (.A(_20535_),
    .B(_18515_),
    .X(_20548_));
 sky130_fd_sc_hd__nor2_2 _25596_ (.A(_20547_),
    .B(_20548_),
    .Y(_01659_));
 sky130_fd_sc_hd__nor2_2 _25597_ (.A(_02576_),
    .B(_19424_),
    .Y(_20549_));
 sky130_fd_sc_hd__nor2_2 _25598_ (.A(_18515_),
    .B(_20536_),
    .Y(_20550_));
 sky130_fd_sc_hd__nor2_2 _25599_ (.A(_20549_),
    .B(_20550_),
    .Y(_20551_));
 sky130_fd_sc_hd__nor2_2 _25600_ (.A(_18518_),
    .B(_20536_),
    .Y(_20552_));
 sky130_fd_sc_hd__a21oi_2 _25601_ (.A1(_20544_),
    .A2(_20539_),
    .B1(_20552_),
    .Y(_20553_));
 sky130_fd_sc_hd__xnor2_2 _25602_ (.A(_20551_),
    .B(_20553_),
    .Y(_01660_));
 sky130_fd_sc_hd__nor2_2 _25603_ (.A(_02577_),
    .B(_20547_),
    .Y(_20554_));
 sky130_fd_sc_hd__nand2_2 _25604_ (.A(_20547_),
    .B(_02577_),
    .Y(_20555_));
 sky130_fd_sc_hd__inv_2 _25605_ (.A(_20555_),
    .Y(_20556_));
 sky130_fd_sc_hd__nor2_2 _25606_ (.A(_20554_),
    .B(_20556_),
    .Y(_01663_));
 sky130_fd_sc_hd__nand3_2 _25607_ (.A(_20544_),
    .B(_20539_),
    .C(_20551_),
    .Y(_20557_));
 sky130_fd_sc_hd__nor2_2 _25608_ (.A(_20552_),
    .B(_20550_),
    .Y(_20558_));
 sky130_fd_sc_hd__nor2_2 _25609_ (.A(_02577_),
    .B(_19424_),
    .Y(_20559_));
 sky130_fd_sc_hd__nor2_2 _25610_ (.A(_18513_),
    .B(_20499_),
    .Y(_20560_));
 sky130_fd_sc_hd__or2_2 _25611_ (.A(_20559_),
    .B(_20560_),
    .X(_20561_));
 sky130_fd_sc_hd__a21oi_2 _25612_ (.A1(_20557_),
    .A2(_20558_),
    .B1(_20561_),
    .Y(_20562_));
 sky130_fd_sc_hd__and3_2 _25613_ (.A(_20557_),
    .B(_20561_),
    .C(_20558_),
    .X(_20563_));
 sky130_fd_sc_hd__nor2_2 _25614_ (.A(_20562_),
    .B(_20563_),
    .Y(_01664_));
 sky130_fd_sc_hd__nor2_2 _25615_ (.A(_18510_),
    .B(_20555_),
    .Y(_20564_));
 sky130_fd_sc_hd__nor2_2 _25616_ (.A(_02578_),
    .B(_20556_),
    .Y(_20565_));
 sky130_fd_sc_hd__nor2_2 _25617_ (.A(_20564_),
    .B(_20565_),
    .Y(_01667_));
 sky130_fd_sc_hd__xnor2_2 _25618_ (.A(_02578_),
    .B(_19424_),
    .Y(_20566_));
 sky130_fd_sc_hd__a211o_2 _25619_ (.A1(_02577_),
    .A2(_19426_),
    .B1(_20566_),
    .C1(_20562_),
    .X(_20567_));
 sky130_fd_sc_hd__o21ai_2 _25620_ (.A1(_20560_),
    .A2(_20562_),
    .B1(_20566_),
    .Y(_20568_));
 sky130_fd_sc_hd__nand2_2 _25621_ (.A(_20567_),
    .B(_20568_),
    .Y(_01668_));
 sky130_fd_sc_hd__nor2_2 _25622_ (.A(_02579_),
    .B(_20564_),
    .Y(_20569_));
 sky130_fd_sc_hd__and2_2 _25623_ (.A(_20564_),
    .B(_02579_),
    .X(_20570_));
 sky130_fd_sc_hd__nor2_2 _25624_ (.A(_20569_),
    .B(_20570_),
    .Y(_01671_));
 sky130_fd_sc_hd__nor2_2 _25625_ (.A(_02579_),
    .B(_20536_),
    .Y(_20571_));
 sky130_fd_sc_hd__nor2_2 _25626_ (.A(_19424_),
    .B(_18507_),
    .Y(_20572_));
 sky130_fd_sc_hd__nor2_2 _25627_ (.A(_20571_),
    .B(_20572_),
    .Y(_20573_));
 sky130_fd_sc_hd__inv_2 _25628_ (.A(_20573_),
    .Y(_20574_));
 sky130_fd_sc_hd__nor2_2 _25629_ (.A(_20566_),
    .B(_20561_),
    .Y(_20575_));
 sky130_fd_sc_hd__o2111ai_2 _25630_ (.A1(_20537_),
    .A2(_20538_),
    .B1(_20551_),
    .C1(_20575_),
    .D1(_20544_),
    .Y(_20576_));
 sky130_fd_sc_hd__a41o_2 _25631_ (.A1(_18510_),
    .A2(_18513_),
    .A3(_18515_),
    .A4(_18518_),
    .B1(_20536_),
    .X(_20577_));
 sky130_fd_sc_hd__nand2_2 _25632_ (.A(_20576_),
    .B(_20577_),
    .Y(_20578_));
 sky130_fd_sc_hd__or2_2 _25633_ (.A(_20574_),
    .B(_20578_),
    .X(_20579_));
 sky130_fd_sc_hd__nand2_2 _25634_ (.A(_20578_),
    .B(_20574_),
    .Y(_20580_));
 sky130_fd_sc_hd__and2_2 _25635_ (.A(_20579_),
    .B(_20580_),
    .X(_01672_));
 sky130_fd_sc_hd__or2_2 _25636_ (.A(_02580_),
    .B(_20570_),
    .X(_20581_));
 sky130_fd_sc_hd__nand2_2 _25637_ (.A(_20570_),
    .B(_02580_),
    .Y(_04073_));
 sky130_fd_sc_hd__and2_2 _25638_ (.A(_20581_),
    .B(_04073_),
    .X(_01675_));
 sky130_fd_sc_hd__nand2_2 _25639_ (.A(_02579_),
    .B(_19426_),
    .Y(_04074_));
 sky130_fd_sc_hd__xor2_2 _25640_ (.A(_02580_),
    .B(_19426_),
    .X(_04075_));
 sky130_fd_sc_hd__a21o_2 _25641_ (.A1(_20580_),
    .A2(_04074_),
    .B1(_04075_),
    .X(_04076_));
 sky130_fd_sc_hd__nand3_2 _25642_ (.A(_20580_),
    .B(_04075_),
    .C(_04074_),
    .Y(_04077_));
 sky130_fd_sc_hd__nand2_2 _25643_ (.A(_04076_),
    .B(_04077_),
    .Y(_01676_));
 sky130_fd_sc_hd__xor2_2 _25644_ (.A(_18502_),
    .B(_04073_),
    .X(_01679_));
 sky130_fd_sc_hd__o21a_2 _25645_ (.A1(_02580_),
    .A2(_02579_),
    .B1(_19426_),
    .X(_04078_));
 sky130_fd_sc_hd__xor2_2 _25646_ (.A(_02581_),
    .B(_19425_),
    .X(_04079_));
 sky130_fd_sc_hd__o21a_2 _25647_ (.A1(_02580_),
    .A2(_19425_),
    .B1(_20574_),
    .X(_04080_));
 sky130_fd_sc_hd__a21boi_2 _25648_ (.A1(_20576_),
    .A2(_20577_),
    .B1_N(_04080_),
    .Y(_04081_));
 sky130_fd_sc_hd__nor3_2 _25649_ (.A(_04078_),
    .B(_04079_),
    .C(_04081_),
    .Y(_04082_));
 sky130_fd_sc_hd__o21a_2 _25650_ (.A1(_04078_),
    .A2(_04081_),
    .B1(_04079_),
    .X(_04083_));
 sky130_fd_sc_hd__nor2_2 _25651_ (.A(_04082_),
    .B(_04083_),
    .Y(_01680_));
 sky130_fd_sc_hd__nor2_2 _25652_ (.A(\mem_wordsize[2] ),
    .B(\mem_wordsize[1] ),
    .Y(_04084_));
 sky130_fd_sc_hd__buf_1 _25653_ (.A(_04084_),
    .X(_04085_));
 sky130_fd_sc_hd__buf_1 _25654_ (.A(_04085_),
    .X(_01683_));
 sky130_fd_sc_hd__buf_1 _25655_ (.A(\mem_wordsize[2] ),
    .X(_04086_));
 sky130_fd_sc_hd__a21oi_2 _25656_ (.A1(_19867_),
    .A2(_04086_),
    .B1(_04084_),
    .Y(_04087_));
 sky130_fd_sc_hd__o21ai_2 _25657_ (.A1(_19534_),
    .A2(_19535_),
    .B1(_04087_),
    .Y(mem_la_wstrb[0]));
 sky130_fd_sc_hd__and2_2 _25658_ (.A(mem_la_wstrb[0]),
    .B(mem_la_write),
    .X(_01684_));
 sky130_fd_sc_hd__and3_2 _25659_ (.A(_00301_),
    .B(_20016_),
    .C(_01685_),
    .X(_01686_));
 sky130_fd_sc_hd__o21ai_2 _25660_ (.A1(_19534_),
    .A2(_19790_),
    .B1(_04087_),
    .Y(mem_la_wstrb[1]));
 sky130_fd_sc_hd__and2_2 _25661_ (.A(mem_la_wstrb[1]),
    .B(mem_la_write),
    .X(_01687_));
 sky130_fd_sc_hd__and3_2 _25662_ (.A(_00301_),
    .B(_20016_),
    .C(_01688_),
    .X(_01689_));
 sky130_fd_sc_hd__nor2_2 _25663_ (.A(_19535_),
    .B(_19867_),
    .Y(_04088_));
 sky130_fd_sc_hd__nor2_2 _25664_ (.A(_19867_),
    .B(_19796_),
    .Y(_04089_));
 sky130_fd_sc_hd__or3_2 _25665_ (.A(_04085_),
    .B(_04088_),
    .C(_04089_),
    .X(mem_la_wstrb[2]));
 sky130_fd_sc_hd__and2_2 _25666_ (.A(mem_la_wstrb[2]),
    .B(mem_la_write),
    .X(_01690_));
 sky130_fd_sc_hd__and3_2 _25667_ (.A(_00301_),
    .B(_20016_),
    .C(_01691_),
    .X(_01692_));
 sky130_fd_sc_hd__nor2_2 _25668_ (.A(_19867_),
    .B(_19789_),
    .Y(_04090_));
 sky130_fd_sc_hd__or3_2 _25669_ (.A(_04085_),
    .B(_04089_),
    .C(_04090_),
    .X(mem_la_wstrb[3]));
 sky130_fd_sc_hd__and2_2 _25670_ (.A(mem_la_wstrb[3]),
    .B(mem_la_write),
    .X(_01693_));
 sky130_fd_sc_hd__and3_2 _25671_ (.A(_00301_),
    .B(_20016_),
    .C(_01694_),
    .X(_01695_));
 sky130_fd_sc_hd__nor2_2 _25672_ (.A(\irq_pending[1] ),
    .B(irq[1]),
    .Y(_01696_));
 sky130_fd_sc_hd__inv_2 _25673_ (.A(_01696_),
    .Y(_01697_));
 sky130_fd_sc_hd__nor2_2 _25674_ (.A(_18327_),
    .B(_01696_),
    .Y(_01698_));
 sky130_fd_sc_hd__or3_2 _25675_ (.A(\cpu_state[0] ),
    .B(_02542_),
    .C(_18255_),
    .X(_04091_));
 sky130_fd_sc_hd__nor2_2 _25676_ (.A(_19852_),
    .B(_04091_),
    .Y(_01700_));
 sky130_fd_sc_hd__nor2_2 _25677_ (.A(_19799_),
    .B(_01697_),
    .Y(_01701_));
 sky130_fd_sc_hd__a2bb2o_2 _25678_ (.A1_N(_18227_),
    .A2_N(_01704_),
    .B1(_01697_),
    .B2(_04091_),
    .X(_01705_));
 sky130_fd_sc_hd__inv_2 _25679_ (.A(mem_rdata[0]),
    .Y(_01707_));
 sky130_fd_sc_hd__nor2_2 _25680_ (.A(_19534_),
    .B(_19790_),
    .Y(_04092_));
 sky130_fd_sc_hd__buf_1 _25681_ (.A(_04092_),
    .X(_04093_));
 sky130_fd_sc_hd__buf_1 _25682_ (.A(_04088_),
    .X(_04094_));
 sky130_fd_sc_hd__buf_1 _25683_ (.A(_04090_),
    .X(_04095_));
 sky130_fd_sc_hd__a22o_2 _25684_ (.A1(_04094_),
    .A2(mem_rdata[16]),
    .B1(_04095_),
    .B2(mem_rdata[24]),
    .X(_04096_));
 sky130_fd_sc_hd__a21oi_2 _25685_ (.A1(mem_rdata[8]),
    .A2(_04093_),
    .B1(_04096_),
    .Y(_01708_));
 sky130_fd_sc_hd__buf_1 _25686_ (.A(_04086_),
    .X(_04097_));
 sky130_fd_sc_hd__o2bb2a_2 _25687_ (.A1_N(_04097_),
    .A2_N(_01710_),
    .B1(_01709_),
    .B2(_20015_),
    .X(_01711_));
 sky130_fd_sc_hd__inv_2 _25688_ (.A(instr_rdinstrh),
    .Y(_04098_));
 sky130_fd_sc_hd__buf_1 _25689_ (.A(_04098_),
    .X(_04099_));
 sky130_fd_sc_hd__inv_2 _25690_ (.A(instr_rdinstr),
    .Y(_04100_));
 sky130_fd_sc_hd__buf_1 _25691_ (.A(_04100_),
    .X(_04101_));
 sky130_fd_sc_hd__inv_2 _25692_ (.A(instr_rdcycleh),
    .Y(_04102_));
 sky130_fd_sc_hd__buf_1 _25693_ (.A(_04102_),
    .X(_04103_));
 sky130_fd_sc_hd__and3_2 _25694_ (.A(_04099_),
    .B(_04101_),
    .C(_04103_),
    .X(_01714_));
 sky130_fd_sc_hd__buf_1 _25695_ (.A(_04100_),
    .X(_04104_));
 sky130_fd_sc_hd__nand2_2 _25696_ (.A(\count_instr[32] ),
    .B(_19474_),
    .Y(_04105_));
 sky130_fd_sc_hd__o221a_2 _25697_ (.A1(_18606_),
    .A2(_04104_),
    .B1(_04103_),
    .B2(_19012_),
    .C1(_04105_),
    .X(_01715_));
 sky130_fd_sc_hd__buf_1 _25698_ (.A(_18199_),
    .X(_04106_));
 sky130_fd_sc_hd__nand2_2 _25699_ (.A(_19439_),
    .B(\timer[0] ),
    .Y(_04107_));
 sky130_fd_sc_hd__o221a_2 _25700_ (.A1(_18332_),
    .A2(_04106_),
    .B1(_18196_),
    .B2(_18330_),
    .C1(_04107_),
    .X(_01718_));
 sky130_fd_sc_hd__buf_1 _25701_ (.A(_18206_),
    .X(_04108_));
 sky130_fd_sc_hd__nand2_2 _25702_ (.A(_20136_),
    .B(_20135_),
    .Y(_04109_));
 sky130_fd_sc_hd__nand2_2 _25703_ (.A(\decoded_imm[0] ),
    .B(\reg_next_pc[0] ),
    .Y(_04110_));
 sky130_fd_sc_hd__buf_1 _25704_ (.A(_18205_),
    .X(_04111_));
 sky130_fd_sc_hd__buf_1 _25705_ (.A(_04111_),
    .X(_04112_));
 sky130_fd_sc_hd__nor2_2 _25706_ (.A(_01712_),
    .B(_04112_),
    .Y(_04113_));
 sky130_fd_sc_hd__buf_1 _25707_ (.A(_18257_),
    .X(_04114_));
 sky130_fd_sc_hd__a2bb2o_2 _25708_ (.A1_N(_01719_),
    .A2_N(_18851_),
    .B1(_04114_),
    .B2(_01713_),
    .X(_04115_));
 sky130_fd_sc_hd__a311o_2 _25709_ (.A1(_04108_),
    .A2(_04109_),
    .A3(_04110_),
    .B1(_04113_),
    .C1(_04115_),
    .X(_01720_));
 sky130_fd_sc_hd__inv_2 _25710_ (.A(mem_rdata[1]),
    .Y(_01721_));
 sky130_fd_sc_hd__a22o_2 _25711_ (.A1(_04094_),
    .A2(mem_rdata[17]),
    .B1(_04095_),
    .B2(mem_rdata[25]),
    .X(_04116_));
 sky130_fd_sc_hd__a21oi_2 _25712_ (.A1(mem_rdata[9]),
    .A2(_04093_),
    .B1(_04116_),
    .Y(_01722_));
 sky130_fd_sc_hd__o2bb2a_2 _25713_ (.A1_N(_04097_),
    .A2_N(_01724_),
    .B1(_01723_),
    .B2(_20015_),
    .X(_01725_));
 sky130_fd_sc_hd__nand2_2 _25714_ (.A(\count_instr[33] ),
    .B(_19474_),
    .Y(_04117_));
 sky130_fd_sc_hd__o221a_2 _25715_ (.A1(_18605_),
    .A2(_04104_),
    .B1(_04103_),
    .B2(_19016_),
    .C1(_04117_),
    .X(_01729_));
 sky130_fd_sc_hd__buf_1 _25716_ (.A(_18197_),
    .X(_04118_));
 sky130_fd_sc_hd__inv_2 _25717_ (.A(\timer[1] ),
    .Y(_04119_));
 sky130_fd_sc_hd__buf_1 _25718_ (.A(_18208_),
    .X(_04120_));
 sky130_fd_sc_hd__buf_1 _25719_ (.A(_04120_),
    .X(_04121_));
 sky130_fd_sc_hd__nand2_2 _25720_ (.A(\cpuregs_rs1[1] ),
    .B(_04121_),
    .Y(_04122_));
 sky130_fd_sc_hd__o221a_2 _25721_ (.A1(_18327_),
    .A2(_04106_),
    .B1(_04118_),
    .B2(_04119_),
    .C1(_04122_),
    .X(_01731_));
 sky130_fd_sc_hd__nor2_2 _25722_ (.A(\reg_pc[1] ),
    .B(\decoded_imm[1] ),
    .Y(_04123_));
 sky130_fd_sc_hd__nand2_2 _25723_ (.A(\reg_pc[1] ),
    .B(\decoded_imm[1] ),
    .Y(_04124_));
 sky130_fd_sc_hd__or2b_2 _25724_ (.A(_04123_),
    .B_N(_04124_),
    .X(_04125_));
 sky130_fd_sc_hd__or2_2 _25725_ (.A(_04110_),
    .B(_04125_),
    .X(_04126_));
 sky130_fd_sc_hd__buf_1 _25726_ (.A(_18206_),
    .X(_04127_));
 sky130_fd_sc_hd__nand2_2 _25727_ (.A(_04125_),
    .B(_04110_),
    .Y(_04128_));
 sky130_fd_sc_hd__buf_1 _25728_ (.A(_18257_),
    .X(_04129_));
 sky130_fd_sc_hd__o22a_2 _25729_ (.A1(_01726_),
    .A2(_04111_),
    .B1(_19771_),
    .B2(_01732_),
    .X(_04130_));
 sky130_fd_sc_hd__a21bo_2 _25730_ (.A1(_04129_),
    .A2(_01727_),
    .B1_N(_04130_),
    .X(_04131_));
 sky130_fd_sc_hd__a31o_2 _25731_ (.A1(_04126_),
    .A2(_04127_),
    .A3(_04128_),
    .B1(_04131_),
    .X(_01733_));
 sky130_fd_sc_hd__inv_2 _25732_ (.A(mem_rdata[2]),
    .Y(_01734_));
 sky130_fd_sc_hd__a22o_2 _25733_ (.A1(_04094_),
    .A2(mem_rdata[18]),
    .B1(_04095_),
    .B2(mem_rdata[26]),
    .X(_04132_));
 sky130_fd_sc_hd__a21oi_2 _25734_ (.A1(mem_rdata[10]),
    .A2(_04093_),
    .B1(_04132_),
    .Y(_01735_));
 sky130_fd_sc_hd__o2bb2a_2 _25735_ (.A1_N(_04097_),
    .A2_N(_01737_),
    .B1(_01736_),
    .B2(_20015_),
    .X(_01738_));
 sky130_fd_sc_hd__nand2_2 _25736_ (.A(_19482_),
    .B(\count_cycle[34] ),
    .Y(_04133_));
 sky130_fd_sc_hd__o221a_2 _25737_ (.A1(_18715_),
    .A2(_04099_),
    .B1(_18604_),
    .B2(_04101_),
    .C1(_04133_),
    .X(_01742_));
 sky130_fd_sc_hd__buf_1 _25738_ (.A(_04120_),
    .X(_04134_));
 sky130_fd_sc_hd__a22o_2 _25739_ (.A1(\irq_mask[2] ),
    .A2(_19454_),
    .B1(_19439_),
    .B2(\timer[2] ),
    .X(_04135_));
 sky130_fd_sc_hd__a21oi_2 _25740_ (.A1(\cpuregs_rs1[2] ),
    .A2(_04134_),
    .B1(_04135_),
    .Y(_01744_));
 sky130_fd_sc_hd__o21ai_2 _25741_ (.A1(_04110_),
    .A2(_04123_),
    .B1(_04124_),
    .Y(_04136_));
 sky130_fd_sc_hd__xor2_2 _25742_ (.A(\reg_pc[2] ),
    .B(\decoded_imm[2] ),
    .X(_04137_));
 sky130_fd_sc_hd__or2_2 _25743_ (.A(_04136_),
    .B(_04137_),
    .X(_04138_));
 sky130_fd_sc_hd__buf_1 _25744_ (.A(_18206_),
    .X(_04139_));
 sky130_fd_sc_hd__nand2_2 _25745_ (.A(_04137_),
    .B(_04136_),
    .Y(_04140_));
 sky130_fd_sc_hd__a2bb2o_2 _25746_ (.A1_N(_01745_),
    .A2_N(_18851_),
    .B1(_04114_),
    .B2(_01740_),
    .X(_04141_));
 sky130_fd_sc_hd__nor2_2 _25747_ (.A(_01739_),
    .B(_20006_),
    .Y(_04142_));
 sky130_fd_sc_hd__a311o_2 _25748_ (.A1(_04138_),
    .A2(_04139_),
    .A3(_04140_),
    .B1(_04141_),
    .C1(_04142_),
    .X(_01746_));
 sky130_fd_sc_hd__inv_2 _25749_ (.A(mem_rdata[3]),
    .Y(_01747_));
 sky130_fd_sc_hd__a22o_2 _25750_ (.A1(_04094_),
    .A2(mem_rdata[19]),
    .B1(_04095_),
    .B2(mem_rdata[27]),
    .X(_04143_));
 sky130_fd_sc_hd__a21oi_2 _25751_ (.A1(mem_rdata[11]),
    .A2(_04093_),
    .B1(_04143_),
    .Y(_01748_));
 sky130_fd_sc_hd__o2bb2a_2 _25752_ (.A1_N(_04097_),
    .A2_N(_01750_),
    .B1(_01749_),
    .B2(_20015_),
    .X(_01751_));
 sky130_fd_sc_hd__nand2_2 _25753_ (.A(\count_instr[35] ),
    .B(_19474_),
    .Y(_04144_));
 sky130_fd_sc_hd__o221a_2 _25754_ (.A1(_18787_),
    .A2(_04104_),
    .B1(_04103_),
    .B2(_19006_),
    .C1(_04144_),
    .X(_01755_));
 sky130_fd_sc_hd__nand2_2 _25755_ (.A(\cpuregs_rs1[3] ),
    .B(_04121_),
    .Y(_04145_));
 sky130_fd_sc_hd__o221a_2 _25756_ (.A1(_18086_),
    .A2(_04106_),
    .B1(_04118_),
    .B2(_20026_),
    .C1(_04145_),
    .X(_01757_));
 sky130_fd_sc_hd__nor2_2 _25757_ (.A(\reg_pc[3] ),
    .B(\decoded_imm[3] ),
    .Y(_04146_));
 sky130_fd_sc_hd__nand2_2 _25758_ (.A(\reg_pc[3] ),
    .B(\decoded_imm[3] ),
    .Y(_04147_));
 sky130_fd_sc_hd__or2b_2 _25759_ (.A(_04146_),
    .B_N(_04147_),
    .X(_04148_));
 sky130_fd_sc_hd__o21ai_2 _25760_ (.A1(\reg_pc[2] ),
    .A2(\decoded_imm[2] ),
    .B1(_04136_),
    .Y(_04149_));
 sky130_fd_sc_hd__o21a_2 _25761_ (.A1(_02073_),
    .A2(_19702_),
    .B1(_04149_),
    .X(_04150_));
 sky130_fd_sc_hd__or2_2 _25762_ (.A(_04148_),
    .B(_04150_),
    .X(_04151_));
 sky130_fd_sc_hd__nand2_2 _25763_ (.A(_04150_),
    .B(_04148_),
    .Y(_04152_));
 sky130_fd_sc_hd__o22a_2 _25764_ (.A1(_01752_),
    .A2(_04111_),
    .B1(_19771_),
    .B2(_01758_),
    .X(_04153_));
 sky130_fd_sc_hd__a21bo_2 _25765_ (.A1(_04129_),
    .A2(_01753_),
    .B1_N(_04153_),
    .X(_04154_));
 sky130_fd_sc_hd__a31o_2 _25766_ (.A1(_04151_),
    .A2(_04127_),
    .A3(_04152_),
    .B1(_04154_),
    .X(_01759_));
 sky130_fd_sc_hd__inv_2 _25767_ (.A(mem_rdata[4]),
    .Y(_01760_));
 sky130_fd_sc_hd__a22o_2 _25768_ (.A1(_04094_),
    .A2(mem_rdata[20]),
    .B1(_04095_),
    .B2(mem_rdata[28]),
    .X(_04155_));
 sky130_fd_sc_hd__a21oi_2 _25769_ (.A1(mem_rdata[12]),
    .A2(_04093_),
    .B1(_04155_),
    .Y(_01761_));
 sky130_fd_sc_hd__buf_1 _25770_ (.A(_04086_),
    .X(_04156_));
 sky130_fd_sc_hd__o2bb2a_2 _25771_ (.A1_N(_04156_),
    .A2_N(_01763_),
    .B1(_01762_),
    .B2(_20015_),
    .X(_01764_));
 sky130_fd_sc_hd__buf_1 _25772_ (.A(instr_rdinstrh),
    .X(_04157_));
 sky130_fd_sc_hd__nand2_2 _25773_ (.A(\count_instr[36] ),
    .B(_04157_),
    .Y(_04158_));
 sky130_fd_sc_hd__o221a_2 _25774_ (.A1(_18789_),
    .A2(_04104_),
    .B1(_04103_),
    .B2(_19005_),
    .C1(_04158_),
    .X(_01768_));
 sky130_fd_sc_hd__a22o_2 _25775_ (.A1(\irq_mask[4] ),
    .A2(_19454_),
    .B1(_19439_),
    .B2(\timer[4] ),
    .X(_04159_));
 sky130_fd_sc_hd__a21oi_2 _25776_ (.A1(\cpuregs_rs1[4] ),
    .A2(_04134_),
    .B1(_04159_),
    .Y(_01770_));
 sky130_fd_sc_hd__nand2_2 _25777_ (.A(_20153_),
    .B(_19713_),
    .Y(_04160_));
 sky130_fd_sc_hd__nand2_2 _25778_ (.A(\reg_pc[4] ),
    .B(\decoded_imm[4] ),
    .Y(_04161_));
 sky130_fd_sc_hd__and2_2 _25779_ (.A(_04160_),
    .B(_04161_),
    .X(_04162_));
 sky130_fd_sc_hd__o21ai_2 _25780_ (.A1(_04146_),
    .A2(_04150_),
    .B1(_04147_),
    .Y(_04163_));
 sky130_fd_sc_hd__or2_2 _25781_ (.A(_04162_),
    .B(_04163_),
    .X(_04164_));
 sky130_fd_sc_hd__nand2_2 _25782_ (.A(_04163_),
    .B(_04162_),
    .Y(_04165_));
 sky130_fd_sc_hd__o22a_2 _25783_ (.A1(_01765_),
    .A2(_04111_),
    .B1(_19771_),
    .B2(_01771_),
    .X(_04166_));
 sky130_fd_sc_hd__a21bo_2 _25784_ (.A1(_04129_),
    .A2(_01766_),
    .B1_N(_04166_),
    .X(_04167_));
 sky130_fd_sc_hd__a31o_2 _25785_ (.A1(_04164_),
    .A2(_04127_),
    .A3(_04165_),
    .B1(_04167_),
    .X(_01772_));
 sky130_fd_sc_hd__inv_2 _25786_ (.A(mem_rdata[5]),
    .Y(_01773_));
 sky130_fd_sc_hd__a22o_2 _25787_ (.A1(_04094_),
    .A2(mem_rdata[21]),
    .B1(_04095_),
    .B2(mem_rdata[29]),
    .X(_04168_));
 sky130_fd_sc_hd__a21oi_2 _25788_ (.A1(mem_rdata[13]),
    .A2(_04093_),
    .B1(_04168_),
    .Y(_01774_));
 sky130_fd_sc_hd__o2bb2a_2 _25789_ (.A1_N(_04156_),
    .A2_N(_01776_),
    .B1(_01775_),
    .B2(_20014_),
    .X(_01777_));
 sky130_fd_sc_hd__buf_1 _25790_ (.A(instr_rdinstrh),
    .X(_04169_));
 sky130_fd_sc_hd__a22o_2 _25791_ (.A1(_18692_),
    .A2(_04169_),
    .B1(\count_instr[5] ),
    .B2(instr_rdinstr),
    .X(_04170_));
 sky130_fd_sc_hd__a21oi_2 _25792_ (.A1(_19482_),
    .A2(\count_cycle[37] ),
    .B1(_04170_),
    .Y(_01781_));
 sky130_fd_sc_hd__a22o_2 _25793_ (.A1(\irq_mask[5] ),
    .A2(_19454_),
    .B1(_19439_),
    .B2(\timer[5] ),
    .X(_04171_));
 sky130_fd_sc_hd__a21oi_2 _25794_ (.A1(\cpuregs_rs1[5] ),
    .A2(_04134_),
    .B1(_04171_),
    .Y(_01783_));
 sky130_fd_sc_hd__nor2_2 _25795_ (.A(\reg_pc[5] ),
    .B(\decoded_imm[5] ),
    .Y(_04172_));
 sky130_fd_sc_hd__nand2_2 _25796_ (.A(\reg_pc[5] ),
    .B(\decoded_imm[5] ),
    .Y(_04173_));
 sky130_fd_sc_hd__and2b_2 _25797_ (.A_N(_04172_),
    .B(_04173_),
    .X(_04174_));
 sky130_fd_sc_hd__nand2_2 _25798_ (.A(_04165_),
    .B(_04161_),
    .Y(_04175_));
 sky130_fd_sc_hd__or2_2 _25799_ (.A(_04174_),
    .B(_04175_),
    .X(_04176_));
 sky130_fd_sc_hd__nand2_2 _25800_ (.A(_04175_),
    .B(_04174_),
    .Y(_04177_));
 sky130_fd_sc_hd__a2bb2o_2 _25801_ (.A1_N(_01784_),
    .A2_N(_18851_),
    .B1(_04114_),
    .B2(_01779_),
    .X(_04178_));
 sky130_fd_sc_hd__buf_1 _25802_ (.A(_18444_),
    .X(_04179_));
 sky130_fd_sc_hd__nor2_2 _25803_ (.A(_01778_),
    .B(_04179_),
    .Y(_04180_));
 sky130_fd_sc_hd__a311o_2 _25804_ (.A1(_04176_),
    .A2(_04139_),
    .A3(_04177_),
    .B1(_04178_),
    .C1(_04180_),
    .X(_01785_));
 sky130_fd_sc_hd__inv_2 _25805_ (.A(mem_rdata[6]),
    .Y(_01786_));
 sky130_fd_sc_hd__a22o_2 _25806_ (.A1(_04088_),
    .A2(mem_rdata[22]),
    .B1(_04090_),
    .B2(mem_rdata[30]),
    .X(_04181_));
 sky130_fd_sc_hd__a21oi_2 _25807_ (.A1(mem_rdata[14]),
    .A2(_04092_),
    .B1(_04181_),
    .Y(_01787_));
 sky130_fd_sc_hd__o2bb2a_2 _25808_ (.A1_N(_04156_),
    .A2_N(_01789_),
    .B1(_01788_),
    .B2(_20014_),
    .X(_01790_));
 sky130_fd_sc_hd__nand2_2 _25809_ (.A(\count_instr[38] ),
    .B(_04157_),
    .Y(_04182_));
 sky130_fd_sc_hd__o221a_2 _25810_ (.A1(_18598_),
    .A2(_04104_),
    .B1(_04103_),
    .B2(_18991_),
    .C1(_04182_),
    .X(_01794_));
 sky130_fd_sc_hd__a22o_2 _25811_ (.A1(\irq_mask[6] ),
    .A2(_19454_),
    .B1(_19439_),
    .B2(\timer[6] ),
    .X(_04183_));
 sky130_fd_sc_hd__a21oi_2 _25812_ (.A1(\cpuregs_rs1[6] ),
    .A2(_04134_),
    .B1(_04183_),
    .Y(_01796_));
 sky130_fd_sc_hd__nand3_2 _25813_ (.A(_04163_),
    .B(_04162_),
    .C(_04174_),
    .Y(_04184_));
 sky130_fd_sc_hd__o21a_2 _25814_ (.A1(_04161_),
    .A2(_04172_),
    .B1(_04173_),
    .X(_04185_));
 sky130_fd_sc_hd__nand2_2 _25815_ (.A(_18564_),
    .B(_20105_),
    .Y(_04186_));
 sky130_fd_sc_hd__nand2_2 _25816_ (.A(\reg_pc[6] ),
    .B(\decoded_imm[6] ),
    .Y(_04187_));
 sky130_fd_sc_hd__nand2_2 _25817_ (.A(_04186_),
    .B(_04187_),
    .Y(_04188_));
 sky130_fd_sc_hd__a31o_2 _25818_ (.A1(_04184_),
    .A2(_04185_),
    .A3(_04188_),
    .B1(_18186_),
    .X(_04189_));
 sky130_fd_sc_hd__nand2_2 _25819_ (.A(_04184_),
    .B(_04185_),
    .Y(_04190_));
 sky130_fd_sc_hd__inv_2 _25820_ (.A(_04190_),
    .Y(_04191_));
 sky130_fd_sc_hd__nor2_2 _25821_ (.A(_04188_),
    .B(_04191_),
    .Y(_04192_));
 sky130_fd_sc_hd__buf_1 _25822_ (.A(_18257_),
    .X(_04193_));
 sky130_fd_sc_hd__buf_1 _25823_ (.A(_18194_),
    .X(_04194_));
 sky130_fd_sc_hd__o2bb2a_2 _25824_ (.A1_N(_04193_),
    .A2_N(_01792_),
    .B1(_01797_),
    .B2(_04194_),
    .X(_04195_));
 sky130_fd_sc_hd__o221ai_2 _25825_ (.A1(_20006_),
    .A2(_01791_),
    .B1(_04189_),
    .B2(_04192_),
    .C1(_04195_),
    .Y(_01798_));
 sky130_fd_sc_hd__inv_2 _25826_ (.A(mem_rdata[7]),
    .Y(_01799_));
 sky130_fd_sc_hd__a22o_2 _25827_ (.A1(_04088_),
    .A2(mem_rdata[23]),
    .B1(_04090_),
    .B2(mem_rdata[31]),
    .X(_04196_));
 sky130_fd_sc_hd__a21oi_2 _25828_ (.A1(mem_rdata[15]),
    .A2(_04092_),
    .B1(_04196_),
    .Y(_01800_));
 sky130_fd_sc_hd__o2bb2a_2 _25829_ (.A1_N(_04156_),
    .A2_N(_01802_),
    .B1(_01801_),
    .B2(_20014_),
    .X(_01803_));
 sky130_fd_sc_hd__buf_1 _25830_ (.A(_04102_),
    .X(_04197_));
 sky130_fd_sc_hd__buf_1 _25831_ (.A(_04197_),
    .X(_04198_));
 sky130_fd_sc_hd__nand2_2 _25832_ (.A(\count_instr[39] ),
    .B(_04157_),
    .Y(_04199_));
 sky130_fd_sc_hd__o221a_2 _25833_ (.A1(_18597_),
    .A2(_04104_),
    .B1(_04198_),
    .B2(_18992_),
    .C1(_04199_),
    .X(_01807_));
 sky130_fd_sc_hd__nand2_2 _25834_ (.A(\cpuregs_rs1[7] ),
    .B(_04121_),
    .Y(_04200_));
 sky130_fd_sc_hd__o221a_2 _25835_ (.A1(_18118_),
    .A2(_04106_),
    .B1(_04118_),
    .B2(_20061_),
    .C1(_04200_),
    .X(_01809_));
 sky130_fd_sc_hd__inv_2 _25836_ (.A(_01804_),
    .Y(_04201_));
 sky130_fd_sc_hd__buf_1 _25837_ (.A(_04193_),
    .X(_04202_));
 sky130_fd_sc_hd__nor2_2 _25838_ (.A(_20172_),
    .B(_20106_),
    .Y(_04203_));
 sky130_fd_sc_hd__inv_2 _25839_ (.A(_04203_),
    .Y(_04204_));
 sky130_fd_sc_hd__nor2_2 _25840_ (.A(\reg_pc[7] ),
    .B(\decoded_imm[7] ),
    .Y(_04205_));
 sky130_fd_sc_hd__inv_2 _25841_ (.A(_04205_),
    .Y(_04206_));
 sky130_fd_sc_hd__nand2_2 _25842_ (.A(_04204_),
    .B(_04206_),
    .Y(_04207_));
 sky130_fd_sc_hd__inv_2 _25843_ (.A(_04207_),
    .Y(_04208_));
 sky130_fd_sc_hd__inv_2 _25844_ (.A(_04187_),
    .Y(_04209_));
 sky130_fd_sc_hd__or2_2 _25845_ (.A(_04209_),
    .B(_04192_),
    .X(_04210_));
 sky130_fd_sc_hd__or2_2 _25846_ (.A(_04208_),
    .B(_04210_),
    .X(_04211_));
 sky130_fd_sc_hd__nand2_2 _25847_ (.A(_04210_),
    .B(_04208_),
    .Y(_04212_));
 sky130_fd_sc_hd__nor2_2 _25848_ (.A(_01810_),
    .B(_19188_),
    .Y(_04213_));
 sky130_fd_sc_hd__a31o_2 _25849_ (.A1(_04211_),
    .A2(_18206_),
    .A3(_04212_),
    .B1(_04213_),
    .X(_04214_));
 sky130_fd_sc_hd__a221o_2 _25850_ (.A1(_18029_),
    .A2(_04201_),
    .B1(_04202_),
    .B2(_01805_),
    .C1(_04214_),
    .X(_01811_));
 sky130_fd_sc_hd__inv_2 _25851_ (.A(mem_rdata[8]),
    .Y(_01812_));
 sky130_fd_sc_hd__buf_1 _25852_ (.A(_04086_),
    .X(_04215_));
 sky130_fd_sc_hd__nand2_2 _25853_ (.A(_04215_),
    .B(_01813_),
    .Y(_01814_));
 sky130_fd_sc_hd__nor2_2 _25854_ (.A(latched_is_lb),
    .B(latched_is_lh),
    .Y(_01816_));
 sky130_fd_sc_hd__inv_2 _25855_ (.A(latched_is_lh),
    .Y(_04216_));
 sky130_fd_sc_hd__buf_1 _25856_ (.A(_04216_),
    .X(_04217_));
 sky130_fd_sc_hd__nand2_2 _25857_ (.A(_04201_),
    .B(latched_is_lb),
    .Y(_04218_));
 sky130_fd_sc_hd__buf_1 _25858_ (.A(_04218_),
    .X(_04219_));
 sky130_fd_sc_hd__o21a_2 _25859_ (.A1(_04217_),
    .A2(_01815_),
    .B1(_04219_),
    .X(_01817_));
 sky130_fd_sc_hd__nand2_2 _25860_ (.A(\count_instr[8] ),
    .B(_19478_),
    .Y(_04220_));
 sky130_fd_sc_hd__o221a_2 _25861_ (.A1(_18697_),
    .A2(_04099_),
    .B1(_04198_),
    .B2(_18998_),
    .C1(_04220_),
    .X(_01821_));
 sky130_fd_sc_hd__nand2_2 _25862_ (.A(\cpuregs_rs1[8] ),
    .B(_04121_),
    .Y(_04221_));
 sky130_fd_sc_hd__o221a_2 _25863_ (.A1(_18115_),
    .A2(_04106_),
    .B1(_04118_),
    .B2(_20063_),
    .C1(_04221_),
    .X(_01823_));
 sky130_fd_sc_hd__nand2_2 _25864_ (.A(_20177_),
    .B(_20107_),
    .Y(_04222_));
 sky130_fd_sc_hd__nand2_2 _25865_ (.A(\reg_pc[8] ),
    .B(\decoded_imm[8] ),
    .Y(_04223_));
 sky130_fd_sc_hd__nand2_2 _25866_ (.A(_04222_),
    .B(_04223_),
    .Y(_04224_));
 sky130_fd_sc_hd__a21oi_2 _25867_ (.A1(_04206_),
    .A2(_04209_),
    .B1(_04203_),
    .Y(_04225_));
 sky130_fd_sc_hd__inv_2 _25868_ (.A(_04225_),
    .Y(_04226_));
 sky130_fd_sc_hd__or2_2 _25869_ (.A(_04188_),
    .B(_04207_),
    .X(_04227_));
 sky130_fd_sc_hd__a21oi_2 _25870_ (.A1(_04184_),
    .A2(_04185_),
    .B1(_04227_),
    .Y(_04228_));
 sky130_fd_sc_hd__nor2_2 _25871_ (.A(_04226_),
    .B(_04228_),
    .Y(_04229_));
 sky130_fd_sc_hd__or2_2 _25872_ (.A(_04224_),
    .B(_04229_),
    .X(_04230_));
 sky130_fd_sc_hd__a21oi_2 _25873_ (.A1(_04229_),
    .A2(_04224_),
    .B1(_18187_),
    .Y(_04231_));
 sky130_fd_sc_hd__buf_1 _25874_ (.A(_18799_),
    .X(_04232_));
 sky130_fd_sc_hd__o22ai_2 _25875_ (.A1(_01818_),
    .A2(_04112_),
    .B1(_04232_),
    .B2(_01824_),
    .Y(_04233_));
 sky130_fd_sc_hd__a221o_2 _25876_ (.A1(_04202_),
    .A2(_01819_),
    .B1(_04230_),
    .B2(_04231_),
    .C1(_04233_),
    .X(_01825_));
 sky130_fd_sc_hd__inv_2 _25877_ (.A(mem_rdata[9]),
    .Y(_01826_));
 sky130_fd_sc_hd__nand2_2 _25878_ (.A(_04215_),
    .B(_01827_),
    .Y(_01828_));
 sky130_fd_sc_hd__o21a_2 _25879_ (.A1(_04217_),
    .A2(_01829_),
    .B1(_04219_),
    .X(_01830_));
 sky130_fd_sc_hd__nand2_2 _25880_ (.A(_19482_),
    .B(_18986_),
    .Y(_04234_));
 sky130_fd_sc_hd__o221a_2 _25881_ (.A1(_18696_),
    .A2(_04099_),
    .B1(_18601_),
    .B2(_04101_),
    .C1(_04234_),
    .X(_01834_));
 sky130_fd_sc_hd__buf_1 _25882_ (.A(_19438_),
    .X(_04235_));
 sky130_fd_sc_hd__a22o_2 _25883_ (.A1(\irq_mask[9] ),
    .A2(_19454_),
    .B1(_04235_),
    .B2(\timer[9] ),
    .X(_04236_));
 sky130_fd_sc_hd__a21oi_2 _25884_ (.A1(\cpuregs_rs1[9] ),
    .A2(_04134_),
    .B1(_04236_),
    .Y(_01836_));
 sky130_fd_sc_hd__nor2_2 _25885_ (.A(\reg_pc[9] ),
    .B(\decoded_imm[9] ),
    .Y(_04237_));
 sky130_fd_sc_hd__nor2_2 _25886_ (.A(_20185_),
    .B(_20108_),
    .Y(_04238_));
 sky130_fd_sc_hd__or2_2 _25887_ (.A(_04237_),
    .B(_04238_),
    .X(_04239_));
 sky130_fd_sc_hd__inv_2 _25888_ (.A(_04239_),
    .Y(_04240_));
 sky130_fd_sc_hd__nand2_2 _25889_ (.A(_04230_),
    .B(_04223_),
    .Y(_04241_));
 sky130_fd_sc_hd__or2_2 _25890_ (.A(_04240_),
    .B(_04241_),
    .X(_04242_));
 sky130_fd_sc_hd__nand2_2 _25891_ (.A(_04241_),
    .B(_04240_),
    .Y(_04243_));
 sky130_fd_sc_hd__a2bb2o_2 _25892_ (.A1_N(_01837_),
    .A2_N(_04194_),
    .B1(_04114_),
    .B2(_01832_),
    .X(_04244_));
 sky130_fd_sc_hd__nor2_2 _25893_ (.A(_01831_),
    .B(_04179_),
    .Y(_04245_));
 sky130_fd_sc_hd__a311o_2 _25894_ (.A1(_04242_),
    .A2(_04139_),
    .A3(_04243_),
    .B1(_04244_),
    .C1(_04245_),
    .X(_01838_));
 sky130_fd_sc_hd__inv_2 _25895_ (.A(mem_rdata[10]),
    .Y(_01839_));
 sky130_fd_sc_hd__nand2_2 _25896_ (.A(_04215_),
    .B(_01840_),
    .Y(_01841_));
 sky130_fd_sc_hd__o21a_2 _25897_ (.A1(_04217_),
    .A2(_01842_),
    .B1(_04219_),
    .X(_01843_));
 sky130_fd_sc_hd__buf_1 _25898_ (.A(instr_rdcycleh),
    .X(_04246_));
 sky130_fd_sc_hd__a22o_2 _25899_ (.A1(\count_instr[10] ),
    .A2(instr_rdinstr),
    .B1(_04246_),
    .B2(\count_cycle[42] ),
    .X(_04247_));
 sky130_fd_sc_hd__a21oi_2 _25900_ (.A1(\count_instr[42] ),
    .A2(_19474_),
    .B1(_04247_),
    .Y(_01847_));
 sky130_fd_sc_hd__buf_1 _25901_ (.A(_18198_),
    .X(_04248_));
 sky130_fd_sc_hd__a22o_2 _25902_ (.A1(\irq_mask[10] ),
    .A2(_04248_),
    .B1(_04235_),
    .B2(\timer[10] ),
    .X(_04249_));
 sky130_fd_sc_hd__a21oi_2 _25903_ (.A1(\cpuregs_rs1[10] ),
    .A2(_04134_),
    .B1(_04249_),
    .Y(_01849_));
 sky130_fd_sc_hd__o22ai_2 _25904_ (.A1(_01844_),
    .A2(_04112_),
    .B1(_04232_),
    .B2(_01850_),
    .Y(_04250_));
 sky130_fd_sc_hd__or2_2 _25905_ (.A(_04224_),
    .B(_04239_),
    .X(_04251_));
 sky130_fd_sc_hd__o21bai_2 _25906_ (.A1(_04226_),
    .A2(_04228_),
    .B1_N(_04251_),
    .Y(_04252_));
 sky130_fd_sc_hd__o21ba_2 _25907_ (.A1(_04223_),
    .A2(_04237_),
    .B1_N(_04238_),
    .X(_04253_));
 sky130_fd_sc_hd__and2_2 _25908_ (.A(_04252_),
    .B(_04253_),
    .X(_04254_));
 sky130_fd_sc_hd__nor2_2 _25909_ (.A(_20191_),
    .B(_20109_),
    .Y(_04255_));
 sky130_fd_sc_hd__nor2_2 _25910_ (.A(\reg_pc[10] ),
    .B(\decoded_imm[10] ),
    .Y(_04256_));
 sky130_fd_sc_hd__or2_2 _25911_ (.A(_04256_),
    .B(_04255_),
    .X(_04257_));
 sky130_fd_sc_hd__a21oi_2 _25912_ (.A1(_04254_),
    .A2(_04257_),
    .B1(_18186_),
    .Y(_04258_));
 sky130_fd_sc_hd__o31a_2 _25913_ (.A1(_04254_),
    .A2(_04255_),
    .A3(_04256_),
    .B1(_04258_),
    .X(_04259_));
 sky130_fd_sc_hd__a211o_2 _25914_ (.A1(_04202_),
    .A2(_01845_),
    .B1(_04250_),
    .C1(_04259_),
    .X(_01851_));
 sky130_fd_sc_hd__inv_2 _25915_ (.A(mem_rdata[11]),
    .Y(_01852_));
 sky130_fd_sc_hd__nand2_2 _25916_ (.A(_04215_),
    .B(_01853_),
    .Y(_01854_));
 sky130_fd_sc_hd__o21a_2 _25917_ (.A1(_04217_),
    .A2(_01855_),
    .B1(_04219_),
    .X(_01856_));
 sky130_fd_sc_hd__nand2_2 _25918_ (.A(_19482_),
    .B(\count_cycle[43] ),
    .Y(_04260_));
 sky130_fd_sc_hd__o221a_2 _25919_ (.A1(_18584_),
    .A2(_04099_),
    .B1(_18596_),
    .B2(_04101_),
    .C1(_04260_),
    .X(_01860_));
 sky130_fd_sc_hd__buf_1 _25920_ (.A(_04120_),
    .X(_04261_));
 sky130_fd_sc_hd__a22o_2 _25921_ (.A1(\irq_mask[11] ),
    .A2(_04248_),
    .B1(_04235_),
    .B2(\timer[11] ),
    .X(_04262_));
 sky130_fd_sc_hd__a21oi_2 _25922_ (.A1(\cpuregs_rs1[11] ),
    .A2(_04261_),
    .B1(_04262_),
    .Y(_01862_));
 sky130_fd_sc_hd__nand2_2 _25923_ (.A(_18552_),
    .B(_20111_),
    .Y(_04263_));
 sky130_fd_sc_hd__nand2_2 _25924_ (.A(\reg_pc[11] ),
    .B(\decoded_imm[11] ),
    .Y(_04264_));
 sky130_fd_sc_hd__nand2_2 _25925_ (.A(_04263_),
    .B(_04264_),
    .Y(_04265_));
 sky130_fd_sc_hd__a21oi_2 _25926_ (.A1(_04252_),
    .A2(_04253_),
    .B1(_04256_),
    .Y(_04266_));
 sky130_fd_sc_hd__nor2_2 _25927_ (.A(_04255_),
    .B(_04266_),
    .Y(_04267_));
 sky130_fd_sc_hd__or2_2 _25928_ (.A(_04265_),
    .B(_04267_),
    .X(_04268_));
 sky130_fd_sc_hd__nand2_2 _25929_ (.A(_04267_),
    .B(_04265_),
    .Y(_04269_));
 sky130_fd_sc_hd__a2bb2o_2 _25930_ (.A1_N(_01863_),
    .A2_N(_04194_),
    .B1(_19851_),
    .B2(_01858_),
    .X(_04270_));
 sky130_fd_sc_hd__nor2_2 _25931_ (.A(_01857_),
    .B(_04179_),
    .Y(_04271_));
 sky130_fd_sc_hd__a311o_2 _25932_ (.A1(_04268_),
    .A2(_04139_),
    .A3(_04269_),
    .B1(_04270_),
    .C1(_04271_),
    .X(_01864_));
 sky130_fd_sc_hd__inv_2 _25933_ (.A(mem_rdata[12]),
    .Y(_01865_));
 sky130_fd_sc_hd__nand2_2 _25934_ (.A(_04215_),
    .B(_01866_),
    .Y(_01867_));
 sky130_fd_sc_hd__o21a_2 _25935_ (.A1(_04217_),
    .A2(_01868_),
    .B1(_04219_),
    .X(_01869_));
 sky130_fd_sc_hd__nand2_2 _25936_ (.A(_19482_),
    .B(\count_cycle[44] ),
    .Y(_04272_));
 sky130_fd_sc_hd__o221a_2 _25937_ (.A1(_18689_),
    .A2(_04099_),
    .B1(_18595_),
    .B2(_04101_),
    .C1(_04272_),
    .X(_01873_));
 sky130_fd_sc_hd__a22o_2 _25938_ (.A1(\irq_mask[12] ),
    .A2(_04248_),
    .B1(_04235_),
    .B2(\timer[12] ),
    .X(_04273_));
 sky130_fd_sc_hd__a21oi_2 _25939_ (.A1(\cpuregs_rs1[12] ),
    .A2(_04261_),
    .B1(_04273_),
    .Y(_01875_));
 sky130_fd_sc_hd__nor2_2 _25940_ (.A(\reg_pc[12] ),
    .B(\decoded_imm[12] ),
    .Y(_04274_));
 sky130_fd_sc_hd__nor2_2 _25941_ (.A(_20208_),
    .B(_20112_),
    .Y(_04275_));
 sky130_fd_sc_hd__nor2_2 _25942_ (.A(_04274_),
    .B(_04275_),
    .Y(_04276_));
 sky130_fd_sc_hd__o21ai_2 _25943_ (.A1(_04255_),
    .A2(_04266_),
    .B1(_04263_),
    .Y(_04277_));
 sky130_fd_sc_hd__nand2_2 _25944_ (.A(_04277_),
    .B(_04264_),
    .Y(_04278_));
 sky130_fd_sc_hd__or2_2 _25945_ (.A(_04276_),
    .B(_04278_),
    .X(_04279_));
 sky130_fd_sc_hd__nand2_2 _25946_ (.A(_04278_),
    .B(_04276_),
    .Y(_04280_));
 sky130_fd_sc_hd__nand2_2 _25947_ (.A(_04193_),
    .B(_01871_),
    .Y(_04281_));
 sky130_fd_sc_hd__o221ai_2 _25948_ (.A1(_01870_),
    .A2(_04112_),
    .B1(_01876_),
    .B2(_04232_),
    .C1(_04281_),
    .Y(_04282_));
 sky130_fd_sc_hd__a31o_2 _25949_ (.A1(_04279_),
    .A2(_04127_),
    .A3(_04280_),
    .B1(_04282_),
    .X(_01877_));
 sky130_fd_sc_hd__inv_2 _25950_ (.A(mem_rdata[13]),
    .Y(_01878_));
 sky130_fd_sc_hd__nand2_2 _25951_ (.A(_04215_),
    .B(_01879_),
    .Y(_01880_));
 sky130_fd_sc_hd__o21a_2 _25952_ (.A1(_04217_),
    .A2(_01881_),
    .B1(_04219_),
    .X(_01882_));
 sky130_fd_sc_hd__buf_1 _25953_ (.A(_04098_),
    .X(_04283_));
 sky130_fd_sc_hd__nand2_2 _25954_ (.A(\count_instr[13] ),
    .B(_19478_),
    .Y(_04284_));
 sky130_fd_sc_hd__o221a_2 _25955_ (.A1(_18681_),
    .A2(_04283_),
    .B1(_04198_),
    .B2(_18978_),
    .C1(_04284_),
    .X(_01886_));
 sky130_fd_sc_hd__a22o_2 _25956_ (.A1(\irq_mask[13] ),
    .A2(_04248_),
    .B1(_04235_),
    .B2(\timer[13] ),
    .X(_04285_));
 sky130_fd_sc_hd__a21oi_2 _25957_ (.A1(\cpuregs_rs1[13] ),
    .A2(_04261_),
    .B1(_04285_),
    .Y(_01888_));
 sky130_fd_sc_hd__nor2_2 _25958_ (.A(_20215_),
    .B(_20113_),
    .Y(_04286_));
 sky130_fd_sc_hd__inv_2 _25959_ (.A(_04286_),
    .Y(_04287_));
 sky130_fd_sc_hd__nor2_2 _25960_ (.A(\reg_pc[13] ),
    .B(\decoded_imm[13] ),
    .Y(_04288_));
 sky130_fd_sc_hd__inv_2 _25961_ (.A(_04288_),
    .Y(_04289_));
 sky130_fd_sc_hd__nand2_2 _25962_ (.A(_04287_),
    .B(_04289_),
    .Y(_04290_));
 sky130_fd_sc_hd__a21oi_2 _25963_ (.A1(_04277_),
    .A2(_04264_),
    .B1(_04274_),
    .Y(_04291_));
 sky130_fd_sc_hd__nor2_2 _25964_ (.A(_04275_),
    .B(_04291_),
    .Y(_04292_));
 sky130_fd_sc_hd__or2_2 _25965_ (.A(_04290_),
    .B(_04292_),
    .X(_04293_));
 sky130_fd_sc_hd__buf_1 _25966_ (.A(_18206_),
    .X(_04294_));
 sky130_fd_sc_hd__nand2_2 _25967_ (.A(_04292_),
    .B(_04290_),
    .Y(_04295_));
 sky130_fd_sc_hd__a2bb2o_2 _25968_ (.A1_N(_01889_),
    .A2_N(_04194_),
    .B1(_19851_),
    .B2(_01884_),
    .X(_04296_));
 sky130_fd_sc_hd__nor2_2 _25969_ (.A(_01883_),
    .B(_04179_),
    .Y(_04297_));
 sky130_fd_sc_hd__a311o_2 _25970_ (.A1(_04293_),
    .A2(_04294_),
    .A3(_04295_),
    .B1(_04296_),
    .C1(_04297_),
    .X(_01890_));
 sky130_fd_sc_hd__inv_2 _25971_ (.A(mem_rdata[14]),
    .Y(_01891_));
 sky130_fd_sc_hd__nand2_2 _25972_ (.A(_04097_),
    .B(_01892_),
    .Y(_01893_));
 sky130_fd_sc_hd__o21a_2 _25973_ (.A1(_04216_),
    .A2(_01894_),
    .B1(_04218_),
    .X(_01895_));
 sky130_fd_sc_hd__inv_2 _25974_ (.A(\count_cycle[14] ),
    .Y(_01898_));
 sky130_fd_sc_hd__buf_1 _25975_ (.A(_04100_),
    .X(_04298_));
 sky130_fd_sc_hd__nand2_2 _25976_ (.A(\count_instr[46] ),
    .B(_04157_),
    .Y(_04299_));
 sky130_fd_sc_hd__o221a_2 _25977_ (.A1(_18759_),
    .A2(_04298_),
    .B1(_04198_),
    .B2(_18981_),
    .C1(_04299_),
    .X(_01899_));
 sky130_fd_sc_hd__nand2_2 _25978_ (.A(\cpuregs_rs1[14] ),
    .B(_04121_),
    .Y(_04300_));
 sky130_fd_sc_hd__o221a_2 _25979_ (.A1(_18139_),
    .A2(_04106_),
    .B1(_04118_),
    .B2(_20039_),
    .C1(_04300_),
    .X(_01901_));
 sky130_fd_sc_hd__nor2_2 _25980_ (.A(\reg_pc[14] ),
    .B(\decoded_imm[14] ),
    .Y(_04301_));
 sky130_fd_sc_hd__nor2_2 _25981_ (.A(_20222_),
    .B(_20114_),
    .Y(_04302_));
 sky130_fd_sc_hd__or2_2 _25982_ (.A(_04301_),
    .B(_04302_),
    .X(_04303_));
 sky130_fd_sc_hd__o21ai_2 _25983_ (.A1(_04275_),
    .A2(_04291_),
    .B1(_04289_),
    .Y(_04304_));
 sky130_fd_sc_hd__and2_2 _25984_ (.A(_04304_),
    .B(_04287_),
    .X(_04305_));
 sky130_fd_sc_hd__or2_2 _25985_ (.A(_04303_),
    .B(_04305_),
    .X(_04306_));
 sky130_fd_sc_hd__nand2_2 _25986_ (.A(_04305_),
    .B(_04303_),
    .Y(_04307_));
 sky130_fd_sc_hd__o22a_2 _25987_ (.A1(_01896_),
    .A2(_04111_),
    .B1(_19771_),
    .B2(_01902_),
    .X(_04308_));
 sky130_fd_sc_hd__a21bo_2 _25988_ (.A1(_04129_),
    .A2(_01897_),
    .B1_N(_04308_),
    .X(_04309_));
 sky130_fd_sc_hd__a31o_2 _25989_ (.A1(_04306_),
    .A2(_04127_),
    .A3(_04307_),
    .B1(_04309_),
    .X(_01903_));
 sky130_fd_sc_hd__inv_2 _25990_ (.A(mem_rdata[15]),
    .Y(_01904_));
 sky130_fd_sc_hd__nand2_2 _25991_ (.A(_04097_),
    .B(_01905_),
    .Y(_01906_));
 sky130_fd_sc_hd__o21a_2 _25992_ (.A1(_04216_),
    .A2(_01907_),
    .B1(_04218_),
    .X(_01908_));
 sky130_fd_sc_hd__a22o_2 _25993_ (.A1(\count_instr[47] ),
    .A2(_04169_),
    .B1(_04246_),
    .B2(\count_cycle[47] ),
    .X(_04310_));
 sky130_fd_sc_hd__a21oi_2 _25994_ (.A1(\count_instr[15] ),
    .A2(_19478_),
    .B1(_04310_),
    .Y(_01912_));
 sky130_fd_sc_hd__a22o_2 _25995_ (.A1(\irq_mask[15] ),
    .A2(_04248_),
    .B1(_04235_),
    .B2(\timer[15] ),
    .X(_04311_));
 sky130_fd_sc_hd__a21oi_2 _25996_ (.A1(\cpuregs_rs1[15] ),
    .A2(_04261_),
    .B1(_04311_),
    .Y(_01914_));
 sky130_fd_sc_hd__nor2_2 _25997_ (.A(\reg_pc[15] ),
    .B(\decoded_imm[15] ),
    .Y(_04312_));
 sky130_fd_sc_hd__nor2_2 _25998_ (.A(_20227_),
    .B(_20115_),
    .Y(_04313_));
 sky130_fd_sc_hd__or2_2 _25999_ (.A(_04312_),
    .B(_04313_),
    .X(_04314_));
 sky130_fd_sc_hd__a21oi_2 _26000_ (.A1(_04304_),
    .A2(_04287_),
    .B1(_04301_),
    .Y(_04315_));
 sky130_fd_sc_hd__nor2_2 _26001_ (.A(_04302_),
    .B(_04315_),
    .Y(_04316_));
 sky130_fd_sc_hd__nor2_2 _26002_ (.A(_04314_),
    .B(_04316_),
    .Y(_04317_));
 sky130_fd_sc_hd__a21o_2 _26003_ (.A1(_04316_),
    .A2(_04314_),
    .B1(_18187_),
    .X(_04318_));
 sky130_fd_sc_hd__o2bb2a_2 _26004_ (.A1_N(_04193_),
    .A2_N(_01910_),
    .B1(_01915_),
    .B2(_19188_),
    .X(_04319_));
 sky130_fd_sc_hd__o221ai_2 _26005_ (.A1(_20006_),
    .A2(_01909_),
    .B1(_04317_),
    .B2(_04318_),
    .C1(_04319_),
    .Y(_01916_));
 sky130_fd_sc_hd__nand2_2 _26006_ (.A(_01683_),
    .B(mem_rdata[16]),
    .Y(_01917_));
 sky130_fd_sc_hd__buf_1 _26007_ (.A(_04246_),
    .X(_04320_));
 sky130_fd_sc_hd__nand2_2 _26008_ (.A(_04320_),
    .B(\count_cycle[48] ),
    .Y(_04321_));
 sky130_fd_sc_hd__o221a_2 _26009_ (.A1(_18586_),
    .A2(_04283_),
    .B1(_18757_),
    .B2(_04101_),
    .C1(_04321_),
    .X(_01921_));
 sky130_fd_sc_hd__buf_1 _26010_ (.A(_18199_),
    .X(_04322_));
 sky130_fd_sc_hd__buf_1 _26011_ (.A(_04120_),
    .X(_04323_));
 sky130_fd_sc_hd__nand2_2 _26012_ (.A(\cpuregs_rs1[16] ),
    .B(_04323_),
    .Y(_04324_));
 sky130_fd_sc_hd__o221a_2 _26013_ (.A1(_18304_),
    .A2(_04322_),
    .B1(_04118_),
    .B2(_20075_),
    .C1(_04324_),
    .X(_01923_));
 sky130_fd_sc_hd__nor2_2 _26014_ (.A(_20235_),
    .B(_20116_),
    .Y(_04325_));
 sky130_fd_sc_hd__inv_2 _26015_ (.A(_04325_),
    .Y(_04326_));
 sky130_fd_sc_hd__nand2_2 _26016_ (.A(_20235_),
    .B(_20116_),
    .Y(_04327_));
 sky130_fd_sc_hd__nand2_2 _26017_ (.A(_04326_),
    .B(_04327_),
    .Y(_04328_));
 sky130_fd_sc_hd__nor2_2 _26018_ (.A(_04313_),
    .B(_04317_),
    .Y(_04329_));
 sky130_fd_sc_hd__nor2_2 _26019_ (.A(_04328_),
    .B(_04329_),
    .Y(_04330_));
 sky130_fd_sc_hd__inv_2 _26020_ (.A(_04330_),
    .Y(_04331_));
 sky130_fd_sc_hd__nand2_2 _26021_ (.A(_04329_),
    .B(_04328_),
    .Y(_04332_));
 sky130_fd_sc_hd__a2bb2o_2 _26022_ (.A1_N(_01924_),
    .A2_N(_04194_),
    .B1(_19851_),
    .B2(_01919_),
    .X(_04333_));
 sky130_fd_sc_hd__nor2_2 _26023_ (.A(_01918_),
    .B(_04179_),
    .Y(_04334_));
 sky130_fd_sc_hd__a311o_2 _26024_ (.A1(_04331_),
    .A2(_04294_),
    .A3(_04332_),
    .B1(_04333_),
    .C1(_04334_),
    .X(_01925_));
 sky130_fd_sc_hd__nand2_2 _26025_ (.A(_01683_),
    .B(mem_rdata[17]),
    .Y(_01926_));
 sky130_fd_sc_hd__nand2_2 _26026_ (.A(\count_instr[49] ),
    .B(_04157_),
    .Y(_04335_));
 sky130_fd_sc_hd__o221a_2 _26027_ (.A1(_18748_),
    .A2(_04298_),
    .B1(_04198_),
    .B2(_18974_),
    .C1(_04335_),
    .X(_01930_));
 sky130_fd_sc_hd__buf_1 _26028_ (.A(_19438_),
    .X(_04336_));
 sky130_fd_sc_hd__a22o_2 _26029_ (.A1(\irq_mask[17] ),
    .A2(_04248_),
    .B1(_04336_),
    .B2(\timer[17] ),
    .X(_04337_));
 sky130_fd_sc_hd__a21oi_2 _26030_ (.A1(\cpuregs_rs1[17] ),
    .A2(_04261_),
    .B1(_04337_),
    .Y(_01932_));
 sky130_fd_sc_hd__nor2_2 _26031_ (.A(\reg_pc[17] ),
    .B(\decoded_imm[17] ),
    .Y(_04338_));
 sky130_fd_sc_hd__nor2_2 _26032_ (.A(_20242_),
    .B(_20118_),
    .Y(_04339_));
 sky130_fd_sc_hd__nor2_2 _26033_ (.A(_04338_),
    .B(_04339_),
    .Y(_04340_));
 sky130_fd_sc_hd__nand2_2 _26034_ (.A(_04331_),
    .B(_04326_),
    .Y(_04341_));
 sky130_fd_sc_hd__or2_2 _26035_ (.A(_04340_),
    .B(_04341_),
    .X(_04342_));
 sky130_fd_sc_hd__nand2_2 _26036_ (.A(_04341_),
    .B(_04340_),
    .Y(_04343_));
 sky130_fd_sc_hd__a2bb2o_2 _26037_ (.A1_N(_01933_),
    .A2_N(_04194_),
    .B1(_19851_),
    .B2(_01928_),
    .X(_04344_));
 sky130_fd_sc_hd__nor2_2 _26038_ (.A(_01927_),
    .B(_04179_),
    .Y(_04345_));
 sky130_fd_sc_hd__a311o_2 _26039_ (.A1(_04342_),
    .A2(_04343_),
    .A3(_04139_),
    .B1(_04344_),
    .C1(_04345_),
    .X(_01934_));
 sky130_fd_sc_hd__nand2_2 _26040_ (.A(_01683_),
    .B(mem_rdata[18]),
    .Y(_01935_));
 sky130_fd_sc_hd__nand2_2 _26041_ (.A(\count_instr[50] ),
    .B(_04157_),
    .Y(_04346_));
 sky130_fd_sc_hd__o221a_2 _26042_ (.A1(_18752_),
    .A2(_04298_),
    .B1(_04198_),
    .B2(_18965_),
    .C1(_04346_),
    .X(_01939_));
 sky130_fd_sc_hd__buf_1 _26043_ (.A(_18197_),
    .X(_04347_));
 sky130_fd_sc_hd__nand2_2 _26044_ (.A(\cpuregs_rs1[18] ),
    .B(_04323_),
    .Y(_04348_));
 sky130_fd_sc_hd__o221a_2 _26045_ (.A1(_18094_),
    .A2(_04322_),
    .B1(_04347_),
    .B2(_20044_),
    .C1(_04348_),
    .X(_01941_));
 sky130_fd_sc_hd__nor2_2 _26046_ (.A(\reg_pc[18] ),
    .B(_20119_),
    .Y(_04349_));
 sky130_fd_sc_hd__nor2_2 _26047_ (.A(\decoded_imm[18] ),
    .B(_20248_),
    .Y(_04350_));
 sky130_fd_sc_hd__o21ba_2 _26048_ (.A1(_04338_),
    .A2(_04326_),
    .B1_N(_04339_),
    .X(_04351_));
 sky130_fd_sc_hd__inv_2 _26049_ (.A(_04351_),
    .Y(_04352_));
 sky130_fd_sc_hd__o22ai_2 _26050_ (.A1(\reg_pc[15] ),
    .A2(\decoded_imm[15] ),
    .B1(_04302_),
    .B2(_04315_),
    .Y(_04353_));
 sky130_fd_sc_hd__inv_2 _26051_ (.A(_04313_),
    .Y(_04354_));
 sky130_fd_sc_hd__or3_2 _26052_ (.A(_04338_),
    .B(_04339_),
    .C(_04328_),
    .X(_04355_));
 sky130_fd_sc_hd__a21oi_2 _26053_ (.A1(_04353_),
    .A2(_04354_),
    .B1(_04355_),
    .Y(_04356_));
 sky130_fd_sc_hd__or4_2 _26054_ (.A(_04349_),
    .B(_04350_),
    .C(_04352_),
    .D(_04356_),
    .X(_04357_));
 sky130_fd_sc_hd__o22ai_2 _26055_ (.A1(_04349_),
    .A2(_04350_),
    .B1(_04352_),
    .B2(_04356_),
    .Y(_04358_));
 sky130_fd_sc_hd__o22ai_2 _26056_ (.A1(_01936_),
    .A2(_18444_),
    .B1(_19188_),
    .B2(_01942_),
    .Y(_04359_));
 sky130_fd_sc_hd__a21o_2 _26057_ (.A1(_19852_),
    .A2(_01937_),
    .B1(_04359_),
    .X(_04360_));
 sky130_fd_sc_hd__a31o_2 _26058_ (.A1(_04357_),
    .A2(_04108_),
    .A3(_04358_),
    .B1(_04360_),
    .X(_01943_));
 sky130_fd_sc_hd__nand2_2 _26059_ (.A(_01683_),
    .B(mem_rdata[19]),
    .Y(_01944_));
 sky130_fd_sc_hd__inv_2 _26060_ (.A(\count_cycle[19] ),
    .Y(_01947_));
 sky130_fd_sc_hd__buf_1 _26061_ (.A(_04100_),
    .X(_04361_));
 sky130_fd_sc_hd__nand2_2 _26062_ (.A(_04320_),
    .B(\count_cycle[51] ),
    .Y(_04362_));
 sky130_fd_sc_hd__o221a_2 _26063_ (.A1(_18672_),
    .A2(_04283_),
    .B1(_18615_),
    .B2(_04361_),
    .C1(_04362_),
    .X(_01948_));
 sky130_fd_sc_hd__nand2_2 _26064_ (.A(\cpuregs_rs1[19] ),
    .B(_04323_),
    .Y(_04363_));
 sky130_fd_sc_hd__o221a_2 _26065_ (.A1(_18092_),
    .A2(_04322_),
    .B1(_04347_),
    .B2(_20043_),
    .C1(_04363_),
    .X(_01950_));
 sky130_fd_sc_hd__nand2_2 _26066_ (.A(_20257_),
    .B(\decoded_imm[19] ),
    .Y(_04364_));
 sky130_fd_sc_hd__nand2_2 _26067_ (.A(_20120_),
    .B(\reg_pc[19] ),
    .Y(_04365_));
 sky130_fd_sc_hd__nand2_2 _26068_ (.A(\reg_pc[18] ),
    .B(\decoded_imm[18] ),
    .Y(_04366_));
 sky130_fd_sc_hd__a22oi_2 _26069_ (.A1(_04364_),
    .A2(_04365_),
    .B1(_04358_),
    .B2(_04366_),
    .Y(_04367_));
 sky130_fd_sc_hd__and4_2 _26070_ (.A(_04358_),
    .B(_04366_),
    .C(_04364_),
    .D(_04365_),
    .X(_04368_));
 sky130_fd_sc_hd__o22a_2 _26071_ (.A1(_01945_),
    .A2(_18444_),
    .B1(_18851_),
    .B2(_01951_),
    .X(_04369_));
 sky130_fd_sc_hd__nand2_2 _26072_ (.A(_19852_),
    .B(_01946_),
    .Y(_04370_));
 sky130_fd_sc_hd__o311ai_2 _26073_ (.A1(_18187_),
    .A2(_04367_),
    .A3(_04368_),
    .B1(_04369_),
    .C1(_04370_),
    .Y(_01952_));
 sky130_fd_sc_hd__nand2_2 _26074_ (.A(_01683_),
    .B(mem_rdata[20]),
    .Y(_01953_));
 sky130_fd_sc_hd__nand2_2 _26075_ (.A(\count_instr[52] ),
    .B(_04169_),
    .Y(_04371_));
 sky130_fd_sc_hd__o221a_2 _26076_ (.A1(_18614_),
    .A2(_04298_),
    .B1(_04197_),
    .B2(_18931_),
    .C1(_04371_),
    .X(_01957_));
 sky130_fd_sc_hd__buf_1 _26077_ (.A(_18198_),
    .X(_04372_));
 sky130_fd_sc_hd__a22o_2 _26078_ (.A1(\irq_mask[20] ),
    .A2(_04372_),
    .B1(_04336_),
    .B2(\timer[20] ),
    .X(_04373_));
 sky130_fd_sc_hd__a21oi_2 _26079_ (.A1(\cpuregs_rs1[20] ),
    .A2(_04261_),
    .B1(_04373_),
    .Y(_01959_));
 sky130_fd_sc_hd__nor2_2 _26080_ (.A(_20263_),
    .B(_20121_),
    .Y(_04374_));
 sky130_fd_sc_hd__inv_2 _26081_ (.A(_04374_),
    .Y(_04375_));
 sky130_fd_sc_hd__nand2_2 _26082_ (.A(_20263_),
    .B(_20121_),
    .Y(_04376_));
 sky130_fd_sc_hd__nand2_2 _26083_ (.A(_04375_),
    .B(_04376_),
    .Y(_04377_));
 sky130_fd_sc_hd__nor2_2 _26084_ (.A(_20257_),
    .B(_20120_),
    .Y(_04378_));
 sky130_fd_sc_hd__or2_2 _26085_ (.A(_04378_),
    .B(_04367_),
    .X(_04379_));
 sky130_fd_sc_hd__inv_2 _26086_ (.A(_04379_),
    .Y(_04380_));
 sky130_fd_sc_hd__or2_2 _26087_ (.A(_04377_),
    .B(_04380_),
    .X(_04381_));
 sky130_fd_sc_hd__nand2_2 _26088_ (.A(_04380_),
    .B(_04377_),
    .Y(_04382_));
 sky130_fd_sc_hd__o22a_2 _26089_ (.A1(_01954_),
    .A2(_04111_),
    .B1(_19771_),
    .B2(_01960_),
    .X(_04383_));
 sky130_fd_sc_hd__a21bo_2 _26090_ (.A1(_04129_),
    .A2(_01955_),
    .B1_N(_04383_),
    .X(_04384_));
 sky130_fd_sc_hd__a31o_2 _26091_ (.A1(_04381_),
    .A2(_04108_),
    .A3(_04382_),
    .B1(_04384_),
    .X(_01961_));
 sky130_fd_sc_hd__buf_1 _26092_ (.A(_04085_),
    .X(_04385_));
 sky130_fd_sc_hd__nand2_2 _26093_ (.A(_04385_),
    .B(mem_rdata[21]),
    .Y(_01962_));
 sky130_fd_sc_hd__a22o_2 _26094_ (.A1(\count_instr[53] ),
    .A2(instr_rdinstrh),
    .B1(_04246_),
    .B2(\count_cycle[53] ),
    .X(_04386_));
 sky130_fd_sc_hd__a21oi_2 _26095_ (.A1(\count_instr[21] ),
    .A2(_19478_),
    .B1(_04386_),
    .Y(_01966_));
 sky130_fd_sc_hd__buf_1 _26096_ (.A(_04120_),
    .X(_04387_));
 sky130_fd_sc_hd__a22o_2 _26097_ (.A1(\irq_mask[21] ),
    .A2(_04372_),
    .B1(_04336_),
    .B2(\timer[21] ),
    .X(_04388_));
 sky130_fd_sc_hd__a21oi_2 _26098_ (.A1(\cpuregs_rs1[21] ),
    .A2(_04387_),
    .B1(_04388_),
    .Y(_01968_));
 sky130_fd_sc_hd__nor2_2 _26099_ (.A(_20272_),
    .B(_20122_),
    .Y(_04389_));
 sky130_fd_sc_hd__inv_2 _26100_ (.A(_04389_),
    .Y(_04390_));
 sky130_fd_sc_hd__nand2_2 _26101_ (.A(_20272_),
    .B(_20122_),
    .Y(_04391_));
 sky130_fd_sc_hd__nand2_2 _26102_ (.A(_04390_),
    .B(_04391_),
    .Y(_04392_));
 sky130_fd_sc_hd__o22ai_2 _26103_ (.A1(\reg_pc[20] ),
    .A2(\decoded_imm[20] ),
    .B1(_04378_),
    .B2(_04367_),
    .Y(_04393_));
 sky130_fd_sc_hd__nand2_2 _26104_ (.A(_04393_),
    .B(_04375_),
    .Y(_04394_));
 sky130_fd_sc_hd__inv_2 _26105_ (.A(_04394_),
    .Y(_04395_));
 sky130_fd_sc_hd__o21a_2 _26106_ (.A1(_04392_),
    .A2(_04395_),
    .B1(_04294_),
    .X(_04396_));
 sky130_fd_sc_hd__nand2_2 _26107_ (.A(_04395_),
    .B(_04392_),
    .Y(_04397_));
 sky130_fd_sc_hd__o22ai_2 _26108_ (.A1(_01963_),
    .A2(_04112_),
    .B1(_04232_),
    .B2(_01969_),
    .Y(_04398_));
 sky130_fd_sc_hd__a221o_2 _26109_ (.A1(_04202_),
    .A2(_01964_),
    .B1(_04396_),
    .B2(_04397_),
    .C1(_04398_),
    .X(_01970_));
 sky130_fd_sc_hd__nand2_2 _26110_ (.A(_04385_),
    .B(mem_rdata[22]),
    .Y(_01971_));
 sky130_fd_sc_hd__nand2_2 _26111_ (.A(_04320_),
    .B(\count_cycle[54] ),
    .Y(_04399_));
 sky130_fd_sc_hd__o221a_2 _26112_ (.A1(_18662_),
    .A2(_04283_),
    .B1(_18733_),
    .B2(_04361_),
    .C1(_04399_),
    .X(_01975_));
 sky130_fd_sc_hd__a22o_2 _26113_ (.A1(\irq_mask[22] ),
    .A2(_04372_),
    .B1(_04336_),
    .B2(\timer[22] ),
    .X(_04400_));
 sky130_fd_sc_hd__a21oi_2 _26114_ (.A1(\cpuregs_rs1[22] ),
    .A2(_04387_),
    .B1(_04400_),
    .Y(_01977_));
 sky130_fd_sc_hd__nor2_2 _26115_ (.A(_20277_),
    .B(_20123_),
    .Y(_04401_));
 sky130_fd_sc_hd__inv_2 _26116_ (.A(_04401_),
    .Y(_04402_));
 sky130_fd_sc_hd__nor2_2 _26117_ (.A(\reg_pc[22] ),
    .B(\decoded_imm[22] ),
    .Y(_04403_));
 sky130_fd_sc_hd__inv_2 _26118_ (.A(_04403_),
    .Y(_04404_));
 sky130_fd_sc_hd__nand2_2 _26119_ (.A(_04402_),
    .B(_04404_),
    .Y(_04405_));
 sky130_fd_sc_hd__a22oi_2 _26120_ (.A1(_20272_),
    .A2(_20122_),
    .B1(_04393_),
    .B2(_04375_),
    .Y(_04406_));
 sky130_fd_sc_hd__inv_2 _26121_ (.A(_04406_),
    .Y(_04407_));
 sky130_fd_sc_hd__nand2_2 _26122_ (.A(_04407_),
    .B(_04390_),
    .Y(_04408_));
 sky130_fd_sc_hd__inv_2 _26123_ (.A(_04408_),
    .Y(_04409_));
 sky130_fd_sc_hd__or2_2 _26124_ (.A(_04405_),
    .B(_04409_),
    .X(_04410_));
 sky130_fd_sc_hd__nand2_2 _26125_ (.A(_04409_),
    .B(_04405_),
    .Y(_04411_));
 sky130_fd_sc_hd__o22a_2 _26126_ (.A1(_01972_),
    .A2(_18205_),
    .B1(_18194_),
    .B2(_01978_),
    .X(_04412_));
 sky130_fd_sc_hd__a21bo_2 _26127_ (.A1(_04129_),
    .A2(_01973_),
    .B1_N(_04412_),
    .X(_04413_));
 sky130_fd_sc_hd__a31o_2 _26128_ (.A1(_04410_),
    .A2(_04108_),
    .A3(_04411_),
    .B1(_04413_),
    .X(_01979_));
 sky130_fd_sc_hd__nand2_2 _26129_ (.A(_04385_),
    .B(mem_rdata[23]),
    .Y(_01980_));
 sky130_fd_sc_hd__a22o_2 _26130_ (.A1(\count_instr[23] ),
    .A2(instr_rdinstr),
    .B1(_04246_),
    .B2(\count_cycle[55] ),
    .X(_04414_));
 sky130_fd_sc_hd__a21oi_2 _26131_ (.A1(\count_instr[55] ),
    .A2(_19474_),
    .B1(_04414_),
    .Y(_01984_));
 sky130_fd_sc_hd__a22o_2 _26132_ (.A1(\irq_mask[23] ),
    .A2(_04372_),
    .B1(_04336_),
    .B2(\timer[23] ),
    .X(_04415_));
 sky130_fd_sc_hd__a21oi_2 _26133_ (.A1(\cpuregs_rs1[23] ),
    .A2(_04387_),
    .B1(_04415_),
    .Y(_01986_));
 sky130_fd_sc_hd__nor2_2 _26134_ (.A(\reg_pc[23] ),
    .B(\decoded_imm[23] ),
    .Y(_04416_));
 sky130_fd_sc_hd__nor2_2 _26135_ (.A(_20286_),
    .B(_20125_),
    .Y(_04417_));
 sky130_fd_sc_hd__or2_2 _26136_ (.A(_04416_),
    .B(_04417_),
    .X(_04418_));
 sky130_fd_sc_hd__o22ai_2 _26137_ (.A1(\reg_pc[22] ),
    .A2(\decoded_imm[22] ),
    .B1(_04389_),
    .B2(_04406_),
    .Y(_04419_));
 sky130_fd_sc_hd__and2_2 _26138_ (.A(_04419_),
    .B(_04402_),
    .X(_04420_));
 sky130_fd_sc_hd__o21a_2 _26139_ (.A1(_04418_),
    .A2(_04420_),
    .B1(_04294_),
    .X(_04421_));
 sky130_fd_sc_hd__nand2_2 _26140_ (.A(_04420_),
    .B(_04418_),
    .Y(_04422_));
 sky130_fd_sc_hd__buf_1 _26141_ (.A(_18205_),
    .X(_04423_));
 sky130_fd_sc_hd__o22ai_2 _26142_ (.A1(_01981_),
    .A2(_04423_),
    .B1(_18800_),
    .B2(_01987_),
    .Y(_04424_));
 sky130_fd_sc_hd__a221o_2 _26143_ (.A1(_04202_),
    .A2(_01982_),
    .B1(_04421_),
    .B2(_04422_),
    .C1(_04424_),
    .X(_01988_));
 sky130_fd_sc_hd__nand2_2 _26144_ (.A(_04385_),
    .B(mem_rdata[24]),
    .Y(_01989_));
 sky130_fd_sc_hd__nand2_2 _26145_ (.A(_04320_),
    .B(\count_cycle[56] ),
    .Y(_04425_));
 sky130_fd_sc_hd__o221a_2 _26146_ (.A1(_18654_),
    .A2(_04283_),
    .B1(_18738_),
    .B2(_04361_),
    .C1(_04425_),
    .X(_01993_));
 sky130_fd_sc_hd__nand2_2 _26147_ (.A(\cpuregs_rs1[24] ),
    .B(_04323_),
    .Y(_04426_));
 sky130_fd_sc_hd__o221a_2 _26148_ (.A1(_18100_),
    .A2(_04322_),
    .B1(_04347_),
    .B2(_20091_),
    .C1(_04426_),
    .X(_01995_));
 sky130_fd_sc_hd__nand2_2 _26149_ (.A(_20291_),
    .B(_20126_),
    .Y(_04427_));
 sky130_fd_sc_hd__nand2_2 _26150_ (.A(\reg_pc[24] ),
    .B(\decoded_imm[24] ),
    .Y(_04428_));
 sky130_fd_sc_hd__nand2_2 _26151_ (.A(_04427_),
    .B(_04428_),
    .Y(_04429_));
 sky130_fd_sc_hd__a22oi_2 _26152_ (.A1(_20286_),
    .A2(_20125_),
    .B1(_04419_),
    .B2(_04402_),
    .Y(_04430_));
 sky130_fd_sc_hd__nor2_2 _26153_ (.A(_04417_),
    .B(_04430_),
    .Y(_04431_));
 sky130_fd_sc_hd__or2_2 _26154_ (.A(_04429_),
    .B(_04431_),
    .X(_04432_));
 sky130_fd_sc_hd__nand2_2 _26155_ (.A(_04431_),
    .B(_04429_),
    .Y(_04433_));
 sky130_fd_sc_hd__o22ai_2 _26156_ (.A1(_01990_),
    .A2(_18444_),
    .B1(_19188_),
    .B2(_01996_),
    .Y(_04434_));
 sky130_fd_sc_hd__a21o_2 _26157_ (.A1(_19852_),
    .A2(_01991_),
    .B1(_04434_),
    .X(_04435_));
 sky130_fd_sc_hd__a31o_2 _26158_ (.A1(_04432_),
    .A2(_04108_),
    .A3(_04433_),
    .B1(_04435_),
    .X(_01997_));
 sky130_fd_sc_hd__nand2_2 _26159_ (.A(_04385_),
    .B(mem_rdata[25]),
    .Y(_01998_));
 sky130_fd_sc_hd__nand2_2 _26160_ (.A(_04320_),
    .B(\count_cycle[57] ),
    .Y(_04436_));
 sky130_fd_sc_hd__o221a_2 _26161_ (.A1(_18653_),
    .A2(_04283_),
    .B1(_18592_),
    .B2(_04361_),
    .C1(_04436_),
    .X(_02002_));
 sky130_fd_sc_hd__a22o_2 _26162_ (.A1(\irq_mask[25] ),
    .A2(_04372_),
    .B1(_04336_),
    .B2(\timer[25] ),
    .X(_04437_));
 sky130_fd_sc_hd__a21oi_2 _26163_ (.A1(\cpuregs_rs1[25] ),
    .A2(_04387_),
    .B1(_04437_),
    .Y(_02004_));
 sky130_fd_sc_hd__nor2_2 _26164_ (.A(\reg_pc[25] ),
    .B(\decoded_imm[25] ),
    .Y(_04438_));
 sky130_fd_sc_hd__nor2_2 _26165_ (.A(_20297_),
    .B(_20127_),
    .Y(_04439_));
 sky130_fd_sc_hd__or2_2 _26166_ (.A(_04438_),
    .B(_04439_),
    .X(_04440_));
 sky130_fd_sc_hd__a21o_2 _26167_ (.A1(_04432_),
    .A2(_04428_),
    .B1(_04440_),
    .X(_04441_));
 sky130_fd_sc_hd__a31oi_2 _26168_ (.A1(_04432_),
    .A2(_04428_),
    .A3(_04440_),
    .B1(_18187_),
    .Y(_04442_));
 sky130_fd_sc_hd__o22ai_2 _26169_ (.A1(_01999_),
    .A2(_04423_),
    .B1(_18800_),
    .B2(_02005_),
    .Y(_04443_));
 sky130_fd_sc_hd__a221o_2 _26170_ (.A1(_04202_),
    .A2(_02000_),
    .B1(_04441_),
    .B2(_04442_),
    .C1(_04443_),
    .X(_02006_));
 sky130_fd_sc_hd__nand2_2 _26171_ (.A(_04385_),
    .B(mem_rdata[26]),
    .Y(_02007_));
 sky130_fd_sc_hd__nand2_2 _26172_ (.A(\count_instr[58] ),
    .B(_04169_),
    .Y(_04444_));
 sky130_fd_sc_hd__o221a_2 _26173_ (.A1(_18591_),
    .A2(_04298_),
    .B1(_04197_),
    .B2(_18887_),
    .C1(_04444_),
    .X(_02011_));
 sky130_fd_sc_hd__a22o_2 _26174_ (.A1(\irq_mask[26] ),
    .A2(_04372_),
    .B1(_19438_),
    .B2(\timer[26] ),
    .X(_04445_));
 sky130_fd_sc_hd__a21oi_2 _26175_ (.A1(\cpuregs_rs1[26] ),
    .A2(_04387_),
    .B1(_04445_),
    .Y(_02013_));
 sky130_fd_sc_hd__o2bb2a_2 _26176_ (.A1_N(_04193_),
    .A2_N(_02009_),
    .B1(_02014_),
    .B2(_19188_),
    .X(_04446_));
 sky130_fd_sc_hd__or2_2 _26177_ (.A(_04429_),
    .B(_04440_),
    .X(_04447_));
 sky130_fd_sc_hd__o21bai_2 _26178_ (.A1(_04417_),
    .A2(_04430_),
    .B1_N(_04447_),
    .Y(_04448_));
 sky130_fd_sc_hd__o21ba_2 _26179_ (.A1(_04428_),
    .A2(_04438_),
    .B1_N(_04439_),
    .X(_04449_));
 sky130_fd_sc_hd__nor2_2 _26180_ (.A(_20303_),
    .B(_20128_),
    .Y(_04450_));
 sky130_fd_sc_hd__inv_2 _26181_ (.A(_04450_),
    .Y(_04451_));
 sky130_fd_sc_hd__nand2_2 _26182_ (.A(_20303_),
    .B(_20128_),
    .Y(_04452_));
 sky130_fd_sc_hd__nand2_2 _26183_ (.A(_04451_),
    .B(_04452_),
    .Y(_04453_));
 sky130_fd_sc_hd__a21oi_2 _26184_ (.A1(_04448_),
    .A2(_04449_),
    .B1(_04453_),
    .Y(_04454_));
 sky130_fd_sc_hd__and3_2 _26185_ (.A(_04448_),
    .B(_04449_),
    .C(_04453_),
    .X(_04455_));
 sky130_fd_sc_hd__or3_2 _26186_ (.A(_18186_),
    .B(_04454_),
    .C(_04455_),
    .X(_04456_));
 sky130_fd_sc_hd__o211ai_2 _26187_ (.A1(_20006_),
    .A2(_02008_),
    .B1(_04446_),
    .C1(_04456_),
    .Y(_02015_));
 sky130_fd_sc_hd__buf_1 _26188_ (.A(_04085_),
    .X(_04457_));
 sky130_fd_sc_hd__nand2_2 _26189_ (.A(_04457_),
    .B(mem_rdata[27]),
    .Y(_02016_));
 sky130_fd_sc_hd__nand2_2 _26190_ (.A(_04320_),
    .B(\count_cycle[59] ),
    .Y(_04458_));
 sky130_fd_sc_hd__o221a_2 _26191_ (.A1(_18580_),
    .A2(_04098_),
    .B1(_18620_),
    .B2(_04361_),
    .C1(_04458_),
    .X(_02020_));
 sky130_fd_sc_hd__a22o_2 _26192_ (.A1(\irq_mask[27] ),
    .A2(_18198_),
    .B1(_19438_),
    .B2(\timer[27] ),
    .X(_04459_));
 sky130_fd_sc_hd__a21oi_2 _26193_ (.A1(\cpuregs_rs1[27] ),
    .A2(_04387_),
    .B1(_04459_),
    .Y(_02022_));
 sky130_fd_sc_hd__nor2_2 _26194_ (.A(\reg_pc[27] ),
    .B(\decoded_imm[27] ),
    .Y(_04460_));
 sky130_fd_sc_hd__nor2_2 _26195_ (.A(_20312_),
    .B(_20129_),
    .Y(_04461_));
 sky130_fd_sc_hd__nor2_2 _26196_ (.A(_04460_),
    .B(_04461_),
    .Y(_04462_));
 sky130_fd_sc_hd__or2_2 _26197_ (.A(_04450_),
    .B(_04454_),
    .X(_04463_));
 sky130_fd_sc_hd__or2_2 _26198_ (.A(_04462_),
    .B(_04463_),
    .X(_04464_));
 sky130_fd_sc_hd__nand2_2 _26199_ (.A(_04463_),
    .B(_04462_),
    .Y(_04465_));
 sky130_fd_sc_hd__o2bb2a_2 _26200_ (.A1_N(_19851_),
    .A2_N(_02018_),
    .B1(_02023_),
    .B2(_18799_),
    .X(_04466_));
 sky130_fd_sc_hd__o21ai_2 _26201_ (.A1(_04112_),
    .A2(_02017_),
    .B1(_04466_),
    .Y(_04467_));
 sky130_fd_sc_hd__a31o_2 _26202_ (.A1(_04464_),
    .A2(_04108_),
    .A3(_04465_),
    .B1(_04467_),
    .X(_02024_));
 sky130_fd_sc_hd__nand2_2 _26203_ (.A(_04457_),
    .B(mem_rdata[28]),
    .Y(_02025_));
 sky130_fd_sc_hd__nand2_2 _26204_ (.A(_04246_),
    .B(\count_cycle[60] ),
    .Y(_04468_));
 sky130_fd_sc_hd__o221a_2 _26205_ (.A1(_18579_),
    .A2(_04098_),
    .B1(_18624_),
    .B2(_04361_),
    .C1(_04468_),
    .X(_02029_));
 sky130_fd_sc_hd__nand2_2 _26206_ (.A(\cpuregs_rs1[28] ),
    .B(_04323_),
    .Y(_04469_));
 sky130_fd_sc_hd__o221a_2 _26207_ (.A1(_18127_),
    .A2(_04322_),
    .B1(_04347_),
    .B2(_20098_),
    .C1(_04469_),
    .X(_02031_));
 sky130_fd_sc_hd__nor2_2 _26208_ (.A(\reg_pc[28] ),
    .B(\decoded_imm[28] ),
    .Y(_04470_));
 sky130_fd_sc_hd__nor2_2 _26209_ (.A(_20317_),
    .B(_20130_),
    .Y(_04471_));
 sky130_fd_sc_hd__nor2_2 _26210_ (.A(_04470_),
    .B(_04471_),
    .Y(_04472_));
 sky130_fd_sc_hd__o21ba_2 _26211_ (.A1(_04460_),
    .A2(_04451_),
    .B1_N(_04461_),
    .X(_04473_));
 sky130_fd_sc_hd__inv_2 _26212_ (.A(_04473_),
    .Y(_04474_));
 sky130_fd_sc_hd__or3_2 _26213_ (.A(_04460_),
    .B(_04461_),
    .C(_04453_),
    .X(_04475_));
 sky130_fd_sc_hd__a21oi_2 _26214_ (.A1(_04448_),
    .A2(_04449_),
    .B1(_04475_),
    .Y(_04476_));
 sky130_fd_sc_hd__or2_2 _26215_ (.A(_04474_),
    .B(_04476_),
    .X(_04477_));
 sky130_fd_sc_hd__or2_2 _26216_ (.A(_04472_),
    .B(_04477_),
    .X(_04478_));
 sky130_fd_sc_hd__nand2_2 _26217_ (.A(_04477_),
    .B(_04472_),
    .Y(_04479_));
 sky130_fd_sc_hd__o22ai_2 _26218_ (.A1(_02026_),
    .A2(_04423_),
    .B1(_18800_),
    .B2(_02032_),
    .Y(_04480_));
 sky130_fd_sc_hd__and2_2 _26219_ (.A(_04114_),
    .B(_02027_),
    .X(_04481_));
 sky130_fd_sc_hd__a311o_2 _26220_ (.A1(_04478_),
    .A2(_04294_),
    .A3(_04479_),
    .B1(_04480_),
    .C1(_04481_),
    .X(_02033_));
 sky130_fd_sc_hd__nand2_2 _26221_ (.A(_04457_),
    .B(mem_rdata[29]),
    .Y(_02034_));
 sky130_fd_sc_hd__nand2_2 _26222_ (.A(\count_instr[61] ),
    .B(_04169_),
    .Y(_04482_));
 sky130_fd_sc_hd__o221a_2 _26223_ (.A1(_18623_),
    .A2(_04298_),
    .B1(_04197_),
    .B2(_18891_),
    .C1(_04482_),
    .X(_02038_));
 sky130_fd_sc_hd__a22o_2 _26224_ (.A1(\irq_mask[29] ),
    .A2(_18198_),
    .B1(_19438_),
    .B2(\timer[29] ),
    .X(_04483_));
 sky130_fd_sc_hd__a21oi_2 _26225_ (.A1(\cpuregs_rs1[29] ),
    .A2(_04121_),
    .B1(_04483_),
    .Y(_02040_));
 sky130_fd_sc_hd__o22ai_2 _26226_ (.A1(\reg_pc[28] ),
    .A2(\decoded_imm[28] ),
    .B1(_04474_),
    .B2(_04476_),
    .Y(_04484_));
 sky130_fd_sc_hd__inv_2 _26227_ (.A(_04471_),
    .Y(_04485_));
 sky130_fd_sc_hd__nor2_2 _26228_ (.A(\reg_pc[29] ),
    .B(\decoded_imm[29] ),
    .Y(_04486_));
 sky130_fd_sc_hd__nor2_2 _26229_ (.A(_20327_),
    .B(_20131_),
    .Y(_04487_));
 sky130_fd_sc_hd__or2_2 _26230_ (.A(_04486_),
    .B(_04487_),
    .X(_04488_));
 sky130_fd_sc_hd__a21oi_2 _26231_ (.A1(_04484_),
    .A2(_04485_),
    .B1(_04488_),
    .Y(_04489_));
 sky130_fd_sc_hd__a31o_2 _26232_ (.A1(_04484_),
    .A2(_04485_),
    .A3(_04488_),
    .B1(_18186_),
    .X(_04490_));
 sky130_fd_sc_hd__o22a_2 _26233_ (.A1(_02035_),
    .A2(_04423_),
    .B1(_18806_),
    .B2(_02041_),
    .X(_04491_));
 sky130_fd_sc_hd__nand2_2 _26234_ (.A(_19852_),
    .B(_02036_),
    .Y(_04492_));
 sky130_fd_sc_hd__o211ai_2 _26235_ (.A1(_04489_),
    .A2(_04490_),
    .B1(_04491_),
    .C1(_04492_),
    .Y(_02042_));
 sky130_fd_sc_hd__nand2_2 _26236_ (.A(_04457_),
    .B(mem_rdata[30]),
    .Y(_02043_));
 sky130_fd_sc_hd__nand2_2 _26237_ (.A(\count_instr[30] ),
    .B(_19478_),
    .Y(_04493_));
 sky130_fd_sc_hd__o221a_2 _26238_ (.A1(_18578_),
    .A2(_04098_),
    .B1(_04197_),
    .B2(_18889_),
    .C1(_04493_),
    .X(_02047_));
 sky130_fd_sc_hd__inv_2 _26239_ (.A(\timer[30] ),
    .Y(_04494_));
 sky130_fd_sc_hd__nand2_2 _26240_ (.A(\cpuregs_rs1[30] ),
    .B(_04323_),
    .Y(_04495_));
 sky130_fd_sc_hd__o221a_2 _26241_ (.A1(_18131_),
    .A2(_04322_),
    .B1(_04347_),
    .B2(_04494_),
    .C1(_04495_),
    .X(_02049_));
 sky130_fd_sc_hd__a21o_2 _26242_ (.A1(_04484_),
    .A2(_04485_),
    .B1(_04486_),
    .X(_04496_));
 sky130_fd_sc_hd__nor2_2 _26243_ (.A(\reg_pc[30] ),
    .B(_20132_),
    .Y(_04497_));
 sky130_fd_sc_hd__nor2_2 _26244_ (.A(\decoded_imm[30] ),
    .B(_18505_),
    .Y(_04498_));
 sky130_fd_sc_hd__nor2_2 _26245_ (.A(_04497_),
    .B(_04498_),
    .Y(_04499_));
 sky130_fd_sc_hd__nand3b_2 _26246_ (.A_N(_04487_),
    .B(_04496_),
    .C(_04499_),
    .Y(_04500_));
 sky130_fd_sc_hd__a22oi_2 _26247_ (.A1(_20327_),
    .A2(_20131_),
    .B1(_04484_),
    .B2(_04485_),
    .Y(_04501_));
 sky130_fd_sc_hd__o22ai_2 _26248_ (.A1(_04497_),
    .A2(_04498_),
    .B1(_04487_),
    .B2(_04501_),
    .Y(_04502_));
 sky130_fd_sc_hd__nor2_2 _26249_ (.A(_02050_),
    .B(_04232_),
    .Y(_04503_));
 sky130_fd_sc_hd__a2bb2o_2 _26250_ (.A1_N(_02044_),
    .A2_N(_04423_),
    .B1(_04114_),
    .B2(_02045_),
    .X(_04504_));
 sky130_fd_sc_hd__a311o_2 _26251_ (.A1(_04500_),
    .A2(_04502_),
    .A3(_04139_),
    .B1(_04503_),
    .C1(_04504_),
    .X(_02051_));
 sky130_fd_sc_hd__nand2_2 _26252_ (.A(_04457_),
    .B(mem_rdata[31]),
    .Y(_02052_));
 sky130_fd_sc_hd__inv_2 _26253_ (.A(\count_cycle[31] ),
    .Y(_02055_));
 sky130_fd_sc_hd__nand2_2 _26254_ (.A(\count_instr[63] ),
    .B(_04169_),
    .Y(_04505_));
 sky130_fd_sc_hd__o221a_2 _26255_ (.A1(_18621_),
    .A2(_04100_),
    .B1(_04197_),
    .B2(_18936_),
    .C1(_04505_),
    .X(_02056_));
 sky130_fd_sc_hd__inv_2 _26256_ (.A(\timer[31] ),
    .Y(_04506_));
 sky130_fd_sc_hd__nand2_2 _26257_ (.A(\cpuregs_rs1[31] ),
    .B(_04120_),
    .Y(_04507_));
 sky130_fd_sc_hd__o221a_2 _26258_ (.A1(_18129_),
    .A2(_18199_),
    .B1(_04347_),
    .B2(_04506_),
    .C1(_04507_),
    .X(_02058_));
 sky130_fd_sc_hd__nand2_2 _26259_ (.A(\reg_pc[30] ),
    .B(\decoded_imm[30] ),
    .Y(_04508_));
 sky130_fd_sc_hd__xnor2_2 _26260_ (.A(\reg_pc[31] ),
    .B(\decoded_imm[31] ),
    .Y(_04509_));
 sky130_fd_sc_hd__a21oi_2 _26261_ (.A1(_04502_),
    .A2(_04508_),
    .B1(_04509_),
    .Y(_04510_));
 sky130_fd_sc_hd__nand3_2 _26262_ (.A(_04502_),
    .B(_04508_),
    .C(_04509_),
    .Y(_04511_));
 sky130_fd_sc_hd__nand2_2 _26263_ (.A(_04511_),
    .B(_04294_),
    .Y(_04512_));
 sky130_fd_sc_hd__nand2_2 _26264_ (.A(_04193_),
    .B(_02054_),
    .Y(_04513_));
 sky130_fd_sc_hd__o221ai_2 _26265_ (.A1(_02053_),
    .A2(_04423_),
    .B1(_02059_),
    .B2(_18800_),
    .C1(_04513_),
    .Y(_04514_));
 sky130_fd_sc_hd__o21bai_2 _26266_ (.A1(_04510_),
    .A2(_04512_),
    .B1_N(_04514_),
    .Y(_02060_));
 sky130_fd_sc_hd__or2_2 _26267_ (.A(\decoded_rd[4] ),
    .B(_00308_),
    .X(_02061_));
 sky130_fd_sc_hd__o21ai_2 _26268_ (.A1(_02064_),
    .A2(_18188_),
    .B1(_04232_),
    .Y(_02065_));
 sky130_fd_sc_hd__nor3_2 _26269_ (.A(_18150_),
    .B(_02410_),
    .C(_00308_),
    .Y(_02066_));
 sky130_fd_sc_hd__and3_2 _26270_ (.A(_18443_),
    .B(_18187_),
    .C(_20006_),
    .X(_02067_));
 sky130_fd_sc_hd__nand2_2 _26271_ (.A(_18338_),
    .B(_00343_),
    .Y(_04515_));
 sky130_fd_sc_hd__a211o_2 _26272_ (.A1(_04515_),
    .A2(_04127_),
    .B1(_18250_),
    .C1(_18029_),
    .X(_02068_));
 sky130_fd_sc_hd__nor2_2 _26273_ (.A(latched_branch),
    .B(_18230_),
    .Y(_04516_));
 sky130_fd_sc_hd__buf_1 _26274_ (.A(_04516_),
    .X(_04517_));
 sky130_fd_sc_hd__buf_1 _26275_ (.A(_04517_),
    .X(_04518_));
 sky130_fd_sc_hd__nor2_2 _26276_ (.A(_04518_),
    .B(_19075_),
    .Y(_02069_));
 sky130_fd_sc_hd__buf_1 _26277_ (.A(_18236_),
    .X(_04519_));
 sky130_fd_sc_hd__nor2_2 _26278_ (.A(_18232_),
    .B(_20135_),
    .Y(_04520_));
 sky130_fd_sc_hd__a221o_2 _26279_ (.A1(_18083_),
    .A2(_04519_),
    .B1(_04518_),
    .B2(_02070_),
    .C1(_04520_),
    .X(_02071_));
 sky130_fd_sc_hd__buf_1 _26280_ (.A(\irq_state[0] ),
    .X(_04521_));
 sky130_fd_sc_hd__and2_2 _26281_ (.A(_04521_),
    .B(\reg_next_pc[1] ),
    .X(_04522_));
 sky130_fd_sc_hd__a221o_2 _26282_ (.A1(_18085_),
    .A2(_04519_),
    .B1(_04518_),
    .B2(_01465_),
    .C1(_04522_),
    .X(_02072_));
 sky130_fd_sc_hd__buf_1 _26283_ (.A(_04517_),
    .X(_04523_));
 sky130_fd_sc_hd__and3_2 _26284_ (.A(_18081_),
    .B(_18236_),
    .C(\irq_pending[2] ),
    .X(_04524_));
 sky130_fd_sc_hd__a221o_2 _26285_ (.A1(_20347_),
    .A2(\reg_next_pc[2] ),
    .B1(_00293_),
    .B2(_04523_),
    .C1(_04524_),
    .X(_02074_));
 sky130_fd_sc_hd__nor2_2 _26286_ (.A(\reg_pc[3] ),
    .B(\reg_pc[2] ),
    .Y(_04525_));
 sky130_fd_sc_hd__nor2_2 _26287_ (.A(_20147_),
    .B(_02073_),
    .Y(_04526_));
 sky130_fd_sc_hd__nor2_2 _26288_ (.A(_04525_),
    .B(_04526_),
    .Y(_02075_));
 sky130_fd_sc_hd__and3_2 _26289_ (.A(_18086_),
    .B(_18236_),
    .C(\irq_pending[3] ),
    .X(_04527_));
 sky130_fd_sc_hd__a221o_2 _26290_ (.A1(_20347_),
    .A2(\reg_next_pc[3] ),
    .B1(_01468_),
    .B2(_04523_),
    .C1(_04527_),
    .X(_02076_));
 sky130_fd_sc_hd__nor2_2 _26291_ (.A(\reg_pc[4] ),
    .B(_04526_),
    .Y(_04528_));
 sky130_fd_sc_hd__nand2_2 _26292_ (.A(_04526_),
    .B(\reg_pc[4] ),
    .Y(_04529_));
 sky130_fd_sc_hd__inv_2 _26293_ (.A(_04529_),
    .Y(_04530_));
 sky130_fd_sc_hd__nor2_2 _26294_ (.A(_04528_),
    .B(_04530_),
    .Y(_02077_));
 sky130_fd_sc_hd__buf_1 _26295_ (.A(\irq_state[1] ),
    .X(_04531_));
 sky130_fd_sc_hd__buf_1 _26296_ (.A(_04531_),
    .X(_04532_));
 sky130_fd_sc_hd__and3_2 _26297_ (.A(_18123_),
    .B(_04532_),
    .C(\irq_pending[4] ),
    .X(_04533_));
 sky130_fd_sc_hd__a221o_2 _26298_ (.A1(_20347_),
    .A2(\reg_next_pc[4] ),
    .B1(_01472_),
    .B2(_04523_),
    .C1(_04533_),
    .X(_02078_));
 sky130_fd_sc_hd__nor2_2 _26299_ (.A(_20161_),
    .B(_04529_),
    .Y(_04534_));
 sky130_fd_sc_hd__nor2_2 _26300_ (.A(\reg_pc[5] ),
    .B(_04530_),
    .Y(_04535_));
 sky130_fd_sc_hd__nor2_2 _26301_ (.A(_04534_),
    .B(_04535_),
    .Y(_02079_));
 sky130_fd_sc_hd__and3_2 _26302_ (.A(_18122_),
    .B(_04532_),
    .C(\irq_pending[5] ),
    .X(_04536_));
 sky130_fd_sc_hd__a221o_2 _26303_ (.A1(_20347_),
    .A2(\reg_next_pc[5] ),
    .B1(_01476_),
    .B2(_04523_),
    .C1(_04536_),
    .X(_02080_));
 sky130_fd_sc_hd__nor2_2 _26304_ (.A(\reg_pc[6] ),
    .B(_04534_),
    .Y(_04537_));
 sky130_fd_sc_hd__nand2_2 _26305_ (.A(_04534_),
    .B(\reg_pc[6] ),
    .Y(_04538_));
 sky130_fd_sc_hd__inv_2 _26306_ (.A(_04538_),
    .Y(_04539_));
 sky130_fd_sc_hd__nor2_2 _26307_ (.A(_04537_),
    .B(_04539_),
    .Y(_02081_));
 sky130_fd_sc_hd__buf_1 _26308_ (.A(_04517_),
    .X(_04540_));
 sky130_fd_sc_hd__and3_2 _26309_ (.A(_18120_),
    .B(_04532_),
    .C(\irq_pending[6] ),
    .X(_04541_));
 sky130_fd_sc_hd__a221o_2 _26310_ (.A1(_20347_),
    .A2(\reg_next_pc[6] ),
    .B1(_01479_),
    .B2(_04540_),
    .C1(_04541_),
    .X(_02082_));
 sky130_fd_sc_hd__nor2_2 _26311_ (.A(_20172_),
    .B(_04538_),
    .Y(_04542_));
 sky130_fd_sc_hd__nor2_2 _26312_ (.A(\reg_pc[7] ),
    .B(_04539_),
    .Y(_04543_));
 sky130_fd_sc_hd__nor2_2 _26313_ (.A(_04542_),
    .B(_04543_),
    .Y(_02083_));
 sky130_fd_sc_hd__buf_1 _26314_ (.A(_18243_),
    .X(_04544_));
 sky130_fd_sc_hd__and3_2 _26315_ (.A(_18118_),
    .B(_04532_),
    .C(\irq_pending[7] ),
    .X(_04545_));
 sky130_fd_sc_hd__a221o_2 _26316_ (.A1(_04544_),
    .A2(\reg_next_pc[7] ),
    .B1(_01482_),
    .B2(_04540_),
    .C1(_04545_),
    .X(_02084_));
 sky130_fd_sc_hd__or2_2 _26317_ (.A(\reg_pc[8] ),
    .B(_04542_),
    .X(_04546_));
 sky130_fd_sc_hd__nand2_2 _26318_ (.A(_04542_),
    .B(\reg_pc[8] ),
    .Y(_04547_));
 sky130_fd_sc_hd__and2_2 _26319_ (.A(_04546_),
    .B(_04547_),
    .X(_02085_));
 sky130_fd_sc_hd__and3_2 _26320_ (.A(_18115_),
    .B(_04532_),
    .C(\irq_pending[8] ),
    .X(_04548_));
 sky130_fd_sc_hd__a221o_2 _26321_ (.A1(_04544_),
    .A2(\reg_next_pc[8] ),
    .B1(_01485_),
    .B2(_04540_),
    .C1(_04548_),
    .X(_02086_));
 sky130_fd_sc_hd__nor2_2 _26322_ (.A(_20185_),
    .B(_04547_),
    .Y(_04549_));
 sky130_fd_sc_hd__and2_2 _26323_ (.A(_04547_),
    .B(_20185_),
    .X(_04550_));
 sky130_fd_sc_hd__nor2_2 _26324_ (.A(_04549_),
    .B(_04550_),
    .Y(_02087_));
 sky130_fd_sc_hd__and3_2 _26325_ (.A(_18114_),
    .B(_04532_),
    .C(\irq_pending[9] ),
    .X(_04551_));
 sky130_fd_sc_hd__a221o_2 _26326_ (.A1(_04544_),
    .A2(\reg_next_pc[9] ),
    .B1(_01488_),
    .B2(_04540_),
    .C1(_04551_),
    .X(_02088_));
 sky130_fd_sc_hd__nor2_2 _26327_ (.A(\reg_pc[10] ),
    .B(_04549_),
    .Y(_04552_));
 sky130_fd_sc_hd__nand2_2 _26328_ (.A(_04549_),
    .B(\reg_pc[10] ),
    .Y(_04553_));
 sky130_fd_sc_hd__inv_2 _26329_ (.A(_04553_),
    .Y(_04554_));
 sky130_fd_sc_hd__nor2_2 _26330_ (.A(_04552_),
    .B(_04554_),
    .Y(_02089_));
 sky130_fd_sc_hd__and2_2 _26331_ (.A(_04521_),
    .B(\reg_next_pc[10] ),
    .X(_04555_));
 sky130_fd_sc_hd__a221o_2 _26332_ (.A1(_18113_),
    .A2(_04519_),
    .B1(_04518_),
    .B2(_01491_),
    .C1(_04555_),
    .X(_02090_));
 sky130_fd_sc_hd__nor2_2 _26333_ (.A(_18552_),
    .B(_04553_),
    .Y(_04556_));
 sky130_fd_sc_hd__nor2_2 _26334_ (.A(\reg_pc[11] ),
    .B(_04554_),
    .Y(_04557_));
 sky130_fd_sc_hd__nor2_2 _26335_ (.A(_04556_),
    .B(_04557_),
    .Y(_02091_));
 sky130_fd_sc_hd__and2_2 _26336_ (.A(_04521_),
    .B(\reg_next_pc[11] ),
    .X(_04558_));
 sky130_fd_sc_hd__a221o_2 _26337_ (.A1(_18112_),
    .A2(_04519_),
    .B1(_04518_),
    .B2(_01494_),
    .C1(_04558_),
    .X(_02092_));
 sky130_fd_sc_hd__nor2_2 _26338_ (.A(\reg_pc[12] ),
    .B(_04556_),
    .Y(_04559_));
 sky130_fd_sc_hd__nand2_2 _26339_ (.A(_04556_),
    .B(\reg_pc[12] ),
    .Y(_04560_));
 sky130_fd_sc_hd__inv_2 _26340_ (.A(_04560_),
    .Y(_04561_));
 sky130_fd_sc_hd__nor2_2 _26341_ (.A(_04559_),
    .B(_04561_),
    .Y(_02093_));
 sky130_fd_sc_hd__buf_1 _26342_ (.A(\irq_state[1] ),
    .X(_04562_));
 sky130_fd_sc_hd__and3_2 _26343_ (.A(_18135_),
    .B(_04562_),
    .C(\irq_pending[12] ),
    .X(_04563_));
 sky130_fd_sc_hd__a221o_2 _26344_ (.A1(_04544_),
    .A2(\reg_next_pc[12] ),
    .B1(_01497_),
    .B2(_04540_),
    .C1(_04563_),
    .X(_02094_));
 sky130_fd_sc_hd__nor2_2 _26345_ (.A(_20215_),
    .B(_04560_),
    .Y(_04564_));
 sky130_fd_sc_hd__nor2_2 _26346_ (.A(\reg_pc[13] ),
    .B(_04561_),
    .Y(_04565_));
 sky130_fd_sc_hd__nor2_2 _26347_ (.A(_04564_),
    .B(_04565_),
    .Y(_02095_));
 sky130_fd_sc_hd__and3_2 _26348_ (.A(_18134_),
    .B(_04562_),
    .C(\irq_pending[13] ),
    .X(_04566_));
 sky130_fd_sc_hd__a221o_2 _26349_ (.A1(_04544_),
    .A2(\reg_next_pc[13] ),
    .B1(_01500_),
    .B2(_04540_),
    .C1(_04566_),
    .X(_02096_));
 sky130_fd_sc_hd__nor2_2 _26350_ (.A(\reg_pc[14] ),
    .B(_04564_),
    .Y(_04567_));
 sky130_fd_sc_hd__and2_2 _26351_ (.A(_04564_),
    .B(\reg_pc[14] ),
    .X(_04568_));
 sky130_fd_sc_hd__nor2_2 _26352_ (.A(_04567_),
    .B(_04568_),
    .Y(_02097_));
 sky130_fd_sc_hd__buf_1 _26353_ (.A(_04516_),
    .X(_04569_));
 sky130_fd_sc_hd__and3_2 _26354_ (.A(_18139_),
    .B(_04562_),
    .C(\irq_pending[14] ),
    .X(_04570_));
 sky130_fd_sc_hd__a221o_2 _26355_ (.A1(_04544_),
    .A2(\reg_next_pc[14] ),
    .B1(_01503_),
    .B2(_04569_),
    .C1(_04570_),
    .X(_02098_));
 sky130_fd_sc_hd__nor2_2 _26356_ (.A(\reg_pc[15] ),
    .B(_04568_),
    .Y(_04571_));
 sky130_fd_sc_hd__nand2_2 _26357_ (.A(_04568_),
    .B(\reg_pc[15] ),
    .Y(_04572_));
 sky130_fd_sc_hd__inv_2 _26358_ (.A(_04572_),
    .Y(_04573_));
 sky130_fd_sc_hd__nor2_2 _26359_ (.A(_04571_),
    .B(_04573_),
    .Y(_02099_));
 sky130_fd_sc_hd__buf_1 _26360_ (.A(_04521_),
    .X(_04574_));
 sky130_fd_sc_hd__and3_2 _26361_ (.A(_18137_),
    .B(_04562_),
    .C(\irq_pending[15] ),
    .X(_04575_));
 sky130_fd_sc_hd__a221o_2 _26362_ (.A1(_04574_),
    .A2(\reg_next_pc[15] ),
    .B1(_01506_),
    .B2(_04569_),
    .C1(_04575_),
    .X(_02100_));
 sky130_fd_sc_hd__nor2_2 _26363_ (.A(_20235_),
    .B(_04572_),
    .Y(_04576_));
 sky130_fd_sc_hd__nor2_2 _26364_ (.A(\reg_pc[16] ),
    .B(_04573_),
    .Y(_04577_));
 sky130_fd_sc_hd__nor2_2 _26365_ (.A(_04576_),
    .B(_04577_),
    .Y(_02101_));
 sky130_fd_sc_hd__and2_2 _26366_ (.A(_04521_),
    .B(\reg_next_pc[16] ),
    .X(_04578_));
 sky130_fd_sc_hd__a221o_2 _26367_ (.A1(_18091_),
    .A2(_04519_),
    .B1(_04518_),
    .B2(_01509_),
    .C1(_04578_),
    .X(_02102_));
 sky130_fd_sc_hd__nor2_2 _26368_ (.A(\reg_pc[17] ),
    .B(_04576_),
    .Y(_04579_));
 sky130_fd_sc_hd__and2_2 _26369_ (.A(_04576_),
    .B(\reg_pc[17] ),
    .X(_04580_));
 sky130_fd_sc_hd__nor2_2 _26370_ (.A(_04579_),
    .B(_04580_),
    .Y(_02103_));
 sky130_fd_sc_hd__and3_2 _26371_ (.A(_18089_),
    .B(_04562_),
    .C(\irq_pending[17] ),
    .X(_04581_));
 sky130_fd_sc_hd__a221o_2 _26372_ (.A1(_04574_),
    .A2(\reg_next_pc[17] ),
    .B1(_01512_),
    .B2(_04569_),
    .C1(_04581_),
    .X(_02104_));
 sky130_fd_sc_hd__or2_2 _26373_ (.A(\reg_pc[18] ),
    .B(_04580_),
    .X(_04582_));
 sky130_fd_sc_hd__nand2_2 _26374_ (.A(_04580_),
    .B(\reg_pc[18] ),
    .Y(_04583_));
 sky130_fd_sc_hd__and2_2 _26375_ (.A(_04582_),
    .B(_04583_),
    .X(_02105_));
 sky130_fd_sc_hd__and3_2 _26376_ (.A(_18094_),
    .B(_04562_),
    .C(\irq_pending[18] ),
    .X(_04584_));
 sky130_fd_sc_hd__a221o_2 _26377_ (.A1(_04574_),
    .A2(\reg_next_pc[18] ),
    .B1(_01515_),
    .B2(_04569_),
    .C1(_04584_),
    .X(_02106_));
 sky130_fd_sc_hd__nor2_2 _26378_ (.A(_20257_),
    .B(_04583_),
    .Y(_04585_));
 sky130_fd_sc_hd__and2_2 _26379_ (.A(_04583_),
    .B(_20257_),
    .X(_04586_));
 sky130_fd_sc_hd__nor2_2 _26380_ (.A(_04585_),
    .B(_04586_),
    .Y(_02107_));
 sky130_fd_sc_hd__buf_1 _26381_ (.A(\irq_state[1] ),
    .X(_04587_));
 sky130_fd_sc_hd__and3_2 _26382_ (.A(_18092_),
    .B(_04587_),
    .C(\irq_pending[19] ),
    .X(_04588_));
 sky130_fd_sc_hd__a221o_2 _26383_ (.A1(_04574_),
    .A2(\reg_next_pc[19] ),
    .B1(_01518_),
    .B2(_04569_),
    .C1(_04588_),
    .X(_02108_));
 sky130_fd_sc_hd__nor2_2 _26384_ (.A(\reg_pc[20] ),
    .B(_04585_),
    .Y(_04589_));
 sky130_fd_sc_hd__nand2_2 _26385_ (.A(_04585_),
    .B(\reg_pc[20] ),
    .Y(_04590_));
 sky130_fd_sc_hd__inv_2 _26386_ (.A(_04590_),
    .Y(_04591_));
 sky130_fd_sc_hd__nor2_2 _26387_ (.A(_04589_),
    .B(_04591_),
    .Y(_02109_));
 sky130_fd_sc_hd__and3_2 _26388_ (.A(_18108_),
    .B(_04587_),
    .C(\irq_pending[20] ),
    .X(_04592_));
 sky130_fd_sc_hd__a221o_2 _26389_ (.A1(_04574_),
    .A2(\reg_next_pc[20] ),
    .B1(_01521_),
    .B2(_04569_),
    .C1(_04592_),
    .X(_02110_));
 sky130_fd_sc_hd__nor2_2 _26390_ (.A(_20272_),
    .B(_04590_),
    .Y(_04593_));
 sky130_fd_sc_hd__nor2_2 _26391_ (.A(\reg_pc[21] ),
    .B(_04591_),
    .Y(_04594_));
 sky130_fd_sc_hd__nor2_2 _26392_ (.A(_04593_),
    .B(_04594_),
    .Y(_02111_));
 sky130_fd_sc_hd__buf_1 _26393_ (.A(_04516_),
    .X(_04595_));
 sky130_fd_sc_hd__and3_2 _26394_ (.A(_18107_),
    .B(_04587_),
    .C(\irq_pending[21] ),
    .X(_04596_));
 sky130_fd_sc_hd__a221o_2 _26395_ (.A1(_04574_),
    .A2(\reg_next_pc[21] ),
    .B1(_01524_),
    .B2(_04595_),
    .C1(_04596_),
    .X(_02112_));
 sky130_fd_sc_hd__or2_2 _26396_ (.A(\reg_pc[22] ),
    .B(_04593_),
    .X(_04597_));
 sky130_fd_sc_hd__nand2_2 _26397_ (.A(_04593_),
    .B(\reg_pc[22] ),
    .Y(_04598_));
 sky130_fd_sc_hd__and2_2 _26398_ (.A(_04597_),
    .B(_04598_),
    .X(_02113_));
 sky130_fd_sc_hd__buf_1 _26399_ (.A(_04521_),
    .X(_04599_));
 sky130_fd_sc_hd__and3_2 _26400_ (.A(_18105_),
    .B(_04587_),
    .C(\irq_pending[22] ),
    .X(_04600_));
 sky130_fd_sc_hd__a221o_2 _26401_ (.A1(_04599_),
    .A2(\reg_next_pc[22] ),
    .B1(_01527_),
    .B2(_04595_),
    .C1(_04600_),
    .X(_02114_));
 sky130_fd_sc_hd__nor2_2 _26402_ (.A(_20286_),
    .B(_04598_),
    .Y(_04601_));
 sky130_fd_sc_hd__and2_2 _26403_ (.A(_04598_),
    .B(_20286_),
    .X(_04602_));
 sky130_fd_sc_hd__nor2_2 _26404_ (.A(_04601_),
    .B(_04602_),
    .Y(_02115_));
 sky130_fd_sc_hd__and3_2 _26405_ (.A(_18103_),
    .B(_04587_),
    .C(\irq_pending[23] ),
    .X(_04603_));
 sky130_fd_sc_hd__a221o_2 _26406_ (.A1(_04599_),
    .A2(\reg_next_pc[23] ),
    .B1(_01530_),
    .B2(_04595_),
    .C1(_04603_),
    .X(_02116_));
 sky130_fd_sc_hd__nor2_2 _26407_ (.A(\reg_pc[24] ),
    .B(_04601_),
    .Y(_04604_));
 sky130_fd_sc_hd__nand2_2 _26408_ (.A(_04601_),
    .B(\reg_pc[24] ),
    .Y(_04605_));
 sky130_fd_sc_hd__inv_2 _26409_ (.A(_04605_),
    .Y(_04606_));
 sky130_fd_sc_hd__nor2_2 _26410_ (.A(_04604_),
    .B(_04606_),
    .Y(_02117_));
 sky130_fd_sc_hd__and3_2 _26411_ (.A(_18100_),
    .B(_04587_),
    .C(\irq_pending[24] ),
    .X(_04607_));
 sky130_fd_sc_hd__a221o_2 _26412_ (.A1(_04599_),
    .A2(\reg_next_pc[24] ),
    .B1(_01533_),
    .B2(_04595_),
    .C1(_04607_),
    .X(_02118_));
 sky130_fd_sc_hd__nor2_2 _26413_ (.A(_20297_),
    .B(_04605_),
    .Y(_04608_));
 sky130_fd_sc_hd__nor2_2 _26414_ (.A(\reg_pc[25] ),
    .B(_04606_),
    .Y(_04609_));
 sky130_fd_sc_hd__nor2_2 _26415_ (.A(_04608_),
    .B(_04609_),
    .Y(_02119_));
 sky130_fd_sc_hd__and3_2 _26416_ (.A(_18099_),
    .B(_04531_),
    .C(\irq_pending[25] ),
    .X(_04610_));
 sky130_fd_sc_hd__a221o_2 _26417_ (.A1(_04599_),
    .A2(\reg_next_pc[25] ),
    .B1(_01536_),
    .B2(_04595_),
    .C1(_04610_),
    .X(_02120_));
 sky130_fd_sc_hd__nor2_2 _26418_ (.A(\reg_pc[26] ),
    .B(_04608_),
    .Y(_04611_));
 sky130_fd_sc_hd__nand2_2 _26419_ (.A(_04608_),
    .B(\reg_pc[26] ),
    .Y(_04612_));
 sky130_fd_sc_hd__inv_2 _26420_ (.A(_04612_),
    .Y(_04613_));
 sky130_fd_sc_hd__nor2_2 _26421_ (.A(_04611_),
    .B(_04613_),
    .Y(_02121_));
 sky130_fd_sc_hd__and2_2 _26422_ (.A(_18240_),
    .B(\reg_next_pc[26] ),
    .X(_04614_));
 sky130_fd_sc_hd__a221o_2 _26423_ (.A1(_18098_),
    .A2(_04519_),
    .B1(_04523_),
    .B2(_01539_),
    .C1(_04614_),
    .X(_02122_));
 sky130_fd_sc_hd__nor2_2 _26424_ (.A(_20312_),
    .B(_04612_),
    .Y(_04615_));
 sky130_fd_sc_hd__nor2_2 _26425_ (.A(\reg_pc[27] ),
    .B(_04613_),
    .Y(_04616_));
 sky130_fd_sc_hd__nor2_2 _26426_ (.A(_04615_),
    .B(_04616_),
    .Y(_02123_));
 sky130_fd_sc_hd__and2_2 _26427_ (.A(_18240_),
    .B(\reg_next_pc[27] ),
    .X(_04617_));
 sky130_fd_sc_hd__a221o_2 _26428_ (.A1(_18097_),
    .A2(_18236_),
    .B1(_04523_),
    .B2(_01542_),
    .C1(_04617_),
    .X(_02124_));
 sky130_fd_sc_hd__nor2_2 _26429_ (.A(\reg_pc[28] ),
    .B(_04615_),
    .Y(_04618_));
 sky130_fd_sc_hd__nand2_2 _26430_ (.A(_04615_),
    .B(\reg_pc[28] ),
    .Y(_04619_));
 sky130_fd_sc_hd__inv_2 _26431_ (.A(_04619_),
    .Y(_04620_));
 sky130_fd_sc_hd__nor2_2 _26432_ (.A(_04618_),
    .B(_04620_),
    .Y(_02125_));
 sky130_fd_sc_hd__and3_2 _26433_ (.A(_18127_),
    .B(_04531_),
    .C(\irq_pending[28] ),
    .X(_04621_));
 sky130_fd_sc_hd__a221o_2 _26434_ (.A1(_04599_),
    .A2(\reg_next_pc[28] ),
    .B1(_01545_),
    .B2(_04595_),
    .C1(_04621_),
    .X(_02126_));
 sky130_fd_sc_hd__nor2_2 _26435_ (.A(_20327_),
    .B(_04619_),
    .Y(_04622_));
 sky130_fd_sc_hd__nor2_2 _26436_ (.A(\reg_pc[29] ),
    .B(_04620_),
    .Y(_04623_));
 sky130_fd_sc_hd__nor2_2 _26437_ (.A(_04622_),
    .B(_04623_),
    .Y(_02127_));
 sky130_fd_sc_hd__and3_2 _26438_ (.A(_18126_),
    .B(_04531_),
    .C(\irq_pending[29] ),
    .X(_04624_));
 sky130_fd_sc_hd__a221o_2 _26439_ (.A1(_04599_),
    .A2(\reg_next_pc[29] ),
    .B1(_01548_),
    .B2(_04517_),
    .C1(_04624_),
    .X(_02128_));
 sky130_fd_sc_hd__nor2_2 _26440_ (.A(\reg_pc[30] ),
    .B(_04622_),
    .Y(_04625_));
 sky130_fd_sc_hd__and2_2 _26441_ (.A(_04622_),
    .B(\reg_pc[30] ),
    .X(_04626_));
 sky130_fd_sc_hd__nor2_2 _26442_ (.A(_04625_),
    .B(_04626_),
    .Y(_02129_));
 sky130_fd_sc_hd__and3_2 _26443_ (.A(_18131_),
    .B(_04531_),
    .C(\irq_pending[30] ),
    .X(_04627_));
 sky130_fd_sc_hd__a221o_2 _26444_ (.A1(_18243_),
    .A2(\reg_next_pc[30] ),
    .B1(_01551_),
    .B2(_04517_),
    .C1(_04627_),
    .X(_02130_));
 sky130_fd_sc_hd__xor2_2 _26445_ (.A(\reg_pc[31] ),
    .B(_04626_),
    .X(_02131_));
 sky130_fd_sc_hd__and3_2 _26446_ (.A(_18129_),
    .B(_04531_),
    .C(\irq_pending[31] ),
    .X(_04628_));
 sky130_fd_sc_hd__a221o_2 _26447_ (.A1(_18243_),
    .A2(\reg_next_pc[31] ),
    .B1(_01554_),
    .B2(_04517_),
    .C1(_04628_),
    .X(_02132_));
 sky130_fd_sc_hd__nor2_2 _26448_ (.A(instr_or),
    .B(instr_ori),
    .Y(_04629_));
 sky130_fd_sc_hd__inv_2 _26449_ (.A(_04629_),
    .Y(_04630_));
 sky130_fd_sc_hd__buf_1 _26450_ (.A(_04630_),
    .X(_04631_));
 sky130_fd_sc_hd__or3_2 _26451_ (.A(is_compare),
    .B(_04631_),
    .C(_18220_),
    .X(_04632_));
 sky130_fd_sc_hd__nor2_2 _26452_ (.A(instr_and),
    .B(instr_andi),
    .Y(_04633_));
 sky130_fd_sc_hd__nor2_2 _26453_ (.A(instr_sll),
    .B(instr_slli),
    .Y(_04634_));
 sky130_fd_sc_hd__nor2_2 _26454_ (.A(instr_xor),
    .B(instr_xori),
    .Y(_04635_));
 sky130_fd_sc_hd__buf_1 _26455_ (.A(_04635_),
    .X(_04636_));
 sky130_fd_sc_hd__and4b_2 _26456_ (.A_N(_04632_),
    .B(_04633_),
    .C(_04634_),
    .D(_04636_),
    .X(_02133_));
 sky130_fd_sc_hd__buf_1 _26457_ (.A(_04629_),
    .X(_04637_));
 sky130_fd_sc_hd__o21ai_2 _26458_ (.A1(_19790_),
    .A2(_04633_),
    .B1(_04637_),
    .Y(_04638_));
 sky130_fd_sc_hd__inv_2 _26459_ (.A(_00343_),
    .Y(_04639_));
 sky130_fd_sc_hd__buf_1 _26460_ (.A(_04630_),
    .X(_04640_));
 sky130_fd_sc_hd__a22o_2 _26461_ (.A1(_04639_),
    .A2(is_compare),
    .B1(_04640_),
    .B2(_19535_),
    .X(_04641_));
 sky130_fd_sc_hd__inv_2 _26462_ (.A(_04634_),
    .Y(_04642_));
 sky130_fd_sc_hd__buf_1 _26463_ (.A(_04642_),
    .X(_04643_));
 sky130_fd_sc_hd__and2_2 _26464_ (.A(_04643_),
    .B(\alu_shl[0] ),
    .X(_04644_));
 sky130_fd_sc_hd__buf_1 _26465_ (.A(_18220_),
    .X(_04645_));
 sky130_fd_sc_hd__inv_2 _26466_ (.A(_04635_),
    .Y(_04646_));
 sky130_fd_sc_hd__buf_1 _26467_ (.A(_04646_),
    .X(_04647_));
 sky130_fd_sc_hd__a22o_2 _26468_ (.A1(_04645_),
    .A2(\alu_shr[0] ),
    .B1(_02591_),
    .B2(_04647_),
    .X(_04648_));
 sky130_fd_sc_hd__a2111o_2 _26469_ (.A1(_19156_),
    .A2(_04638_),
    .B1(_04641_),
    .C1(_04644_),
    .D1(_04648_),
    .X(_02134_));
 sky130_fd_sc_hd__buf_1 _26470_ (.A(_04643_),
    .X(_04649_));
 sky130_fd_sc_hd__buf_1 _26471_ (.A(_04649_),
    .X(_04650_));
 sky130_fd_sc_hd__inv_2 _26472_ (.A(_04633_),
    .Y(_04651_));
 sky130_fd_sc_hd__nor2_2 _26473_ (.A(_04630_),
    .B(_04651_),
    .Y(_04652_));
 sky130_fd_sc_hd__inv_2 _26474_ (.A(_04652_),
    .Y(_04653_));
 sky130_fd_sc_hd__o211a_2 _26475_ (.A1(_04640_),
    .A2(_19868_),
    .B1(_19869_),
    .C1(_04653_),
    .X(_04654_));
 sky130_fd_sc_hd__buf_1 _26476_ (.A(_18220_),
    .X(_04655_));
 sky130_fd_sc_hd__nor2_2 _26477_ (.A(_04636_),
    .B(_19870_),
    .Y(_04656_));
 sky130_fd_sc_hd__a21o_2 _26478_ (.A1(\alu_shr[1] ),
    .A2(_04655_),
    .B1(_04656_),
    .X(_04657_));
 sky130_fd_sc_hd__a211o_2 _26479_ (.A1(\alu_shl[1] ),
    .A2(_04650_),
    .B1(_04654_),
    .C1(_04657_),
    .X(_02135_));
 sky130_fd_sc_hd__buf_1 _26480_ (.A(_04645_),
    .X(_04658_));
 sky130_fd_sc_hd__buf_1 _26481_ (.A(_04646_),
    .X(_04659_));
 sky130_fd_sc_hd__buf_1 _26482_ (.A(_04659_),
    .X(_04660_));
 sky130_fd_sc_hd__nor2_2 _26483_ (.A(_19914_),
    .B(_04629_),
    .Y(_04661_));
 sky130_fd_sc_hd__and2_2 _26484_ (.A(_19916_),
    .B(_04651_),
    .X(_04662_));
 sky130_fd_sc_hd__a211o_2 _26485_ (.A1(\alu_shl[2] ),
    .A2(_04649_),
    .B1(_04661_),
    .C1(_04662_),
    .X(_04663_));
 sky130_fd_sc_hd__a221o_2 _26486_ (.A1(\alu_shr[2] ),
    .A2(_04658_),
    .B1(_19917_),
    .B2(_04660_),
    .C1(_04663_),
    .X(_02136_));
 sky130_fd_sc_hd__buf_1 _26487_ (.A(_04651_),
    .X(_04664_));
 sky130_fd_sc_hd__buf_1 _26488_ (.A(_04664_),
    .X(_04665_));
 sky130_fd_sc_hd__buf_1 _26489_ (.A(_04629_),
    .X(_04666_));
 sky130_fd_sc_hd__nor2_2 _26490_ (.A(_19910_),
    .B(_04666_),
    .Y(_04667_));
 sky130_fd_sc_hd__a21o_2 _26491_ (.A1(_19912_),
    .A2(_04665_),
    .B1(_04667_),
    .X(_04668_));
 sky130_fd_sc_hd__a22o_2 _26492_ (.A1(_19913_),
    .A2(_04660_),
    .B1(_04655_),
    .B2(\alu_shr[3] ),
    .X(_04669_));
 sky130_fd_sc_hd__a211o_2 _26493_ (.A1(\alu_shl[3] ),
    .A2(_04650_),
    .B1(_04668_),
    .C1(_04669_),
    .X(_02137_));
 sky130_fd_sc_hd__buf_1 _26494_ (.A(_04659_),
    .X(_04670_));
 sky130_fd_sc_hd__buf_1 _26495_ (.A(_04645_),
    .X(_04671_));
 sky130_fd_sc_hd__buf_1 _26496_ (.A(_04643_),
    .X(_04672_));
 sky130_fd_sc_hd__nand2_2 _26497_ (.A(_04672_),
    .B(\alu_shl[4] ),
    .Y(_04673_));
 sky130_fd_sc_hd__nand2_2 _26498_ (.A(_19908_),
    .B(_04665_),
    .Y(_04674_));
 sky130_fd_sc_hd__o211ai_2 _26499_ (.A1(_19906_),
    .A2(_04637_),
    .B1(_04673_),
    .C1(_04674_),
    .Y(_04675_));
 sky130_fd_sc_hd__a221o_2 _26500_ (.A1(_19909_),
    .A2(_04670_),
    .B1(_04671_),
    .B2(\alu_shr[4] ),
    .C1(_04675_),
    .X(_02138_));
 sky130_fd_sc_hd__nor2_2 _26501_ (.A(_19920_),
    .B(_04633_),
    .Y(_04676_));
 sky130_fd_sc_hd__a21o_2 _26502_ (.A1(_04640_),
    .A2(_19919_),
    .B1(_04676_),
    .X(_04677_));
 sky130_fd_sc_hd__a22o_2 _26503_ (.A1(_19922_),
    .A2(_04647_),
    .B1(_04655_),
    .B2(\alu_shr[5] ),
    .X(_04678_));
 sky130_fd_sc_hd__a211o_2 _26504_ (.A1(\alu_shl[5] ),
    .A2(_04650_),
    .B1(_04677_),
    .C1(_04678_),
    .X(_02139_));
 sky130_fd_sc_hd__nand2_2 _26505_ (.A(_04672_),
    .B(\alu_shl[6] ),
    .Y(_04679_));
 sky130_fd_sc_hd__nand2_2 _26506_ (.A(_19859_),
    .B(_04665_),
    .Y(_04680_));
 sky130_fd_sc_hd__o211ai_2 _26507_ (.A1(_19857_),
    .A2(_04637_),
    .B1(_04679_),
    .C1(_04680_),
    .Y(_04681_));
 sky130_fd_sc_hd__a221o_2 _26508_ (.A1(_19860_),
    .A2(_04670_),
    .B1(_04671_),
    .B2(\alu_shr[6] ),
    .C1(_04681_),
    .X(_02140_));
 sky130_fd_sc_hd__o211a_2 _26509_ (.A1(_04640_),
    .A2(_19863_),
    .B1(_19864_),
    .C1(_04653_),
    .X(_04682_));
 sky130_fd_sc_hd__nor2_2 _26510_ (.A(_04636_),
    .B(_19865_),
    .Y(_04683_));
 sky130_fd_sc_hd__a21o_2 _26511_ (.A1(\alu_shr[7] ),
    .A2(_04655_),
    .B1(_04683_),
    .X(_04684_));
 sky130_fd_sc_hd__a211o_2 _26512_ (.A1(\alu_shl[7] ),
    .A2(_04650_),
    .B1(_04682_),
    .C1(_04684_),
    .X(_02141_));
 sky130_fd_sc_hd__nand2_2 _26513_ (.A(_04672_),
    .B(\alu_shl[8] ),
    .Y(_04685_));
 sky130_fd_sc_hd__nand2_2 _26514_ (.A(_19899_),
    .B(_04665_),
    .Y(_04686_));
 sky130_fd_sc_hd__o211ai_2 _26515_ (.A1(_19897_),
    .A2(_04637_),
    .B1(_04685_),
    .C1(_04686_),
    .Y(_04687_));
 sky130_fd_sc_hd__a221o_2 _26516_ (.A1(_19900_),
    .A2(_04670_),
    .B1(_04671_),
    .B2(\alu_shr[8] ),
    .C1(_04687_),
    .X(_02142_));
 sky130_fd_sc_hd__nand2_2 _26517_ (.A(_04672_),
    .B(\alu_shl[9] ),
    .Y(_04688_));
 sky130_fd_sc_hd__nand2_2 _26518_ (.A(_19895_),
    .B(_04665_),
    .Y(_04689_));
 sky130_fd_sc_hd__o211ai_2 _26519_ (.A1(_19893_),
    .A2(_04637_),
    .B1(_04688_),
    .C1(_04689_),
    .Y(_04690_));
 sky130_fd_sc_hd__a221o_2 _26520_ (.A1(_19896_),
    .A2(_04670_),
    .B1(_04671_),
    .B2(\alu_shr[9] ),
    .C1(_04690_),
    .X(_02143_));
 sky130_fd_sc_hd__buf_1 _26521_ (.A(_04645_),
    .X(_04691_));
 sky130_fd_sc_hd__buf_1 _26522_ (.A(_04652_),
    .X(_04692_));
 sky130_fd_sc_hd__buf_1 _26523_ (.A(_04692_),
    .X(_04693_));
 sky130_fd_sc_hd__nor2_2 _26524_ (.A(_19901_),
    .B(_04693_),
    .Y(_04694_));
 sky130_fd_sc_hd__or2_2 _26525_ (.A(_19903_),
    .B(_04631_),
    .X(_04695_));
 sky130_fd_sc_hd__buf_1 _26526_ (.A(_04642_),
    .X(_04696_));
 sky130_fd_sc_hd__a22o_2 _26527_ (.A1(\alu_shl[10] ),
    .A2(_04696_),
    .B1(_19904_),
    .B2(_04647_),
    .X(_04697_));
 sky130_fd_sc_hd__a221o_2 _26528_ (.A1(\alu_shr[10] ),
    .A2(_04691_),
    .B1(_04694_),
    .B2(_04695_),
    .C1(_04697_),
    .X(_02144_));
 sky130_fd_sc_hd__nor2_2 _26529_ (.A(_19889_),
    .B(_04629_),
    .Y(_04698_));
 sky130_fd_sc_hd__and2_2 _26530_ (.A(_19891_),
    .B(_04651_),
    .X(_04699_));
 sky130_fd_sc_hd__a211o_2 _26531_ (.A1(\alu_shl[11] ),
    .A2(_04649_),
    .B1(_04698_),
    .C1(_04699_),
    .X(_04700_));
 sky130_fd_sc_hd__a221o_2 _26532_ (.A1(\alu_shr[11] ),
    .A2(_04691_),
    .B1(_19892_),
    .B2(_04660_),
    .C1(_04700_),
    .X(_02145_));
 sky130_fd_sc_hd__nand2_2 _26533_ (.A(_04672_),
    .B(\alu_shl[12] ),
    .Y(_04701_));
 sky130_fd_sc_hd__nand2_2 _26534_ (.A(_19882_),
    .B(_04664_),
    .Y(_04702_));
 sky130_fd_sc_hd__o211ai_2 _26535_ (.A1(_19880_),
    .A2(_04666_),
    .B1(_04701_),
    .C1(_04702_),
    .Y(_04703_));
 sky130_fd_sc_hd__a221o_2 _26536_ (.A1(_19883_),
    .A2(_04670_),
    .B1(_04658_),
    .B2(\alu_shr[12] ),
    .C1(_04703_),
    .X(_02146_));
 sky130_fd_sc_hd__nor2_2 _26537_ (.A(_19876_),
    .B(_04693_),
    .Y(_04704_));
 sky130_fd_sc_hd__or2_2 _26538_ (.A(_19878_),
    .B(_04631_),
    .X(_04705_));
 sky130_fd_sc_hd__a22o_2 _26539_ (.A1(\alu_shl[13] ),
    .A2(_04696_),
    .B1(_19879_),
    .B2(_04647_),
    .X(_04706_));
 sky130_fd_sc_hd__a221o_2 _26540_ (.A1(\alu_shr[13] ),
    .A2(_04691_),
    .B1(_04704_),
    .B2(_04705_),
    .C1(_04706_),
    .X(_02147_));
 sky130_fd_sc_hd__nor2_2 _26541_ (.A(_19884_),
    .B(_04693_),
    .Y(_04707_));
 sky130_fd_sc_hd__or2_2 _26542_ (.A(_19886_),
    .B(_04631_),
    .X(_04708_));
 sky130_fd_sc_hd__buf_1 _26543_ (.A(_04659_),
    .X(_04709_));
 sky130_fd_sc_hd__a22o_2 _26544_ (.A1(\alu_shl[14] ),
    .A2(_04696_),
    .B1(_19887_),
    .B2(_04709_),
    .X(_04710_));
 sky130_fd_sc_hd__a221o_2 _26545_ (.A1(\alu_shr[14] ),
    .A2(_04691_),
    .B1(_04707_),
    .B2(_04708_),
    .C1(_04710_),
    .X(_02148_));
 sky130_fd_sc_hd__nor2_2 _26546_ (.A(_19872_),
    .B(_04629_),
    .Y(_04711_));
 sky130_fd_sc_hd__and2_2 _26547_ (.A(_19874_),
    .B(_04651_),
    .X(_04712_));
 sky130_fd_sc_hd__a211o_2 _26548_ (.A1(\alu_shl[15] ),
    .A2(_04672_),
    .B1(_04711_),
    .C1(_04712_),
    .X(_04713_));
 sky130_fd_sc_hd__a221o_2 _26549_ (.A1(\alu_shr[15] ),
    .A2(_04691_),
    .B1(_19875_),
    .B2(_04660_),
    .C1(_04713_),
    .X(_02149_));
 sky130_fd_sc_hd__inv_2 _26550_ (.A(pcpi_rs2[16]),
    .Y(_02363_));
 sky130_fd_sc_hd__a21oi_2 _26551_ (.A1(_02363_),
    .A2(_20237_),
    .B1(_04637_),
    .Y(_04714_));
 sky130_fd_sc_hd__nor2_2 _26552_ (.A(_04636_),
    .B(_19997_),
    .Y(_04715_));
 sky130_fd_sc_hd__a32o_2 _26553_ (.A1(_04664_),
    .A2(pcpi_rs2[16]),
    .A3(_19519_),
    .B1(\alu_shl[16] ),
    .B2(_04649_),
    .X(_04716_));
 sky130_fd_sc_hd__a2111o_2 _26554_ (.A1(_04658_),
    .A2(\alu_shr[16] ),
    .B1(_04714_),
    .C1(_04715_),
    .D1(_04716_),
    .X(_02150_));
 sky130_fd_sc_hd__nand2_2 _26555_ (.A(_04696_),
    .B(\alu_shl[17] ),
    .Y(_04717_));
 sky130_fd_sc_hd__nand2_2 _26556_ (.A(_19984_),
    .B(_04664_),
    .Y(_04718_));
 sky130_fd_sc_hd__o211ai_2 _26557_ (.A1(_19982_),
    .A2(_04666_),
    .B1(_04717_),
    .C1(_04718_),
    .Y(_04719_));
 sky130_fd_sc_hd__a221o_2 _26558_ (.A1(_19985_),
    .A2(_04670_),
    .B1(_04658_),
    .B2(\alu_shr[17] ),
    .C1(_04719_),
    .X(_02151_));
 sky130_fd_sc_hd__nor2_2 _26559_ (.A(_19992_),
    .B(_04693_),
    .Y(_04720_));
 sky130_fd_sc_hd__or2_2 _26560_ (.A(_19994_),
    .B(_04631_),
    .X(_04721_));
 sky130_fd_sc_hd__buf_1 _26561_ (.A(_04643_),
    .X(_04722_));
 sky130_fd_sc_hd__a22o_2 _26562_ (.A1(\alu_shl[18] ),
    .A2(_04722_),
    .B1(_19995_),
    .B2(_04709_),
    .X(_04723_));
 sky130_fd_sc_hd__a221o_2 _26563_ (.A1(\alu_shr[18] ),
    .A2(_04691_),
    .B1(_04720_),
    .B2(_04721_),
    .C1(_04723_),
    .X(_02152_));
 sky130_fd_sc_hd__nand2_2 _26564_ (.A(_04696_),
    .B(\alu_shl[19] ),
    .Y(_04724_));
 sky130_fd_sc_hd__nand2_2 _26565_ (.A(_19989_),
    .B(_04664_),
    .Y(_04725_));
 sky130_fd_sc_hd__o211ai_2 _26566_ (.A1(_19987_),
    .A2(_04666_),
    .B1(_04724_),
    .C1(_04725_),
    .Y(_04726_));
 sky130_fd_sc_hd__a221o_2 _26567_ (.A1(_19990_),
    .A2(_04660_),
    .B1(_04658_),
    .B2(\alu_shr[19] ),
    .C1(_04726_),
    .X(_02153_));
 sky130_fd_sc_hd__o211a_2 _26568_ (.A1(_04640_),
    .A2(_19940_),
    .B1(_19941_),
    .C1(_04653_),
    .X(_04727_));
 sky130_fd_sc_hd__nor2_2 _26569_ (.A(_04636_),
    .B(_19942_),
    .Y(_04728_));
 sky130_fd_sc_hd__a21o_2 _26570_ (.A1(\alu_shl[20] ),
    .A2(_04649_),
    .B1(_04728_),
    .X(_04729_));
 sky130_fd_sc_hd__a211o_2 _26571_ (.A1(\alu_shr[20] ),
    .A2(_04671_),
    .B1(_04727_),
    .C1(_04729_),
    .X(_02154_));
 sky130_fd_sc_hd__buf_1 _26572_ (.A(_04645_),
    .X(_04730_));
 sky130_fd_sc_hd__nor2_2 _26573_ (.A(_19925_),
    .B(_04693_),
    .Y(_04731_));
 sky130_fd_sc_hd__buf_1 _26574_ (.A(_04630_),
    .X(_04732_));
 sky130_fd_sc_hd__or2_2 _26575_ (.A(_19927_),
    .B(_04732_),
    .X(_04733_));
 sky130_fd_sc_hd__a22o_2 _26576_ (.A1(\alu_shl[21] ),
    .A2(_04722_),
    .B1(_19928_),
    .B2(_04709_),
    .X(_04734_));
 sky130_fd_sc_hd__a221o_2 _26577_ (.A1(\alu_shr[21] ),
    .A2(_04730_),
    .B1(_04731_),
    .B2(_04733_),
    .C1(_04734_),
    .X(_02155_));
 sky130_fd_sc_hd__nor2_2 _26578_ (.A(_19934_),
    .B(_04693_),
    .Y(_04735_));
 sky130_fd_sc_hd__or2_2 _26579_ (.A(_19936_),
    .B(_04732_),
    .X(_04736_));
 sky130_fd_sc_hd__a22o_2 _26580_ (.A1(\alu_shl[22] ),
    .A2(_04722_),
    .B1(_19937_),
    .B2(_04709_),
    .X(_04737_));
 sky130_fd_sc_hd__a221o_2 _26581_ (.A1(\alu_shr[22] ),
    .A2(_04730_),
    .B1(_04735_),
    .B2(_04736_),
    .C1(_04737_),
    .X(_02156_));
 sky130_fd_sc_hd__nor2_2 _26582_ (.A(_19929_),
    .B(_04692_),
    .Y(_04738_));
 sky130_fd_sc_hd__or2_2 _26583_ (.A(_19931_),
    .B(_04732_),
    .X(_04739_));
 sky130_fd_sc_hd__a22o_2 _26584_ (.A1(\alu_shl[23] ),
    .A2(_04722_),
    .B1(_19932_),
    .B2(_04709_),
    .X(_04740_));
 sky130_fd_sc_hd__a221o_2 _26585_ (.A1(\alu_shr[23] ),
    .A2(_04730_),
    .B1(_04738_),
    .B2(_04739_),
    .C1(_04740_),
    .X(_02157_));
 sky130_fd_sc_hd__o211a_2 _26586_ (.A1(_04631_),
    .A2(_19958_),
    .B1(_19959_),
    .C1(_04653_),
    .X(_04741_));
 sky130_fd_sc_hd__nor2_2 _26587_ (.A(_04636_),
    .B(_19960_),
    .Y(_04742_));
 sky130_fd_sc_hd__a21o_2 _26588_ (.A1(\alu_shl[24] ),
    .A2(_04649_),
    .B1(_04742_),
    .X(_04743_));
 sky130_fd_sc_hd__a211o_2 _26589_ (.A1(\alu_shr[24] ),
    .A2(_04671_),
    .B1(_04741_),
    .C1(_04743_),
    .X(_02158_));
 sky130_fd_sc_hd__nor2_2 _26590_ (.A(_19944_),
    .B(_04692_),
    .Y(_04744_));
 sky130_fd_sc_hd__or2_2 _26591_ (.A(_19946_),
    .B(_04732_),
    .X(_04745_));
 sky130_fd_sc_hd__a22o_2 _26592_ (.A1(\alu_shl[25] ),
    .A2(_04722_),
    .B1(_19947_),
    .B2(_04709_),
    .X(_04746_));
 sky130_fd_sc_hd__a221o_2 _26593_ (.A1(\alu_shr[25] ),
    .A2(_04730_),
    .B1(_04744_),
    .B2(_04745_),
    .C1(_04746_),
    .X(_02159_));
 sky130_fd_sc_hd__nor2_2 _26594_ (.A(_19954_),
    .B(_04633_),
    .Y(_04747_));
 sky130_fd_sc_hd__a21o_2 _26595_ (.A1(_04640_),
    .A2(_19953_),
    .B1(_04747_),
    .X(_04748_));
 sky130_fd_sc_hd__a22o_2 _26596_ (.A1(_19956_),
    .A2(_04647_),
    .B1(_04655_),
    .B2(\alu_shr[26] ),
    .X(_04749_));
 sky130_fd_sc_hd__a211o_2 _26597_ (.A1(\alu_shl[26] ),
    .A2(_04650_),
    .B1(_04748_),
    .C1(_04749_),
    .X(_02160_));
 sky130_fd_sc_hd__nor2_2 _26598_ (.A(_19966_),
    .B(_04692_),
    .Y(_04750_));
 sky130_fd_sc_hd__or2_2 _26599_ (.A(_19968_),
    .B(_04732_),
    .X(_04751_));
 sky130_fd_sc_hd__a22o_2 _26600_ (.A1(\alu_shl[27] ),
    .A2(_04722_),
    .B1(_19969_),
    .B2(_04659_),
    .X(_04752_));
 sky130_fd_sc_hd__a221o_2 _26601_ (.A1(\alu_shr[27] ),
    .A2(_04730_),
    .B1(_04750_),
    .B2(_04751_),
    .C1(_04752_),
    .X(_02161_));
 sky130_fd_sc_hd__nor2_2 _26602_ (.A(_19948_),
    .B(_04692_),
    .Y(_04753_));
 sky130_fd_sc_hd__or2_2 _26603_ (.A(_19950_),
    .B(_04732_),
    .X(_04754_));
 sky130_fd_sc_hd__a22o_2 _26604_ (.A1(\alu_shl[28] ),
    .A2(_04643_),
    .B1(_19951_),
    .B2(_04659_),
    .X(_04755_));
 sky130_fd_sc_hd__a221o_2 _26605_ (.A1(\alu_shr[28] ),
    .A2(_04730_),
    .B1(_04753_),
    .B2(_04754_),
    .C1(_04755_),
    .X(_02162_));
 sky130_fd_sc_hd__nor2_2 _26606_ (.A(_19962_),
    .B(_04692_),
    .Y(_04756_));
 sky130_fd_sc_hd__or2_2 _26607_ (.A(_19964_),
    .B(_04630_),
    .X(_04757_));
 sky130_fd_sc_hd__a22o_2 _26608_ (.A1(\alu_shl[29] ),
    .A2(_04643_),
    .B1(_19965_),
    .B2(_04659_),
    .X(_04758_));
 sky130_fd_sc_hd__a221o_2 _26609_ (.A1(\alu_shr[29] ),
    .A2(_04655_),
    .B1(_04756_),
    .B2(_04757_),
    .C1(_04758_),
    .X(_02163_));
 sky130_fd_sc_hd__nand2_2 _26610_ (.A(_04696_),
    .B(\alu_shl[30] ),
    .Y(_04759_));
 sky130_fd_sc_hd__nand2_2 _26611_ (.A(_19976_),
    .B(_04664_),
    .Y(_04760_));
 sky130_fd_sc_hd__o211ai_2 _26612_ (.A1(_19974_),
    .A2(_04666_),
    .B1(_04759_),
    .C1(_04760_),
    .Y(_04761_));
 sky130_fd_sc_hd__a221o_2 _26613_ (.A1(_19977_),
    .A2(_04660_),
    .B1(_04658_),
    .B2(\alu_shr[30] ),
    .C1(_04761_),
    .X(_02164_));
 sky130_fd_sc_hd__nor2_2 _26614_ (.A(_19970_),
    .B(_04666_),
    .Y(_04762_));
 sky130_fd_sc_hd__a21o_2 _26615_ (.A1(_19972_),
    .A2(_04665_),
    .B1(_04762_),
    .X(_04763_));
 sky130_fd_sc_hd__a22o_2 _26616_ (.A1(_19973_),
    .A2(_04647_),
    .B1(_04645_),
    .B2(\alu_shr[31] ),
    .X(_04764_));
 sky130_fd_sc_hd__a211o_2 _26617_ (.A1(\alu_shl[31] ),
    .A2(_04650_),
    .B1(_04763_),
    .C1(_04764_),
    .X(_02165_));
 sky130_fd_sc_hd__and3_2 _26618_ (.A(_00289_),
    .B(_18012_),
    .C(_20016_),
    .X(_02166_));
 sky130_fd_sc_hd__buf_1 _26619_ (.A(\mem_wordsize[1] ),
    .X(_04765_));
 sky130_fd_sc_hd__a22o_2 _26620_ (.A1(pcpi_rs2[8]),
    .A2(_04156_),
    .B1(_19156_),
    .B2(_04765_),
    .X(_02167_));
 sky130_fd_sc_hd__buf_1 _26621_ (.A(_04086_),
    .X(_04766_));
 sky130_fd_sc_hd__a22o_2 _26622_ (.A1(_19147_),
    .A2(_04766_),
    .B1(_19155_),
    .B2(_04765_),
    .X(_02168_));
 sky130_fd_sc_hd__a22o_2 _26623_ (.A1(pcpi_rs2[10]),
    .A2(_04766_),
    .B1(_19154_),
    .B2(_04765_),
    .X(_02169_));
 sky130_fd_sc_hd__a22o_2 _26624_ (.A1(_19146_),
    .A2(_04766_),
    .B1(_19778_),
    .B2(_04765_),
    .X(_02170_));
 sky130_fd_sc_hd__a22o_2 _26625_ (.A1(pcpi_rs2[12]),
    .A2(_04766_),
    .B1(_19152_),
    .B2(_04765_),
    .X(_02171_));
 sky130_fd_sc_hd__a22o_2 _26626_ (.A1(_19145_),
    .A2(_04766_),
    .B1(_19151_),
    .B2(\mem_wordsize[1] ),
    .X(_02172_));
 sky130_fd_sc_hd__a22o_2 _26627_ (.A1(_19143_),
    .A2(_04766_),
    .B1(_19150_),
    .B2(\mem_wordsize[1] ),
    .X(_02173_));
 sky130_fd_sc_hd__a22o_2 _26628_ (.A1(_19142_),
    .A2(_04086_),
    .B1(_19149_),
    .B2(\mem_wordsize[1] ),
    .X(_02174_));
 sky130_fd_sc_hd__o21a_2 _26629_ (.A1(_04156_),
    .A2(_04765_),
    .B1(_19156_),
    .X(_02175_));
 sky130_fd_sc_hd__nor2_2 _26630_ (.A(_02318_),
    .B(_04457_),
    .Y(_02176_));
 sky130_fd_sc_hd__buf_1 _26631_ (.A(_04085_),
    .X(_04767_));
 sky130_fd_sc_hd__nor2_2 _26632_ (.A(_02321_),
    .B(_04767_),
    .Y(_02177_));
 sky130_fd_sc_hd__nor2_2 _26633_ (.A(_02324_),
    .B(_04767_),
    .Y(_02178_));
 sky130_fd_sc_hd__nor2_2 _26634_ (.A(_02327_),
    .B(_04767_),
    .Y(_02179_));
 sky130_fd_sc_hd__nor2_2 _26635_ (.A(_02330_),
    .B(_04767_),
    .Y(_02180_));
 sky130_fd_sc_hd__nor2_2 _26636_ (.A(_02333_),
    .B(_04767_),
    .Y(_02181_));
 sky130_fd_sc_hd__nor2_2 _26637_ (.A(_02336_),
    .B(_04767_),
    .Y(_02182_));
 sky130_fd_sc_hd__nand2_2 _26638_ (.A(_20020_),
    .B(latched_store),
    .Y(_02183_));
 sky130_fd_sc_hd__or2_2 _26639_ (.A(\irq_pending[3] ),
    .B(irq[3]),
    .X(_02214_));
 sky130_fd_sc_hd__and2_2 _26640_ (.A(_02214_),
    .B(\irq_mask[3] ),
    .X(_02215_));
 sky130_fd_sc_hd__inv_2 _26641_ (.A(_01700_),
    .Y(_02217_));
 sky130_fd_sc_hd__or2_2 _26642_ (.A(\irq_pending[4] ),
    .B(irq[4]),
    .X(_02218_));
 sky130_fd_sc_hd__and2_2 _26643_ (.A(_02218_),
    .B(\irq_mask[4] ),
    .X(_02219_));
 sky130_fd_sc_hd__or2_2 _26644_ (.A(\irq_pending[5] ),
    .B(irq[5]),
    .X(_02221_));
 sky130_fd_sc_hd__and2_2 _26645_ (.A(_02221_),
    .B(\irq_mask[5] ),
    .X(_02222_));
 sky130_fd_sc_hd__or2_2 _26646_ (.A(\irq_pending[6] ),
    .B(irq[6]),
    .X(_02224_));
 sky130_fd_sc_hd__and2_2 _26647_ (.A(_02224_),
    .B(\irq_mask[6] ),
    .X(_02225_));
 sky130_fd_sc_hd__or2_2 _26648_ (.A(\irq_pending[7] ),
    .B(irq[7]),
    .X(_02227_));
 sky130_fd_sc_hd__and2_2 _26649_ (.A(_02227_),
    .B(\irq_mask[7] ),
    .X(_02228_));
 sky130_fd_sc_hd__or2_2 _26650_ (.A(\irq_pending[8] ),
    .B(irq[8]),
    .X(_02230_));
 sky130_fd_sc_hd__and2_2 _26651_ (.A(_02230_),
    .B(\irq_mask[8] ),
    .X(_02231_));
 sky130_fd_sc_hd__or2_2 _26652_ (.A(\irq_pending[9] ),
    .B(irq[9]),
    .X(_02233_));
 sky130_fd_sc_hd__and2_2 _26653_ (.A(_02233_),
    .B(\irq_mask[9] ),
    .X(_02234_));
 sky130_fd_sc_hd__or2_2 _26654_ (.A(\irq_pending[10] ),
    .B(irq[10]),
    .X(_02236_));
 sky130_fd_sc_hd__and2_2 _26655_ (.A(_02236_),
    .B(\irq_mask[10] ),
    .X(_02237_));
 sky130_fd_sc_hd__or2_2 _26656_ (.A(\irq_pending[11] ),
    .B(irq[11]),
    .X(_02239_));
 sky130_fd_sc_hd__and2_2 _26657_ (.A(_02239_),
    .B(\irq_mask[11] ),
    .X(_02240_));
 sky130_fd_sc_hd__or2_2 _26658_ (.A(\irq_pending[12] ),
    .B(irq[12]),
    .X(_02242_));
 sky130_fd_sc_hd__and2_2 _26659_ (.A(_02242_),
    .B(\irq_mask[12] ),
    .X(_02243_));
 sky130_fd_sc_hd__or2_2 _26660_ (.A(\irq_pending[13] ),
    .B(irq[13]),
    .X(_02245_));
 sky130_fd_sc_hd__and2_2 _26661_ (.A(_02245_),
    .B(\irq_mask[13] ),
    .X(_02246_));
 sky130_fd_sc_hd__or2_2 _26662_ (.A(\irq_pending[14] ),
    .B(irq[14]),
    .X(_02248_));
 sky130_fd_sc_hd__and2_2 _26663_ (.A(_02248_),
    .B(\irq_mask[14] ),
    .X(_02249_));
 sky130_fd_sc_hd__or2_2 _26664_ (.A(\irq_pending[15] ),
    .B(irq[15]),
    .X(_02251_));
 sky130_fd_sc_hd__and2_2 _26665_ (.A(_02251_),
    .B(\irq_mask[15] ),
    .X(_02252_));
 sky130_fd_sc_hd__or2_2 _26666_ (.A(\irq_pending[16] ),
    .B(irq[16]),
    .X(_02254_));
 sky130_fd_sc_hd__and2_2 _26667_ (.A(_02254_),
    .B(\irq_mask[16] ),
    .X(_02255_));
 sky130_fd_sc_hd__or2_2 _26668_ (.A(\irq_pending[17] ),
    .B(irq[17]),
    .X(_02257_));
 sky130_fd_sc_hd__and2_2 _26669_ (.A(_02257_),
    .B(\irq_mask[17] ),
    .X(_02258_));
 sky130_fd_sc_hd__or2_2 _26670_ (.A(\irq_pending[18] ),
    .B(irq[18]),
    .X(_02260_));
 sky130_fd_sc_hd__and2_2 _26671_ (.A(_02260_),
    .B(\irq_mask[18] ),
    .X(_02261_));
 sky130_fd_sc_hd__or2_2 _26672_ (.A(\irq_pending[19] ),
    .B(irq[19]),
    .X(_02263_));
 sky130_fd_sc_hd__and2_2 _26673_ (.A(_02263_),
    .B(\irq_mask[19] ),
    .X(_02264_));
 sky130_fd_sc_hd__or2_2 _26674_ (.A(\irq_pending[20] ),
    .B(irq[20]),
    .X(_02266_));
 sky130_fd_sc_hd__and2_2 _26675_ (.A(_02266_),
    .B(\irq_mask[20] ),
    .X(_02267_));
 sky130_fd_sc_hd__or2_2 _26676_ (.A(\irq_pending[21] ),
    .B(irq[21]),
    .X(_02269_));
 sky130_fd_sc_hd__and2_2 _26677_ (.A(_02269_),
    .B(\irq_mask[21] ),
    .X(_02270_));
 sky130_fd_sc_hd__or2_2 _26678_ (.A(\irq_pending[22] ),
    .B(irq[22]),
    .X(_02272_));
 sky130_fd_sc_hd__and2_2 _26679_ (.A(_02272_),
    .B(\irq_mask[22] ),
    .X(_02273_));
 sky130_fd_sc_hd__or2_2 _26680_ (.A(\irq_pending[23] ),
    .B(irq[23]),
    .X(_02275_));
 sky130_fd_sc_hd__and2_2 _26681_ (.A(_02275_),
    .B(\irq_mask[23] ),
    .X(_02276_));
 sky130_fd_sc_hd__or2_2 _26682_ (.A(\irq_pending[24] ),
    .B(irq[24]),
    .X(_02278_));
 sky130_fd_sc_hd__and2_2 _26683_ (.A(_02278_),
    .B(\irq_mask[24] ),
    .X(_02279_));
 sky130_fd_sc_hd__or2_2 _26684_ (.A(\irq_pending[25] ),
    .B(irq[25]),
    .X(_02281_));
 sky130_fd_sc_hd__and2_2 _26685_ (.A(_02281_),
    .B(\irq_mask[25] ),
    .X(_02282_));
 sky130_fd_sc_hd__or2_2 _26686_ (.A(\irq_pending[26] ),
    .B(irq[26]),
    .X(_02284_));
 sky130_fd_sc_hd__and2_2 _26687_ (.A(_02284_),
    .B(\irq_mask[26] ),
    .X(_02285_));
 sky130_fd_sc_hd__or2_2 _26688_ (.A(\irq_pending[27] ),
    .B(irq[27]),
    .X(_02287_));
 sky130_fd_sc_hd__and2_2 _26689_ (.A(_02287_),
    .B(\irq_mask[27] ),
    .X(_02288_));
 sky130_fd_sc_hd__or2_2 _26690_ (.A(\irq_pending[28] ),
    .B(irq[28]),
    .X(_02290_));
 sky130_fd_sc_hd__and2_2 _26691_ (.A(_02290_),
    .B(\irq_mask[28] ),
    .X(_02291_));
 sky130_fd_sc_hd__or2_2 _26692_ (.A(\irq_pending[29] ),
    .B(irq[29]),
    .X(_02293_));
 sky130_fd_sc_hd__and2_2 _26693_ (.A(_02293_),
    .B(\irq_mask[29] ),
    .X(_02294_));
 sky130_fd_sc_hd__or2_2 _26694_ (.A(\irq_pending[30] ),
    .B(irq[30]),
    .X(_02296_));
 sky130_fd_sc_hd__and2_2 _26695_ (.A(_02296_),
    .B(\irq_mask[30] ),
    .X(_02297_));
 sky130_fd_sc_hd__or2_2 _26696_ (.A(\irq_pending[31] ),
    .B(irq[31]),
    .X(_02299_));
 sky130_fd_sc_hd__and2_2 _26697_ (.A(_02299_),
    .B(\irq_mask[31] ),
    .X(_02300_));
 sky130_fd_sc_hd__nor2_2 _26698_ (.A(\timer[27] ),
    .B(\timer[26] ),
    .Y(_04768_));
 sky130_fd_sc_hd__and3b_2 _26699_ (.A_N(_20021_),
    .B(_20052_),
    .C(_04768_),
    .X(_04769_));
 sky130_fd_sc_hd__or2_2 _26700_ (.A(\timer[11] ),
    .B(\timer[10] ),
    .X(_04770_));
 sky130_fd_sc_hd__or2_2 _26701_ (.A(\timer[13] ),
    .B(\timer[12] ),
    .X(_04771_));
 sky130_fd_sc_hd__or4_2 _26702_ (.A(\timer[3] ),
    .B(\timer[2] ),
    .C(\timer[7] ),
    .D(\timer[6] ),
    .X(_04772_));
 sky130_fd_sc_hd__nor3_2 _26703_ (.A(_04770_),
    .B(_04771_),
    .C(_04772_),
    .Y(_04773_));
 sky130_fd_sc_hd__and4_2 _26704_ (.A(_20045_),
    .B(_04506_),
    .C(_04494_),
    .D(_20048_),
    .X(_04774_));
 sky130_fd_sc_hd__nor2_2 _26705_ (.A(\timer[15] ),
    .B(\timer[14] ),
    .Y(_04775_));
 sky130_fd_sc_hd__and3_2 _26706_ (.A(_04775_),
    .B(_04119_),
    .C(\timer[0] ),
    .X(_04776_));
 sky130_fd_sc_hd__and3_2 _26707_ (.A(_04776_),
    .B(_20022_),
    .C(_20033_),
    .X(_04777_));
 sky130_fd_sc_hd__a41o_2 _26708_ (.A1(_04769_),
    .A2(_04773_),
    .A3(_04774_),
    .A4(_04777_),
    .B1(\irq_pending[0] ),
    .X(_02302_));
 sky130_fd_sc_hd__or2_2 _26709_ (.A(_02303_),
    .B(irq[0]),
    .X(_02304_));
 sky130_fd_sc_hd__and2_2 _26710_ (.A(_02304_),
    .B(\irq_mask[0] ),
    .X(_02305_));
 sky130_fd_sc_hd__nor2_2 _26711_ (.A(\irq_pending[2] ),
    .B(irq[2]),
    .Y(_02307_));
 sky130_fd_sc_hd__or2_2 _26712_ (.A(_18081_),
    .B(_02307_),
    .X(_02308_));
 sky130_fd_sc_hd__nor2_2 _26713_ (.A(_02310_),
    .B(_18278_),
    .Y(_02311_));
 sky130_fd_sc_hd__or2_2 _26714_ (.A(_19805_),
    .B(_02311_),
    .X(_02312_));
 sky130_fd_sc_hd__or2_2 _26715_ (.A(_02313_),
    .B(_19805_),
    .X(_02314_));
 sky130_fd_sc_hd__or2_2 _26716_ (.A(_02316_),
    .B(_19805_),
    .X(_02317_));
 sky130_fd_sc_hd__nor2_2 _26717_ (.A(pcpi_rs1[31]),
    .B(_19971_),
    .Y(_04778_));
 sky130_fd_sc_hd__or2_2 _26718_ (.A(_19787_),
    .B(_00048_),
    .X(_04779_));
 sky130_fd_sc_hd__inv_2 _26719_ (.A(_19788_),
    .Y(_04780_));
 sky130_fd_sc_hd__nor2_2 _26720_ (.A(_19789_),
    .B(_04780_),
    .Y(_00049_));
 sky130_fd_sc_hd__a2111o_2 _26721_ (.A1(_04779_),
    .A2(_19533_),
    .B1(_00049_),
    .C1(_19913_),
    .D1(_19917_),
    .X(_04781_));
 sky130_fd_sc_hd__nand2_2 _26722_ (.A(_19911_),
    .B(_19153_),
    .Y(_04782_));
 sky130_fd_sc_hd__nand2_2 _26723_ (.A(_19915_),
    .B(mem_la_wdata[2]),
    .Y(_04783_));
 sky130_fd_sc_hd__or2_2 _26724_ (.A(_04783_),
    .B(_19913_),
    .X(_04784_));
 sky130_fd_sc_hd__a311o_2 _26725_ (.A1(_04781_),
    .A2(_04782_),
    .A3(_04784_),
    .B1(_19922_),
    .C1(_19909_),
    .X(_04785_));
 sky130_fd_sc_hd__nand2_2 _26726_ (.A(_19918_),
    .B(_19151_),
    .Y(_04786_));
 sky130_fd_sc_hd__or3_2 _26727_ (.A(_19777_),
    .B(_19530_),
    .C(_19922_),
    .X(_04787_));
 sky130_fd_sc_hd__a31o_2 _26728_ (.A1(_04785_),
    .A2(_04786_),
    .A3(_04787_),
    .B1(_19860_),
    .X(_04788_));
 sky130_fd_sc_hd__nand2_2 _26729_ (.A(_19858_),
    .B(_19150_),
    .Y(_04789_));
 sky130_fd_sc_hd__a21bo_2 _26730_ (.A1(_04788_),
    .A2(_04789_),
    .B1_N(_19865_),
    .X(_04790_));
 sky130_fd_sc_hd__nand2_2 _26731_ (.A(_19862_),
    .B(_19149_),
    .Y(_04791_));
 sky130_fd_sc_hd__a21o_2 _26732_ (.A1(_04790_),
    .A2(_04791_),
    .B1(_19905_),
    .X(_04792_));
 sky130_fd_sc_hd__nand2_2 _26733_ (.A(_19890_),
    .B(_19146_),
    .Y(_04793_));
 sky130_fd_sc_hd__or3_2 _26734_ (.A(_02339_),
    .B(_19526_),
    .C(_19896_),
    .X(_04794_));
 sky130_fd_sc_hd__nand2_2 _26735_ (.A(_19894_),
    .B(_19147_),
    .Y(_04795_));
 sky130_fd_sc_hd__a21o_2 _26736_ (.A1(_04794_),
    .A2(_04795_),
    .B1(_19904_),
    .X(_04796_));
 sky130_fd_sc_hd__nand2_2 _26737_ (.A(_19902_),
    .B(pcpi_rs2[10]),
    .Y(_04797_));
 sky130_fd_sc_hd__a21o_2 _26738_ (.A1(_04796_),
    .A2(_04797_),
    .B1(_19892_),
    .X(_04798_));
 sky130_fd_sc_hd__a31o_2 _26739_ (.A1(_04792_),
    .A2(_04793_),
    .A3(_04798_),
    .B1(_19888_),
    .X(_04799_));
 sky130_fd_sc_hd__nand2_2 _26740_ (.A(_19873_),
    .B(_19142_),
    .Y(_04800_));
 sky130_fd_sc_hd__or3_2 _26741_ (.A(_02351_),
    .B(_19523_),
    .C(_19879_),
    .X(_04801_));
 sky130_fd_sc_hd__nand2_2 _26742_ (.A(_19877_),
    .B(_19145_),
    .Y(_04802_));
 sky130_fd_sc_hd__a21o_2 _26743_ (.A1(_04801_),
    .A2(_04802_),
    .B1(_19887_),
    .X(_04803_));
 sky130_fd_sc_hd__nand2_2 _26744_ (.A(_19885_),
    .B(_19143_),
    .Y(_04804_));
 sky130_fd_sc_hd__a21o_2 _26745_ (.A1(_04803_),
    .A2(_04804_),
    .B1(_19875_),
    .X(_04805_));
 sky130_fd_sc_hd__nand2_2 _26746_ (.A(_19998_),
    .B(_19943_),
    .Y(_04806_));
 sky130_fd_sc_hd__a31o_2 _26747_ (.A1(_04799_),
    .A2(_04800_),
    .A3(_04805_),
    .B1(_04806_),
    .X(_04807_));
 sky130_fd_sc_hd__nor2_2 _26748_ (.A(_19518_),
    .B(_02366_),
    .Y(_04808_));
 sky130_fd_sc_hd__and3_2 _26749_ (.A(_19986_),
    .B(pcpi_rs2[16]),
    .C(_20237_),
    .X(_04809_));
 sky130_fd_sc_hd__o21ai_2 _26750_ (.A1(_04808_),
    .A2(_04809_),
    .B1(_19996_),
    .Y(_04810_));
 sky130_fd_sc_hd__nand2_2 _26751_ (.A(_19993_),
    .B(_19141_),
    .Y(_04811_));
 sky130_fd_sc_hd__a21o_2 _26752_ (.A1(_04810_),
    .A2(_04811_),
    .B1(_19990_),
    .X(_04812_));
 sky130_fd_sc_hd__o21ai_2 _26753_ (.A1(_02372_),
    .A2(_19515_),
    .B1(_04812_),
    .Y(_04813_));
 sky130_fd_sc_hd__nor2_2 _26754_ (.A(_02375_),
    .B(_19928_),
    .Y(_04814_));
 sky130_fd_sc_hd__a22o_2 _26755_ (.A1(_19139_),
    .A2(_19926_),
    .B1(_04814_),
    .B2(_19939_),
    .X(_04815_));
 sky130_fd_sc_hd__nor2_2 _26756_ (.A(_19513_),
    .B(_02381_),
    .Y(_04816_));
 sky130_fd_sc_hd__a21oi_2 _26757_ (.A1(_04815_),
    .A2(_19938_),
    .B1(_04816_),
    .Y(_04817_));
 sky130_fd_sc_hd__nor2_2 _26758_ (.A(_19932_),
    .B(_04817_),
    .Y(_04818_));
 sky130_fd_sc_hd__a221oi_2 _26759_ (.A1(_19138_),
    .A2(_19930_),
    .B1(_04813_),
    .B2(_19943_),
    .C1(_04818_),
    .Y(_04819_));
 sky130_fd_sc_hd__a21bo_2 _26760_ (.A1(_04807_),
    .A2(_04819_),
    .B1_N(_19981_),
    .X(_04820_));
 sky130_fd_sc_hd__or3_2 _26761_ (.A(_02387_),
    .B(_19511_),
    .C(_19947_),
    .X(_04821_));
 sky130_fd_sc_hd__nand2_2 _26762_ (.A(_19945_),
    .B(_19137_),
    .Y(_04822_));
 sky130_fd_sc_hd__a21o_2 _26763_ (.A1(_04821_),
    .A2(_04822_),
    .B1(_19956_),
    .X(_04823_));
 sky130_fd_sc_hd__nand2_2 _26764_ (.A(_19952_),
    .B(pcpi_rs2[26]),
    .Y(_04824_));
 sky130_fd_sc_hd__a21o_2 _26765_ (.A1(_04823_),
    .A2(_04824_),
    .B1(_19969_),
    .X(_04825_));
 sky130_fd_sc_hd__nand2_2 _26766_ (.A(_19967_),
    .B(_19135_),
    .Y(_04826_));
 sky130_fd_sc_hd__a211o_2 _26767_ (.A1(_04825_),
    .A2(_04826_),
    .B1(_19951_),
    .C1(_19965_),
    .X(_04827_));
 sky130_fd_sc_hd__nand2_2 _26768_ (.A(_19963_),
    .B(_19134_),
    .Y(_04828_));
 sky130_fd_sc_hd__or3_2 _26769_ (.A(_02399_),
    .B(_19507_),
    .C(_19965_),
    .X(_04829_));
 sky130_fd_sc_hd__a31o_2 _26770_ (.A1(_04827_),
    .A2(_04828_),
    .A3(_04829_),
    .B1(_19979_),
    .X(_04830_));
 sky130_fd_sc_hd__o31a_2 _26771_ (.A1(_02405_),
    .A2(_19505_),
    .A3(_19973_),
    .B1(_04830_),
    .X(_04831_));
 sky130_fd_sc_hd__nand2_2 _26772_ (.A(_04820_),
    .B(_04831_),
    .Y(_04832_));
 sky130_fd_sc_hd__o21ba_2 _26773_ (.A1(_04778_),
    .A2(_04832_),
    .B1_N(_00000_),
    .X(_00002_));
 sky130_fd_sc_hd__nor2_2 _26774_ (.A(_04778_),
    .B(_00000_),
    .Y(_04833_));
 sky130_fd_sc_hd__o21a_2 _26775_ (.A1(_19973_),
    .A2(_04832_),
    .B1(_04833_),
    .X(_00001_));
 sky130_fd_sc_hd__buf_1 _26776_ (.A(\pcpi_mul.rs2[0] ),
    .X(_04834_));
 sky130_fd_sc_hd__inv_2 _26777_ (.A(_04834_),
    .Y(_04835_));
 sky130_fd_sc_hd__buf_1 _26778_ (.A(_04835_),
    .X(_04836_));
 sky130_fd_sc_hd__inv_2 _26779_ (.A(\pcpi_mul.rs1[0] ),
    .Y(_04837_));
 sky130_fd_sc_hd__buf_1 _26780_ (.A(_04837_),
    .X(_04838_));
 sky130_fd_sc_hd__buf_1 _26781_ (.A(_04838_),
    .X(_04839_));
 sky130_fd_sc_hd__buf_1 _26782_ (.A(_04839_),
    .X(_04840_));
 sky130_fd_sc_hd__nor2_2 _26783_ (.A(_04836_),
    .B(_04840_),
    .Y(_02623_));
 sky130_fd_sc_hd__nand2_2 _26784_ (.A(_19155_),
    .B(mem_la_wdata[0]),
    .Y(_04841_));
 sky130_fd_sc_hd__nand2_2 _26785_ (.A(_04780_),
    .B(_04841_),
    .Y(_02319_));
 sky130_fd_sc_hd__nor2_2 _26786_ (.A(_19533_),
    .B(_02320_),
    .Y(_04842_));
 sky130_fd_sc_hd__nand2_2 _26787_ (.A(_19533_),
    .B(_02320_),
    .Y(_04843_));
 sky130_fd_sc_hd__or2b_2 _26788_ (.A(_04842_),
    .B_N(_04843_),
    .X(_04844_));
 sky130_fd_sc_hd__xor2_2 _26789_ (.A(_19855_),
    .B(_04844_),
    .X(_02602_));
 sky130_fd_sc_hd__nor2_2 _26790_ (.A(_19154_),
    .B(_04780_),
    .Y(_04845_));
 sky130_fd_sc_hd__inv_2 _26791_ (.A(_04845_),
    .Y(_04846_));
 sky130_fd_sc_hd__nand2_2 _26792_ (.A(_04780_),
    .B(_19154_),
    .Y(_04847_));
 sky130_fd_sc_hd__nand2_2 _26793_ (.A(_04846_),
    .B(_04847_),
    .Y(_02322_));
 sky130_fd_sc_hd__or2_2 _26794_ (.A(_19532_),
    .B(_02323_),
    .X(_04848_));
 sky130_fd_sc_hd__nand2_2 _26795_ (.A(_19532_),
    .B(_02323_),
    .Y(_04849_));
 sky130_fd_sc_hd__nand2_2 _26796_ (.A(_04848_),
    .B(_04849_),
    .Y(_04850_));
 sky130_fd_sc_hd__o21ai_2 _26797_ (.A1(_04842_),
    .A2(_19855_),
    .B1(_04843_),
    .Y(_04851_));
 sky130_fd_sc_hd__xnor2_2 _26798_ (.A(_04850_),
    .B(_04851_),
    .Y(_02613_));
 sky130_fd_sc_hd__nand2_2 _26799_ (.A(_04846_),
    .B(_19778_),
    .Y(_04852_));
 sky130_fd_sc_hd__nand2_2 _26800_ (.A(_04852_),
    .B(_19791_),
    .Y(_02325_));
 sky130_fd_sc_hd__nor2_2 _26801_ (.A(_19531_),
    .B(_02326_),
    .Y(_04853_));
 sky130_fd_sc_hd__nand2_2 _26802_ (.A(_19531_),
    .B(_02326_),
    .Y(_04854_));
 sky130_fd_sc_hd__inv_2 _26803_ (.A(_04854_),
    .Y(_04855_));
 sky130_fd_sc_hd__nor2_2 _26804_ (.A(_04853_),
    .B(_04855_),
    .Y(_04856_));
 sky130_fd_sc_hd__nand2_2 _26805_ (.A(_04851_),
    .B(_04848_),
    .Y(_04857_));
 sky130_fd_sc_hd__nand2_2 _26806_ (.A(_04857_),
    .B(_04849_),
    .Y(_04858_));
 sky130_fd_sc_hd__xor2_2 _26807_ (.A(_04856_),
    .B(_04858_),
    .X(_02616_));
 sky130_fd_sc_hd__nand2_2 _26808_ (.A(_19791_),
    .B(_19152_),
    .Y(_04859_));
 sky130_fd_sc_hd__nand2_2 _26809_ (.A(_19793_),
    .B(_04859_),
    .Y(_02328_));
 sky130_fd_sc_hd__inv_2 _26810_ (.A(_02329_),
    .Y(_04860_));
 sky130_fd_sc_hd__nor2_2 _26811_ (.A(_19907_),
    .B(_04860_),
    .Y(_04861_));
 sky130_fd_sc_hd__inv_2 _26812_ (.A(_04861_),
    .Y(_04862_));
 sky130_fd_sc_hd__nor2_2 _26813_ (.A(_19530_),
    .B(_02329_),
    .Y(_04863_));
 sky130_fd_sc_hd__inv_2 _26814_ (.A(_04863_),
    .Y(_04864_));
 sky130_fd_sc_hd__nand2_2 _26815_ (.A(_04862_),
    .B(_04864_),
    .Y(_04865_));
 sky130_fd_sc_hd__a21oi_2 _26816_ (.A1(_04857_),
    .A2(_04849_),
    .B1(_04853_),
    .Y(_04866_));
 sky130_fd_sc_hd__nor2_2 _26817_ (.A(_04855_),
    .B(_04866_),
    .Y(_04867_));
 sky130_fd_sc_hd__xor2_2 _26818_ (.A(_04865_),
    .B(_04867_),
    .X(_02617_));
 sky130_fd_sc_hd__nand2_2 _26819_ (.A(_19793_),
    .B(_19151_),
    .Y(_04868_));
 sky130_fd_sc_hd__nand2_2 _26820_ (.A(_19792_),
    .B(_02330_),
    .Y(_04869_));
 sky130_fd_sc_hd__nand2_2 _26821_ (.A(_04868_),
    .B(_04869_),
    .Y(_02331_));
 sky130_fd_sc_hd__nor2_2 _26822_ (.A(_19529_),
    .B(_02332_),
    .Y(_04870_));
 sky130_fd_sc_hd__nand2_2 _26823_ (.A(_19529_),
    .B(_02332_),
    .Y(_04871_));
 sky130_fd_sc_hd__inv_2 _26824_ (.A(_04871_),
    .Y(_04872_));
 sky130_fd_sc_hd__nor2_2 _26825_ (.A(_04870_),
    .B(_04872_),
    .Y(_04873_));
 sky130_fd_sc_hd__o21ai_2 _26826_ (.A1(_04855_),
    .A2(_04866_),
    .B1(_04864_),
    .Y(_04874_));
 sky130_fd_sc_hd__nand2_2 _26827_ (.A(_04874_),
    .B(_04862_),
    .Y(_04875_));
 sky130_fd_sc_hd__xor2_2 _26828_ (.A(_04873_),
    .B(_04875_),
    .X(_02618_));
 sky130_fd_sc_hd__or2_2 _26829_ (.A(mem_la_wdata[6]),
    .B(_04869_),
    .X(_04876_));
 sky130_fd_sc_hd__nand2_2 _26830_ (.A(_04869_),
    .B(_19150_),
    .Y(_04877_));
 sky130_fd_sc_hd__nand2_2 _26831_ (.A(_04876_),
    .B(_04877_),
    .Y(_02334_));
 sky130_fd_sc_hd__xor2_2 _26832_ (.A(pcpi_rs1[6]),
    .B(_02335_),
    .X(_04878_));
 sky130_fd_sc_hd__a21oi_2 _26833_ (.A1(_04874_),
    .A2(_04862_),
    .B1(_04870_),
    .Y(_04879_));
 sky130_fd_sc_hd__or2_2 _26834_ (.A(_04872_),
    .B(_04879_),
    .X(_04880_));
 sky130_fd_sc_hd__or2_2 _26835_ (.A(_04878_),
    .B(_04880_),
    .X(_04881_));
 sky130_fd_sc_hd__nand2_2 _26836_ (.A(_04880_),
    .B(_04878_),
    .Y(_04882_));
 sky130_fd_sc_hd__and2_2 _26837_ (.A(_04881_),
    .B(_04882_),
    .X(_02619_));
 sky130_fd_sc_hd__nor2_2 _26838_ (.A(mem_la_wdata[7]),
    .B(_04876_),
    .Y(_04883_));
 sky130_fd_sc_hd__and2_2 _26839_ (.A(_04876_),
    .B(_19149_),
    .X(_04884_));
 sky130_fd_sc_hd__or2_2 _26840_ (.A(_04883_),
    .B(_04884_),
    .X(_02337_));
 sky130_fd_sc_hd__nor2_2 _26841_ (.A(pcpi_rs1[7]),
    .B(_02338_),
    .Y(_04885_));
 sky130_fd_sc_hd__inv_2 _26842_ (.A(_02338_),
    .Y(_04886_));
 sky130_fd_sc_hd__nor2_2 _26843_ (.A(_19862_),
    .B(_04886_),
    .Y(_04887_));
 sky130_fd_sc_hd__nor2_2 _26844_ (.A(_04885_),
    .B(_04887_),
    .Y(_04888_));
 sky130_fd_sc_hd__inv_2 _26845_ (.A(_02335_),
    .Y(_04889_));
 sky130_fd_sc_hd__o21ai_2 _26846_ (.A1(_19858_),
    .A2(_04889_),
    .B1(_04882_),
    .Y(_04890_));
 sky130_fd_sc_hd__xor2_2 _26847_ (.A(_04888_),
    .B(_04890_),
    .X(_02620_));
 sky130_fd_sc_hd__or2_2 _26848_ (.A(_02339_),
    .B(_04883_),
    .X(_04891_));
 sky130_fd_sc_hd__nand2_2 _26849_ (.A(_04883_),
    .B(_02339_),
    .Y(_04892_));
 sky130_fd_sc_hd__nand2_2 _26850_ (.A(_04891_),
    .B(_04892_),
    .Y(_02340_));
 sky130_fd_sc_hd__or2_2 _26851_ (.A(pcpi_rs1[8]),
    .B(_02341_),
    .X(_04893_));
 sky130_fd_sc_hd__nand2_2 _26852_ (.A(pcpi_rs1[8]),
    .B(_02341_),
    .Y(_04894_));
 sky130_fd_sc_hd__nand2_2 _26853_ (.A(_04893_),
    .B(_04894_),
    .Y(_04895_));
 sky130_fd_sc_hd__inv_2 _26854_ (.A(_04895_),
    .Y(_04896_));
 sky130_fd_sc_hd__and2_2 _26855_ (.A(_04888_),
    .B(_04878_),
    .X(_04897_));
 sky130_fd_sc_hd__o21ai_2 _26856_ (.A1(_04872_),
    .A2(_04879_),
    .B1(_04897_),
    .Y(_04898_));
 sky130_fd_sc_hd__nor2_2 _26857_ (.A(_04889_),
    .B(_04885_),
    .Y(_04899_));
 sky130_fd_sc_hd__a21oi_2 _26858_ (.A1(_04899_),
    .A2(_19528_),
    .B1(_04887_),
    .Y(_04900_));
 sky130_fd_sc_hd__nand2_2 _26859_ (.A(_04898_),
    .B(_04900_),
    .Y(_04901_));
 sky130_fd_sc_hd__or2_2 _26860_ (.A(_04896_),
    .B(_04901_),
    .X(_04902_));
 sky130_fd_sc_hd__nand2_2 _26861_ (.A(_04901_),
    .B(_04896_),
    .Y(_04903_));
 sky130_fd_sc_hd__and2_2 _26862_ (.A(_04902_),
    .B(_04903_),
    .X(_02621_));
 sky130_fd_sc_hd__nor2_2 _26863_ (.A(pcpi_rs2[9]),
    .B(_04892_),
    .Y(_04904_));
 sky130_fd_sc_hd__and2_2 _26864_ (.A(_04892_),
    .B(_19147_),
    .X(_04905_));
 sky130_fd_sc_hd__or2_2 _26865_ (.A(_04904_),
    .B(_04905_),
    .X(_02343_));
 sky130_fd_sc_hd__nor2_2 _26866_ (.A(_19525_),
    .B(_02344_),
    .Y(_04906_));
 sky130_fd_sc_hd__and2_2 _26867_ (.A(_19525_),
    .B(_02344_),
    .X(_04907_));
 sky130_fd_sc_hd__nor2_2 _26868_ (.A(_04906_),
    .B(_04907_),
    .Y(_04908_));
 sky130_fd_sc_hd__nand2_2 _26869_ (.A(_04903_),
    .B(_04894_),
    .Y(_04909_));
 sky130_fd_sc_hd__xor2_2 _26870_ (.A(_04908_),
    .B(_04909_),
    .X(_02622_));
 sky130_fd_sc_hd__or2_2 _26871_ (.A(_02345_),
    .B(_04904_),
    .X(_04910_));
 sky130_fd_sc_hd__nand2_2 _26872_ (.A(_04904_),
    .B(_02345_),
    .Y(_04911_));
 sky130_fd_sc_hd__nand2_2 _26873_ (.A(_04910_),
    .B(_04911_),
    .Y(_02346_));
 sky130_fd_sc_hd__inv_2 _26874_ (.A(_02347_),
    .Y(_04912_));
 sky130_fd_sc_hd__nor2_2 _26875_ (.A(pcpi_rs1[10]),
    .B(_04912_),
    .Y(_04913_));
 sky130_fd_sc_hd__nor2_2 _26876_ (.A(_02347_),
    .B(_19902_),
    .Y(_04914_));
 sky130_fd_sc_hd__or2_2 _26877_ (.A(_04913_),
    .B(_04914_),
    .X(_04915_));
 sky130_fd_sc_hd__o21bai_2 _26878_ (.A1(_04894_),
    .A2(_04906_),
    .B1_N(_04907_),
    .Y(_04916_));
 sky130_fd_sc_hd__nand2_2 _26879_ (.A(_04896_),
    .B(_04908_),
    .Y(_04917_));
 sky130_fd_sc_hd__a21oi_2 _26880_ (.A1(_04898_),
    .A2(_04900_),
    .B1(_04917_),
    .Y(_04918_));
 sky130_fd_sc_hd__nor3_2 _26881_ (.A(_04915_),
    .B(_04916_),
    .C(_04918_),
    .Y(_04919_));
 sky130_fd_sc_hd__o22ai_2 _26882_ (.A1(_04913_),
    .A2(_04914_),
    .B1(_04916_),
    .B2(_04918_),
    .Y(_04920_));
 sky130_fd_sc_hd__nor2b_2 _26883_ (.A(_04919_),
    .B_N(_04920_),
    .Y(_02592_));
 sky130_fd_sc_hd__nor2_2 _26884_ (.A(pcpi_rs2[11]),
    .B(_04911_),
    .Y(_04921_));
 sky130_fd_sc_hd__and2_2 _26885_ (.A(_04911_),
    .B(_19146_),
    .X(_04922_));
 sky130_fd_sc_hd__or2_2 _26886_ (.A(_04921_),
    .B(_04922_),
    .X(_02349_));
 sky130_fd_sc_hd__nor2_2 _26887_ (.A(_19902_),
    .B(_04912_),
    .Y(_04923_));
 sky130_fd_sc_hd__inv_2 _26888_ (.A(_04923_),
    .Y(_04924_));
 sky130_fd_sc_hd__nor2_2 _26889_ (.A(_19524_),
    .B(_02350_),
    .Y(_04925_));
 sky130_fd_sc_hd__and2_2 _26890_ (.A(_19524_),
    .B(_02350_),
    .X(_04926_));
 sky130_fd_sc_hd__or2_2 _26891_ (.A(_04925_),
    .B(_04926_),
    .X(_04927_));
 sky130_fd_sc_hd__a21oi_2 _26892_ (.A1(_04920_),
    .A2(_04924_),
    .B1(_04927_),
    .Y(_04928_));
 sky130_fd_sc_hd__and3_2 _26893_ (.A(_04920_),
    .B(_04924_),
    .C(_04927_),
    .X(_04929_));
 sky130_fd_sc_hd__nor2_2 _26894_ (.A(_04928_),
    .B(_04929_),
    .Y(_02593_));
 sky130_fd_sc_hd__or2_2 _26895_ (.A(_02351_),
    .B(_04921_),
    .X(_04930_));
 sky130_fd_sc_hd__nand2_2 _26896_ (.A(_04921_),
    .B(_02351_),
    .Y(_04931_));
 sky130_fd_sc_hd__nand2_2 _26897_ (.A(_04930_),
    .B(_04931_),
    .Y(_02352_));
 sky130_fd_sc_hd__inv_2 _26898_ (.A(_02353_),
    .Y(_04932_));
 sky130_fd_sc_hd__nor2_2 _26899_ (.A(_19523_),
    .B(_04932_),
    .Y(_04933_));
 sky130_fd_sc_hd__nor2_2 _26900_ (.A(_02353_),
    .B(_19881_),
    .Y(_04934_));
 sky130_fd_sc_hd__or4_2 _26901_ (.A(_04926_),
    .B(_04933_),
    .C(_04934_),
    .D(_04928_),
    .X(_04935_));
 sky130_fd_sc_hd__o22ai_2 _26902_ (.A1(_04933_),
    .A2(_04934_),
    .B1(_04926_),
    .B2(_04928_),
    .Y(_04936_));
 sky130_fd_sc_hd__and2_2 _26903_ (.A(_04935_),
    .B(_04936_),
    .X(_02594_));
 sky130_fd_sc_hd__nor2_2 _26904_ (.A(pcpi_rs2[13]),
    .B(_04931_),
    .Y(_04937_));
 sky130_fd_sc_hd__inv_2 _26905_ (.A(_04937_),
    .Y(_04938_));
 sky130_fd_sc_hd__nand2_2 _26906_ (.A(_04931_),
    .B(_19145_),
    .Y(_04939_));
 sky130_fd_sc_hd__nand2_2 _26907_ (.A(_04938_),
    .B(_04939_),
    .Y(_02355_));
 sky130_fd_sc_hd__nor2_2 _26908_ (.A(_19881_),
    .B(_04932_),
    .Y(_04940_));
 sky130_fd_sc_hd__inv_2 _26909_ (.A(_04940_),
    .Y(_04941_));
 sky130_fd_sc_hd__nor2_2 _26910_ (.A(_19521_),
    .B(_02356_),
    .Y(_04942_));
 sky130_fd_sc_hd__and2_2 _26911_ (.A(_19521_),
    .B(_02356_),
    .X(_04943_));
 sky130_fd_sc_hd__or2_2 _26912_ (.A(_04942_),
    .B(_04943_),
    .X(_04944_));
 sky130_fd_sc_hd__a21oi_2 _26913_ (.A1(_04936_),
    .A2(_04941_),
    .B1(_04944_),
    .Y(_04945_));
 sky130_fd_sc_hd__and3_2 _26914_ (.A(_04936_),
    .B(_04941_),
    .C(_04944_),
    .X(_04946_));
 sky130_fd_sc_hd__nor2_2 _26915_ (.A(_04945_),
    .B(_04946_),
    .Y(_02595_));
 sky130_fd_sc_hd__nand2_2 _26916_ (.A(_04938_),
    .B(_19143_),
    .Y(_04947_));
 sky130_fd_sc_hd__nand2_2 _26917_ (.A(_04937_),
    .B(_02357_),
    .Y(_04948_));
 sky130_fd_sc_hd__nand2_2 _26918_ (.A(_04947_),
    .B(_04948_),
    .Y(_02358_));
 sky130_fd_sc_hd__inv_2 _26919_ (.A(_02359_),
    .Y(_04949_));
 sky130_fd_sc_hd__nor2_2 _26920_ (.A(pcpi_rs1[14]),
    .B(_04949_),
    .Y(_04950_));
 sky130_fd_sc_hd__nor2_2 _26921_ (.A(_02359_),
    .B(_19885_),
    .Y(_04951_));
 sky130_fd_sc_hd__or4_2 _26922_ (.A(_04943_),
    .B(_04950_),
    .C(_04951_),
    .D(_04945_),
    .X(_04952_));
 sky130_fd_sc_hd__o22ai_2 _26923_ (.A1(_04950_),
    .A2(_04951_),
    .B1(_04943_),
    .B2(_04945_),
    .Y(_04953_));
 sky130_fd_sc_hd__and2_2 _26924_ (.A(_04952_),
    .B(_04953_),
    .X(_02596_));
 sky130_fd_sc_hd__nor2_2 _26925_ (.A(pcpi_rs2[15]),
    .B(_04948_),
    .Y(_04954_));
 sky130_fd_sc_hd__and2_2 _26926_ (.A(_04948_),
    .B(_19142_),
    .X(_04955_));
 sky130_fd_sc_hd__or2_2 _26927_ (.A(_04954_),
    .B(_04955_),
    .X(_02361_));
 sky130_fd_sc_hd__nor2_2 _26928_ (.A(_19885_),
    .B(_04949_),
    .Y(_04956_));
 sky130_fd_sc_hd__inv_2 _26929_ (.A(_04956_),
    .Y(_04957_));
 sky130_fd_sc_hd__nor2_2 _26930_ (.A(_19520_),
    .B(_02362_),
    .Y(_04958_));
 sky130_fd_sc_hd__and2_2 _26931_ (.A(_19520_),
    .B(_02362_),
    .X(_04959_));
 sky130_fd_sc_hd__nor2_2 _26932_ (.A(_04958_),
    .B(_04959_),
    .Y(_04960_));
 sky130_fd_sc_hd__inv_2 _26933_ (.A(_04960_),
    .Y(_04961_));
 sky130_fd_sc_hd__a21oi_2 _26934_ (.A1(_04953_),
    .A2(_04957_),
    .B1(_04961_),
    .Y(_04962_));
 sky130_fd_sc_hd__and3_2 _26935_ (.A(_04953_),
    .B(_04957_),
    .C(_04961_),
    .X(_04963_));
 sky130_fd_sc_hd__nor2_2 _26936_ (.A(_04962_),
    .B(_04963_),
    .Y(_02597_));
 sky130_fd_sc_hd__or2_2 _26937_ (.A(_02363_),
    .B(_04954_),
    .X(_04964_));
 sky130_fd_sc_hd__nand2_2 _26938_ (.A(_04954_),
    .B(_02363_),
    .Y(_04965_));
 sky130_fd_sc_hd__nand2_2 _26939_ (.A(_04964_),
    .B(_04965_),
    .Y(_02364_));
 sky130_fd_sc_hd__nor2_2 _26940_ (.A(_19519_),
    .B(_02365_),
    .Y(_04966_));
 sky130_fd_sc_hd__inv_2 _26941_ (.A(_02365_),
    .Y(_04967_));
 sky130_fd_sc_hd__nor2_2 _26942_ (.A(_20237_),
    .B(_04967_),
    .Y(_04968_));
 sky130_fd_sc_hd__or2_2 _26943_ (.A(_04966_),
    .B(_04968_),
    .X(_04969_));
 sky130_fd_sc_hd__nor2_2 _26944_ (.A(_04959_),
    .B(_04962_),
    .Y(_04970_));
 sky130_fd_sc_hd__xor2_2 _26945_ (.A(_04969_),
    .B(_04970_),
    .X(_02598_));
 sky130_fd_sc_hd__or2_2 _26946_ (.A(pcpi_rs2[17]),
    .B(_04965_),
    .X(_04971_));
 sky130_fd_sc_hd__nand2_2 _26947_ (.A(_04965_),
    .B(pcpi_rs2[17]),
    .Y(_04972_));
 sky130_fd_sc_hd__nand2_2 _26948_ (.A(_04971_),
    .B(_04972_),
    .Y(_02367_));
 sky130_fd_sc_hd__nor2_2 _26949_ (.A(_19518_),
    .B(_02368_),
    .Y(_04973_));
 sky130_fd_sc_hd__nand2_2 _26950_ (.A(pcpi_rs1[17]),
    .B(_02368_),
    .Y(_04974_));
 sky130_fd_sc_hd__and2b_2 _26951_ (.A_N(_04973_),
    .B(_04974_),
    .X(_04975_));
 sky130_fd_sc_hd__inv_2 _26952_ (.A(_04975_),
    .Y(_04976_));
 sky130_fd_sc_hd__o21ba_2 _26953_ (.A1(_04966_),
    .A2(_04970_),
    .B1_N(_04968_),
    .X(_04977_));
 sky130_fd_sc_hd__xor2_2 _26954_ (.A(_04976_),
    .B(_04977_),
    .X(_02599_));
 sky130_fd_sc_hd__or2_2 _26955_ (.A(pcpi_rs2[18]),
    .B(_04971_),
    .X(_04978_));
 sky130_fd_sc_hd__nand2_2 _26956_ (.A(_04971_),
    .B(_19141_),
    .Y(_04979_));
 sky130_fd_sc_hd__nand2_2 _26957_ (.A(_04978_),
    .B(_04979_),
    .Y(_02370_));
 sky130_fd_sc_hd__nor2_2 _26958_ (.A(_19517_),
    .B(_02371_),
    .Y(_04980_));
 sky130_fd_sc_hd__and2_2 _26959_ (.A(_19517_),
    .B(_02371_),
    .X(_04981_));
 sky130_fd_sc_hd__nor2_2 _26960_ (.A(_04980_),
    .B(_04981_),
    .Y(_04982_));
 sky130_fd_sc_hd__nor2_2 _26961_ (.A(_04976_),
    .B(_04969_),
    .Y(_04983_));
 sky130_fd_sc_hd__o21ai_2 _26962_ (.A1(_04959_),
    .A2(_04962_),
    .B1(_04983_),
    .Y(_04984_));
 sky130_fd_sc_hd__o31a_2 _26963_ (.A1(_20237_),
    .A2(_04967_),
    .A3(_04973_),
    .B1(_04974_),
    .X(_04985_));
 sky130_fd_sc_hd__nand2_2 _26964_ (.A(_04984_),
    .B(_04985_),
    .Y(_04986_));
 sky130_fd_sc_hd__xor2_2 _26965_ (.A(_04982_),
    .B(_04986_),
    .X(_02600_));
 sky130_fd_sc_hd__nor2_2 _26966_ (.A(pcpi_rs2[19]),
    .B(_04978_),
    .Y(_04987_));
 sky130_fd_sc_hd__and2_2 _26967_ (.A(_04978_),
    .B(pcpi_rs2[19]),
    .X(_04988_));
 sky130_fd_sc_hd__or2_2 _26968_ (.A(_04987_),
    .B(_04988_),
    .X(_02373_));
 sky130_fd_sc_hd__inv_2 _26969_ (.A(_02374_),
    .Y(_04989_));
 sky130_fd_sc_hd__nor2_2 _26970_ (.A(_19515_),
    .B(_04989_),
    .Y(_04990_));
 sky130_fd_sc_hd__nor2_2 _26971_ (.A(_02374_),
    .B(_19988_),
    .Y(_04991_));
 sky130_fd_sc_hd__a21oi_2 _26972_ (.A1(_04984_),
    .A2(_04985_),
    .B1(_04980_),
    .Y(_04992_));
 sky130_fd_sc_hd__or4_2 _26973_ (.A(_04981_),
    .B(_04990_),
    .C(_04991_),
    .D(_04992_),
    .X(_04993_));
 sky130_fd_sc_hd__o22ai_2 _26974_ (.A1(_04990_),
    .A2(_04991_),
    .B1(_04981_),
    .B2(_04992_),
    .Y(_04994_));
 sky130_fd_sc_hd__and2_2 _26975_ (.A(_04993_),
    .B(_04994_),
    .X(_02601_));
 sky130_fd_sc_hd__or2_2 _26976_ (.A(_02375_),
    .B(_04987_),
    .X(_04995_));
 sky130_fd_sc_hd__nand2_2 _26977_ (.A(_04987_),
    .B(_02375_),
    .Y(_04996_));
 sky130_fd_sc_hd__nand2_2 _26978_ (.A(_04995_),
    .B(_04996_),
    .Y(_02376_));
 sky130_fd_sc_hd__nor2_2 _26979_ (.A(_19988_),
    .B(_04989_),
    .Y(_04997_));
 sky130_fd_sc_hd__inv_2 _26980_ (.A(_04997_),
    .Y(_04998_));
 sky130_fd_sc_hd__nor2_2 _26981_ (.A(pcpi_rs1[20]),
    .B(_02377_),
    .Y(_04999_));
 sky130_fd_sc_hd__and2_2 _26982_ (.A(pcpi_rs1[20]),
    .B(_02377_),
    .X(_05000_));
 sky130_fd_sc_hd__nor2_2 _26983_ (.A(_04999_),
    .B(_05000_),
    .Y(_05001_));
 sky130_fd_sc_hd__inv_2 _26984_ (.A(_05001_),
    .Y(_05002_));
 sky130_fd_sc_hd__a21oi_2 _26985_ (.A1(_04994_),
    .A2(_04998_),
    .B1(_05002_),
    .Y(_05003_));
 sky130_fd_sc_hd__and3_2 _26986_ (.A(_04994_),
    .B(_04998_),
    .C(_05002_),
    .X(_05004_));
 sky130_fd_sc_hd__nor2_2 _26987_ (.A(_05003_),
    .B(_05004_),
    .Y(_02603_));
 sky130_fd_sc_hd__or2_2 _26988_ (.A(pcpi_rs2[21]),
    .B(_04996_),
    .X(_05005_));
 sky130_fd_sc_hd__nand2_2 _26989_ (.A(_04996_),
    .B(_19139_),
    .Y(_05006_));
 sky130_fd_sc_hd__nand2_2 _26990_ (.A(_05005_),
    .B(_05006_),
    .Y(_02379_));
 sky130_fd_sc_hd__and2_2 _26991_ (.A(_19926_),
    .B(_02380_),
    .X(_05007_));
 sky130_fd_sc_hd__nor2_2 _26992_ (.A(_02380_),
    .B(_19926_),
    .Y(_05008_));
 sky130_fd_sc_hd__or4_2 _26993_ (.A(_05000_),
    .B(_05007_),
    .C(_05008_),
    .D(_05003_),
    .X(_05009_));
 sky130_fd_sc_hd__o22ai_2 _26994_ (.A1(_05007_),
    .A2(_05008_),
    .B1(_05000_),
    .B2(_05003_),
    .Y(_05010_));
 sky130_fd_sc_hd__and2_2 _26995_ (.A(_05009_),
    .B(_05010_),
    .X(_02604_));
 sky130_fd_sc_hd__or2_2 _26996_ (.A(pcpi_rs2[22]),
    .B(_05005_),
    .X(_05011_));
 sky130_fd_sc_hd__nand2_2 _26997_ (.A(_05005_),
    .B(pcpi_rs2[22]),
    .Y(_05012_));
 sky130_fd_sc_hd__nand2_2 _26998_ (.A(_05011_),
    .B(_05012_),
    .Y(_02382_));
 sky130_fd_sc_hd__nand2_2 _26999_ (.A(_19514_),
    .B(_02380_),
    .Y(_05013_));
 sky130_fd_sc_hd__nor2_2 _27000_ (.A(_19513_),
    .B(_02383_),
    .Y(_05014_));
 sky130_fd_sc_hd__and2_2 _27001_ (.A(_19513_),
    .B(_02383_),
    .X(_05015_));
 sky130_fd_sc_hd__nor2_2 _27002_ (.A(_05014_),
    .B(_05015_),
    .Y(_05016_));
 sky130_fd_sc_hd__a21boi_2 _27003_ (.A1(_05010_),
    .A2(_05013_),
    .B1_N(_05016_),
    .Y(_05017_));
 sky130_fd_sc_hd__o211a_2 _27004_ (.A1(_05015_),
    .A2(_05014_),
    .B1(_05013_),
    .C1(_05010_),
    .X(_05018_));
 sky130_fd_sc_hd__nor2_2 _27005_ (.A(_05017_),
    .B(_05018_),
    .Y(_02605_));
 sky130_fd_sc_hd__nor2_2 _27006_ (.A(_19138_),
    .B(_05011_),
    .Y(_05019_));
 sky130_fd_sc_hd__and2_2 _27007_ (.A(_05011_),
    .B(_19138_),
    .X(_05020_));
 sky130_fd_sc_hd__or2_2 _27008_ (.A(_05019_),
    .B(_05020_),
    .X(_02385_));
 sky130_fd_sc_hd__and2_2 _27009_ (.A(_19930_),
    .B(_02386_),
    .X(_05021_));
 sky130_fd_sc_hd__nor2_2 _27010_ (.A(_02386_),
    .B(_19930_),
    .Y(_05022_));
 sky130_fd_sc_hd__or4_2 _27011_ (.A(_05015_),
    .B(_05021_),
    .C(_05022_),
    .D(_05017_),
    .X(_05023_));
 sky130_fd_sc_hd__o22ai_2 _27012_ (.A1(_05021_),
    .A2(_05022_),
    .B1(_05015_),
    .B2(_05017_),
    .Y(_05024_));
 sky130_fd_sc_hd__and2_2 _27013_ (.A(_05023_),
    .B(_05024_),
    .X(_02606_));
 sky130_fd_sc_hd__or2_2 _27014_ (.A(_02387_),
    .B(_05019_),
    .X(_05025_));
 sky130_fd_sc_hd__nand2_2 _27015_ (.A(_05019_),
    .B(_02387_),
    .Y(_05026_));
 sky130_fd_sc_hd__nand2_2 _27016_ (.A(_05025_),
    .B(_05026_),
    .Y(_02388_));
 sky130_fd_sc_hd__or2_2 _27017_ (.A(pcpi_rs1[24]),
    .B(_02389_),
    .X(_05027_));
 sky130_fd_sc_hd__nand2_2 _27018_ (.A(_19511_),
    .B(_02389_),
    .Y(_05028_));
 sky130_fd_sc_hd__and2_2 _27019_ (.A(_05027_),
    .B(_05028_),
    .X(_05029_));
 sky130_fd_sc_hd__nand2_2 _27020_ (.A(_19512_),
    .B(_02386_),
    .Y(_05030_));
 sky130_fd_sc_hd__nand2_2 _27021_ (.A(_05024_),
    .B(_05030_),
    .Y(_05031_));
 sky130_fd_sc_hd__or2_2 _27022_ (.A(_05029_),
    .B(_05031_),
    .X(_05032_));
 sky130_fd_sc_hd__nand2_2 _27023_ (.A(_05031_),
    .B(_05029_),
    .Y(_05033_));
 sky130_fd_sc_hd__and2_2 _27024_ (.A(_05032_),
    .B(_05033_),
    .X(_02607_));
 sky130_fd_sc_hd__nor2_2 _27025_ (.A(_19137_),
    .B(_05026_),
    .Y(_05034_));
 sky130_fd_sc_hd__inv_2 _27026_ (.A(_05034_),
    .Y(_05035_));
 sky130_fd_sc_hd__nand2_2 _27027_ (.A(_05026_),
    .B(_19137_),
    .Y(_05036_));
 sky130_fd_sc_hd__nand2_2 _27028_ (.A(_05035_),
    .B(_05036_),
    .Y(_02391_));
 sky130_fd_sc_hd__nor2_2 _27029_ (.A(_19509_),
    .B(_02392_),
    .Y(_05037_));
 sky130_fd_sc_hd__inv_2 _27030_ (.A(_05037_),
    .Y(_05038_));
 sky130_fd_sc_hd__nand2_2 _27031_ (.A(_19509_),
    .B(_02392_),
    .Y(_05039_));
 sky130_fd_sc_hd__nand2_2 _27032_ (.A(_05038_),
    .B(_05039_),
    .Y(_05040_));
 sky130_fd_sc_hd__inv_2 _27033_ (.A(_05040_),
    .Y(_05041_));
 sky130_fd_sc_hd__nand2_2 _27034_ (.A(_05033_),
    .B(_05028_),
    .Y(_05042_));
 sky130_fd_sc_hd__xor2_2 _27035_ (.A(_05041_),
    .B(_05042_),
    .X(_02608_));
 sky130_fd_sc_hd__nand2_2 _27036_ (.A(_05035_),
    .B(pcpi_rs2[26]),
    .Y(_05043_));
 sky130_fd_sc_hd__nand2_2 _27037_ (.A(_05034_),
    .B(_02393_),
    .Y(_05044_));
 sky130_fd_sc_hd__nand2_2 _27038_ (.A(_05043_),
    .B(_05044_),
    .Y(_02394_));
 sky130_fd_sc_hd__nor2_2 _27039_ (.A(_19508_),
    .B(_02395_),
    .Y(_05045_));
 sky130_fd_sc_hd__inv_2 _27040_ (.A(_02395_),
    .Y(_05046_));
 sky130_fd_sc_hd__nor2_2 _27041_ (.A(_19952_),
    .B(_05046_),
    .Y(_05047_));
 sky130_fd_sc_hd__nor2_2 _27042_ (.A(_05045_),
    .B(_05047_),
    .Y(_05048_));
 sky130_fd_sc_hd__o21ai_2 _27043_ (.A1(_05028_),
    .A2(_05037_),
    .B1(_05039_),
    .Y(_05049_));
 sky130_fd_sc_hd__nand2_2 _27044_ (.A(_05041_),
    .B(_05029_),
    .Y(_05050_));
 sky130_fd_sc_hd__a21oi_2 _27045_ (.A1(_05024_),
    .A2(_05030_),
    .B1(_05050_),
    .Y(_05051_));
 sky130_fd_sc_hd__or2_2 _27046_ (.A(_05049_),
    .B(_05051_),
    .X(_05052_));
 sky130_fd_sc_hd__xor2_2 _27047_ (.A(_05048_),
    .B(_05052_),
    .X(_02609_));
 sky130_fd_sc_hd__nor2_2 _27048_ (.A(_19135_),
    .B(_05044_),
    .Y(_05053_));
 sky130_fd_sc_hd__and2_2 _27049_ (.A(_05044_),
    .B(_19135_),
    .X(_05054_));
 sky130_fd_sc_hd__or2_2 _27050_ (.A(_05053_),
    .B(_05054_),
    .X(_02397_));
 sky130_fd_sc_hd__nor2_2 _27051_ (.A(pcpi_rs1[27]),
    .B(_02398_),
    .Y(_05055_));
 sky130_fd_sc_hd__inv_2 _27052_ (.A(_02398_),
    .Y(_05056_));
 sky130_fd_sc_hd__nor2_2 _27053_ (.A(_19967_),
    .B(_05056_),
    .Y(_05057_));
 sky130_fd_sc_hd__nor2_2 _27054_ (.A(_05055_),
    .B(_05057_),
    .Y(_05058_));
 sky130_fd_sc_hd__a21oi_2 _27055_ (.A1(_05052_),
    .A2(_05048_),
    .B1(_05047_),
    .Y(_05059_));
 sky130_fd_sc_hd__xnor2_2 _27056_ (.A(_05058_),
    .B(_05059_),
    .Y(_02610_));
 sky130_fd_sc_hd__or2_2 _27057_ (.A(_02399_),
    .B(_05053_),
    .X(_05060_));
 sky130_fd_sc_hd__nand2_2 _27058_ (.A(_05053_),
    .B(_02399_),
    .Y(_05061_));
 sky130_fd_sc_hd__nand2_2 _27059_ (.A(_05060_),
    .B(_05061_),
    .Y(_02400_));
 sky130_fd_sc_hd__and2_2 _27060_ (.A(_05048_),
    .B(_05058_),
    .X(_05062_));
 sky130_fd_sc_hd__o21ai_2 _27061_ (.A1(_05049_),
    .A2(_05051_),
    .B1(_05062_),
    .Y(_05063_));
 sky130_fd_sc_hd__nor2_2 _27062_ (.A(_05046_),
    .B(_05055_),
    .Y(_05064_));
 sky130_fd_sc_hd__a21oi_2 _27063_ (.A1(_05064_),
    .A2(_19508_),
    .B1(_05057_),
    .Y(_05065_));
 sky130_fd_sc_hd__nor2_2 _27064_ (.A(_19507_),
    .B(_02401_),
    .Y(_05066_));
 sky130_fd_sc_hd__inv_2 _27065_ (.A(_02401_),
    .Y(_05067_));
 sky130_fd_sc_hd__nor2_2 _27066_ (.A(_19949_),
    .B(_05067_),
    .Y(_05068_));
 sky130_fd_sc_hd__or2_2 _27067_ (.A(_05066_),
    .B(_05068_),
    .X(_05069_));
 sky130_fd_sc_hd__a21oi_2 _27068_ (.A1(_05063_),
    .A2(_05065_),
    .B1(_05069_),
    .Y(_05070_));
 sky130_fd_sc_hd__and3_2 _27069_ (.A(_05063_),
    .B(_05065_),
    .C(_05069_),
    .X(_05071_));
 sky130_fd_sc_hd__nor2_2 _27070_ (.A(_05070_),
    .B(_05071_),
    .Y(_02611_));
 sky130_fd_sc_hd__or2_2 _27071_ (.A(_19134_),
    .B(_05061_),
    .X(_05072_));
 sky130_fd_sc_hd__nand2_2 _27072_ (.A(_05061_),
    .B(_19134_),
    .Y(_05073_));
 sky130_fd_sc_hd__nand2_2 _27073_ (.A(_05072_),
    .B(_05073_),
    .Y(_02403_));
 sky130_fd_sc_hd__or2_2 _27074_ (.A(pcpi_rs1[29]),
    .B(_02404_),
    .X(_05074_));
 sky130_fd_sc_hd__nand2_2 _27075_ (.A(_19506_),
    .B(_02404_),
    .Y(_05075_));
 sky130_fd_sc_hd__nand2_2 _27076_ (.A(_05074_),
    .B(_05075_),
    .Y(_05076_));
 sky130_fd_sc_hd__a22oi_2 _27077_ (.A1(_19949_),
    .A2(_05067_),
    .B1(_05063_),
    .B2(_05065_),
    .Y(_05077_));
 sky130_fd_sc_hd__or3_2 _27078_ (.A(_05068_),
    .B(_05076_),
    .C(_05077_),
    .X(_05078_));
 sky130_fd_sc_hd__o21ai_2 _27079_ (.A1(_05068_),
    .A2(_05077_),
    .B1(_05076_),
    .Y(_05079_));
 sky130_fd_sc_hd__nand2_2 _27080_ (.A(_05078_),
    .B(_05079_),
    .Y(_02612_));
 sky130_fd_sc_hd__nor2_2 _27081_ (.A(pcpi_rs2[30]),
    .B(_05072_),
    .Y(_05080_));
 sky130_fd_sc_hd__and2_2 _27082_ (.A(_05072_),
    .B(pcpi_rs2[30]),
    .X(_05081_));
 sky130_fd_sc_hd__or2_2 _27083_ (.A(_05080_),
    .B(_05081_),
    .X(_02406_));
 sky130_fd_sc_hd__o22ai_2 _27084_ (.A1(_19506_),
    .A2(_02404_),
    .B1(_05068_),
    .B2(_05077_),
    .Y(_05082_));
 sky130_fd_sc_hd__nor2_2 _27085_ (.A(_19505_),
    .B(_02407_),
    .Y(_05083_));
 sky130_fd_sc_hd__and2_2 _27086_ (.A(_19505_),
    .B(_02407_),
    .X(_05084_));
 sky130_fd_sc_hd__nor2_2 _27087_ (.A(_05083_),
    .B(_05084_),
    .Y(_05085_));
 sky130_fd_sc_hd__inv_2 _27088_ (.A(_05085_),
    .Y(_05086_));
 sky130_fd_sc_hd__a21oi_2 _27089_ (.A1(_05082_),
    .A2(_05075_),
    .B1(_05086_),
    .Y(_05087_));
 sky130_fd_sc_hd__nand2_2 _27090_ (.A(_05082_),
    .B(_05075_),
    .Y(_05088_));
 sky130_fd_sc_hd__nor2_2 _27091_ (.A(_05085_),
    .B(_05088_),
    .Y(_05089_));
 sky130_fd_sc_hd__nor2_2 _27092_ (.A(_05087_),
    .B(_05089_),
    .Y(_02614_));
 sky130_fd_sc_hd__xor2_2 _27093_ (.A(_19971_),
    .B(_05080_),
    .X(_02408_));
 sky130_fd_sc_hd__and2_2 _27094_ (.A(_18173_),
    .B(_02409_),
    .X(_05090_));
 sky130_fd_sc_hd__nor2_2 _27095_ (.A(_02409_),
    .B(_18173_),
    .Y(_05091_));
 sky130_fd_sc_hd__o22ai_2 _27096_ (.A1(_05090_),
    .A2(_05091_),
    .B1(_05084_),
    .B2(_05087_),
    .Y(_05092_));
 sky130_fd_sc_hd__or3_2 _27097_ (.A(_05084_),
    .B(_05091_),
    .C(_05090_),
    .X(_05093_));
 sky130_fd_sc_hd__a21o_2 _27098_ (.A1(_05088_),
    .A2(_05085_),
    .B1(_05093_),
    .X(_05094_));
 sky130_fd_sc_hd__nand2_2 _27099_ (.A(_05092_),
    .B(_05094_),
    .Y(_02615_));
 sky130_fd_sc_hd__nand2_2 _27100_ (.A(_19404_),
    .B(_19638_),
    .Y(_05095_));
 sky130_fd_sc_hd__nand2_2 _27101_ (.A(_19402_),
    .B(_19642_),
    .Y(_05096_));
 sky130_fd_sc_hd__nor2_2 _27102_ (.A(_05095_),
    .B(_05096_),
    .Y(_05097_));
 sky130_fd_sc_hd__and2_2 _27103_ (.A(_05095_),
    .B(_05096_),
    .X(_05098_));
 sky130_fd_sc_hd__nor2_2 _27104_ (.A(_05097_),
    .B(_05098_),
    .Y(_02624_));
 sky130_fd_sc_hd__inv_2 _27105_ (.A(_05097_),
    .Y(_05099_));
 sky130_fd_sc_hd__inv_2 _27106_ (.A(\pcpi_mul.rs1[2] ),
    .Y(_05100_));
 sky130_fd_sc_hd__buf_1 _27107_ (.A(_05100_),
    .X(_05101_));
 sky130_fd_sc_hd__nand2_2 _27108_ (.A(\pcpi_mul.rs2[2] ),
    .B(\pcpi_mul.rs2[1] ),
    .Y(_05102_));
 sky130_fd_sc_hd__buf_1 _27109_ (.A(_05102_),
    .X(_05103_));
 sky130_fd_sc_hd__buf_1 _27110_ (.A(\pcpi_mul.rs1[1] ),
    .X(_05104_));
 sky130_fd_sc_hd__buf_1 _27111_ (.A(_05104_),
    .X(_05105_));
 sky130_fd_sc_hd__inv_2 _27112_ (.A(_05105_),
    .Y(_05106_));
 sky130_fd_sc_hd__or3_2 _27113_ (.A(_05103_),
    .B(_05106_),
    .C(_04839_),
    .X(_05107_));
 sky130_fd_sc_hd__a22o_2 _27114_ (.A1(_19399_),
    .A2(_19642_),
    .B1(_19402_),
    .B2(_19638_),
    .X(_05108_));
 sky130_fd_sc_hd__nand2_2 _27115_ (.A(_05107_),
    .B(_05108_),
    .Y(_05109_));
 sky130_fd_sc_hd__or3_2 _27116_ (.A(_04836_),
    .B(_05101_),
    .C(_05109_),
    .X(_05110_));
 sky130_fd_sc_hd__o21ai_2 _27117_ (.A1(_04836_),
    .A2(_05101_),
    .B1(_05109_),
    .Y(_05111_));
 sky130_fd_sc_hd__nand2_2 _27118_ (.A(_05110_),
    .B(_05111_),
    .Y(_05112_));
 sky130_fd_sc_hd__nor2_2 _27119_ (.A(_05099_),
    .B(_05112_),
    .Y(_05113_));
 sky130_fd_sc_hd__and2_2 _27120_ (.A(_05112_),
    .B(_05099_),
    .X(_05114_));
 sky130_fd_sc_hd__nor2_2 _27121_ (.A(_05113_),
    .B(_05114_),
    .Y(_02625_));
 sky130_fd_sc_hd__buf_1 _27122_ (.A(\pcpi_mul.rs2[3] ),
    .X(_05115_));
 sky130_fd_sc_hd__buf_1 _27123_ (.A(_05115_),
    .X(_05116_));
 sky130_fd_sc_hd__nand2_2 _27124_ (.A(_05116_),
    .B(_19641_),
    .Y(_05117_));
 sky130_fd_sc_hd__buf_1 _27125_ (.A(_19400_),
    .X(_05118_));
 sky130_fd_sc_hd__buf_1 _27126_ (.A(_19632_),
    .X(_05119_));
 sky130_fd_sc_hd__buf_1 _27127_ (.A(_05119_),
    .X(_05120_));
 sky130_fd_sc_hd__nand2_2 _27128_ (.A(_05118_),
    .B(_05120_),
    .Y(_05121_));
 sky130_fd_sc_hd__buf_1 _27129_ (.A(\pcpi_mul.rs2[2] ),
    .X(_05122_));
 sky130_fd_sc_hd__buf_1 _27130_ (.A(_05122_),
    .X(_05123_));
 sky130_fd_sc_hd__buf_1 _27131_ (.A(_05105_),
    .X(_05124_));
 sky130_fd_sc_hd__nand2_2 _27132_ (.A(_05123_),
    .B(_05124_),
    .Y(_05125_));
 sky130_fd_sc_hd__nor2_2 _27133_ (.A(_05121_),
    .B(_05125_),
    .Y(_05126_));
 sky130_fd_sc_hd__nand2_2 _27134_ (.A(_05121_),
    .B(_05125_),
    .Y(_05127_));
 sky130_fd_sc_hd__or3b_2 _27135_ (.A(_05117_),
    .B(_05126_),
    .C_N(_05127_),
    .X(_05128_));
 sky130_fd_sc_hd__inv_2 _27136_ (.A(_05126_),
    .Y(_05129_));
 sky130_fd_sc_hd__a21bo_2 _27137_ (.A1(_05129_),
    .A2(_05127_),
    .B1_N(_05117_),
    .X(_05130_));
 sky130_fd_sc_hd__nand2_2 _27138_ (.A(_19404_),
    .B(_19631_),
    .Y(_05131_));
 sky130_fd_sc_hd__inv_2 _27139_ (.A(_05131_),
    .Y(_05132_));
 sky130_fd_sc_hd__a21o_2 _27140_ (.A1(_05128_),
    .A2(_05130_),
    .B1(_05132_),
    .X(_05133_));
 sky130_fd_sc_hd__nand3_2 _27141_ (.A(_05128_),
    .B(_05130_),
    .C(_05132_),
    .Y(_05134_));
 sky130_fd_sc_hd__nand2_2 _27142_ (.A(_05133_),
    .B(_05134_),
    .Y(_05135_));
 sky130_fd_sc_hd__nand3_2 _27143_ (.A(_05135_),
    .B(_05107_),
    .C(_05110_),
    .Y(_05136_));
 sky130_fd_sc_hd__a21oi_2 _27144_ (.A1(_05107_),
    .A2(_05110_),
    .B1(_05135_),
    .Y(_05137_));
 sky130_fd_sc_hd__inv_2 _27145_ (.A(_05137_),
    .Y(_05138_));
 sky130_fd_sc_hd__a21oi_2 _27146_ (.A1(_05136_),
    .A2(_05138_),
    .B1(_05113_),
    .Y(_05139_));
 sky130_fd_sc_hd__nand3_2 _27147_ (.A(_05138_),
    .B(_05113_),
    .C(_05136_),
    .Y(_05140_));
 sky130_fd_sc_hd__nor2b_2 _27148_ (.A(_05139_),
    .B_N(_05140_),
    .Y(_02626_));
 sky130_fd_sc_hd__buf_1 _27149_ (.A(_19398_),
    .X(_05141_));
 sky130_fd_sc_hd__buf_1 _27150_ (.A(\pcpi_mul.rs2[1] ),
    .X(_05142_));
 sky130_fd_sc_hd__buf_1 _27151_ (.A(_05142_),
    .X(_05143_));
 sky130_fd_sc_hd__buf_1 _27152_ (.A(_05143_),
    .X(_05144_));
 sky130_fd_sc_hd__a22o_2 _27153_ (.A1(_05141_),
    .A2(_19634_),
    .B1(_05144_),
    .B2(_19631_),
    .X(_05145_));
 sky130_fd_sc_hd__buf_1 _27154_ (.A(\pcpi_mul.rs1[3] ),
    .X(_05146_));
 sky130_fd_sc_hd__nand2_2 _27155_ (.A(_05146_),
    .B(\pcpi_mul.rs1[2] ),
    .Y(_05147_));
 sky130_fd_sc_hd__or2_2 _27156_ (.A(_05102_),
    .B(_05147_),
    .X(_05148_));
 sky130_fd_sc_hd__inv_2 _27157_ (.A(\pcpi_mul.rs2[3] ),
    .Y(_05149_));
 sky130_fd_sc_hd__buf_1 _27158_ (.A(_05149_),
    .X(_05150_));
 sky130_fd_sc_hd__buf_1 _27159_ (.A(_05150_),
    .X(_05151_));
 sky130_fd_sc_hd__o2bb2ai_2 _27160_ (.A1_N(_05145_),
    .A2_N(_05148_),
    .B1(_05151_),
    .B2(_05106_),
    .Y(_05152_));
 sky130_fd_sc_hd__o2111ai_2 _27161_ (.A1(_05103_),
    .A2(_05147_),
    .B1(_19395_),
    .C1(_19638_),
    .D1(_05145_),
    .Y(_05153_));
 sky130_fd_sc_hd__nand2_2 _27162_ (.A(_05152_),
    .B(_05153_),
    .Y(_05154_));
 sky130_fd_sc_hd__buf_1 _27163_ (.A(\pcpi_mul.rs2[4] ),
    .X(_05155_));
 sky130_fd_sc_hd__nand2_2 _27164_ (.A(_05155_),
    .B(_19639_),
    .Y(_05156_));
 sky130_fd_sc_hd__buf_1 _27165_ (.A(\pcpi_mul.rs2[0] ),
    .X(_05157_));
 sky130_fd_sc_hd__buf_1 _27166_ (.A(\pcpi_mul.rs1[4] ),
    .X(_05158_));
 sky130_fd_sc_hd__nand2_2 _27167_ (.A(_05157_),
    .B(_05158_),
    .Y(_05159_));
 sky130_fd_sc_hd__nor2_2 _27168_ (.A(_05156_),
    .B(_05159_),
    .Y(_05160_));
 sky130_fd_sc_hd__inv_2 _27169_ (.A(_05160_),
    .Y(_05161_));
 sky130_fd_sc_hd__nand2_2 _27170_ (.A(_05156_),
    .B(_05159_),
    .Y(_05162_));
 sky130_fd_sc_hd__nand2_2 _27171_ (.A(_05161_),
    .B(_05162_),
    .Y(_05163_));
 sky130_fd_sc_hd__nand2_2 _27172_ (.A(_05154_),
    .B(_05163_),
    .Y(_05164_));
 sky130_fd_sc_hd__nand3b_2 _27173_ (.A_N(_05163_),
    .B(_05152_),
    .C(_05153_),
    .Y(_05165_));
 sky130_fd_sc_hd__nand2_2 _27174_ (.A(_05164_),
    .B(_05165_),
    .Y(_05166_));
 sky130_fd_sc_hd__nand2_2 _27175_ (.A(_05166_),
    .B(_05134_),
    .Y(_05167_));
 sky130_fd_sc_hd__nand3b_2 _27176_ (.A_N(_05134_),
    .B(_05164_),
    .C(_05165_),
    .Y(_05168_));
 sky130_fd_sc_hd__nand2_2 _27177_ (.A(_05167_),
    .B(_05168_),
    .Y(_05169_));
 sky130_fd_sc_hd__nand2_2 _27178_ (.A(_05128_),
    .B(_05129_),
    .Y(_05170_));
 sky130_fd_sc_hd__inv_2 _27179_ (.A(_05170_),
    .Y(_05171_));
 sky130_fd_sc_hd__nand2_2 _27180_ (.A(_05169_),
    .B(_05171_),
    .Y(_05172_));
 sky130_fd_sc_hd__nand3_2 _27181_ (.A(_05167_),
    .B(_05168_),
    .C(_05170_),
    .Y(_05173_));
 sky130_fd_sc_hd__nand2_2 _27182_ (.A(_05172_),
    .B(_05173_),
    .Y(_05174_));
 sky130_fd_sc_hd__inv_2 _27183_ (.A(_05174_),
    .Y(_05175_));
 sky130_fd_sc_hd__nand2_2 _27184_ (.A(_05140_),
    .B(_05138_),
    .Y(_05176_));
 sky130_fd_sc_hd__or2_2 _27185_ (.A(_05175_),
    .B(_05176_),
    .X(_05177_));
 sky130_fd_sc_hd__nand2_2 _27186_ (.A(_05176_),
    .B(_05175_),
    .Y(_05178_));
 sky130_fd_sc_hd__and2_2 _27187_ (.A(_05177_),
    .B(_05178_),
    .X(_02627_));
 sky130_fd_sc_hd__nand2_2 _27188_ (.A(_19390_),
    .B(_19635_),
    .Y(_05179_));
 sky130_fd_sc_hd__buf_1 _27189_ (.A(\pcpi_mul.rs2[5] ),
    .X(_05180_));
 sky130_fd_sc_hd__nand2_2 _27190_ (.A(_05180_),
    .B(_19639_),
    .Y(_05181_));
 sky130_fd_sc_hd__nor2_2 _27191_ (.A(_05179_),
    .B(_05181_),
    .Y(_05182_));
 sky130_fd_sc_hd__nand2_2 _27192_ (.A(_05179_),
    .B(_05181_),
    .Y(_05183_));
 sky130_fd_sc_hd__buf_1 _27193_ (.A(_19624_),
    .X(_05184_));
 sky130_fd_sc_hd__and2_2 _27194_ (.A(_04834_),
    .B(_05184_),
    .X(_05185_));
 sky130_fd_sc_hd__nand3b_2 _27195_ (.A_N(_05182_),
    .B(_05183_),
    .C(_05185_),
    .Y(_05186_));
 sky130_fd_sc_hd__buf_1 _27196_ (.A(_19387_),
    .X(_05187_));
 sky130_fd_sc_hd__buf_1 _27197_ (.A(\pcpi_mul.rs1[0] ),
    .X(_05188_));
 sky130_fd_sc_hd__buf_1 _27198_ (.A(_19390_),
    .X(_05189_));
 sky130_fd_sc_hd__buf_1 _27199_ (.A(_05104_),
    .X(_05190_));
 sky130_fd_sc_hd__a22oi_2 _27200_ (.A1(_05187_),
    .A2(_05188_),
    .B1(_05189_),
    .B2(_05190_),
    .Y(_05191_));
 sky130_fd_sc_hd__buf_1 _27201_ (.A(_05157_),
    .X(_05192_));
 sky130_fd_sc_hd__buf_1 _27202_ (.A(\pcpi_mul.rs1[5] ),
    .X(_05193_));
 sky130_fd_sc_hd__buf_1 _27203_ (.A(_05193_),
    .X(_05194_));
 sky130_fd_sc_hd__nand2_2 _27204_ (.A(_05192_),
    .B(_05194_),
    .Y(_05195_));
 sky130_fd_sc_hd__o21ai_2 _27205_ (.A1(_05191_),
    .A2(_05182_),
    .B1(_05195_),
    .Y(_05196_));
 sky130_fd_sc_hd__nand3_2 _27206_ (.A(_05186_),
    .B(_05160_),
    .C(_05196_),
    .Y(_05197_));
 sky130_fd_sc_hd__o21ai_2 _27207_ (.A1(_05191_),
    .A2(_05182_),
    .B1(_05185_),
    .Y(_05198_));
 sky130_fd_sc_hd__nand3_2 _27208_ (.A(_05187_),
    .B(_05189_),
    .C(_05105_),
    .Y(_05199_));
 sky130_fd_sc_hd__o211ai_2 _27209_ (.A1(_04838_),
    .A2(_05199_),
    .B1(_05195_),
    .C1(_05183_),
    .Y(_05200_));
 sky130_fd_sc_hd__nand3_2 _27210_ (.A(_05198_),
    .B(_05161_),
    .C(_05200_),
    .Y(_05201_));
 sky130_fd_sc_hd__nand2_2 _27211_ (.A(_05197_),
    .B(_05201_),
    .Y(_05202_));
 sky130_fd_sc_hd__buf_1 _27212_ (.A(_19397_),
    .X(_05203_));
 sky130_fd_sc_hd__buf_1 _27213_ (.A(_19629_),
    .X(_05204_));
 sky130_fd_sc_hd__buf_1 _27214_ (.A(_05142_),
    .X(_05205_));
 sky130_fd_sc_hd__buf_1 _27215_ (.A(\pcpi_mul.rs1[4] ),
    .X(_05206_));
 sky130_fd_sc_hd__buf_1 _27216_ (.A(_05206_),
    .X(_05207_));
 sky130_fd_sc_hd__a22oi_2 _27217_ (.A1(_05203_),
    .A2(_05204_),
    .B1(_05205_),
    .B2(_05207_),
    .Y(_05208_));
 sky130_fd_sc_hd__buf_1 _27218_ (.A(_19397_),
    .X(_05209_));
 sky130_fd_sc_hd__buf_1 _27219_ (.A(_05142_),
    .X(_05210_));
 sky130_fd_sc_hd__buf_1 _27220_ (.A(\pcpi_mul.rs1[4] ),
    .X(_05211_));
 sky130_fd_sc_hd__buf_1 _27221_ (.A(_05211_),
    .X(_05212_));
 sky130_fd_sc_hd__buf_1 _27222_ (.A(_19629_),
    .X(_05213_));
 sky130_fd_sc_hd__and4_2 _27223_ (.A(_05209_),
    .B(_05210_),
    .C(_05212_),
    .D(_05213_),
    .X(_05214_));
 sky130_fd_sc_hd__buf_1 _27224_ (.A(_19632_),
    .X(_05215_));
 sky130_fd_sc_hd__nand2_2 _27225_ (.A(\pcpi_mul.rs2[3] ),
    .B(_05215_),
    .Y(_05216_));
 sky130_fd_sc_hd__o21bai_2 _27226_ (.A1(_05208_),
    .A2(_05214_),
    .B1_N(_05216_),
    .Y(_05217_));
 sky130_fd_sc_hd__buf_1 _27227_ (.A(_05146_),
    .X(_05218_));
 sky130_fd_sc_hd__nand2_2 _27228_ (.A(_05122_),
    .B(_05218_),
    .Y(_05219_));
 sky130_fd_sc_hd__nand3b_2 _27229_ (.A_N(_05219_),
    .B(_05205_),
    .C(_05207_),
    .Y(_05220_));
 sky130_fd_sc_hd__buf_1 _27230_ (.A(_05142_),
    .X(_05221_));
 sky130_fd_sc_hd__buf_1 _27231_ (.A(_05211_),
    .X(_05222_));
 sky130_fd_sc_hd__a22o_2 _27232_ (.A1(_05209_),
    .A2(_05213_),
    .B1(_05221_),
    .B2(_05222_),
    .X(_05223_));
 sky130_fd_sc_hd__nand3_2 _27233_ (.A(_05220_),
    .B(_05216_),
    .C(_05223_),
    .Y(_05224_));
 sky130_fd_sc_hd__and2_2 _27234_ (.A(_05217_),
    .B(_05224_),
    .X(_05225_));
 sky130_fd_sc_hd__nand2_2 _27235_ (.A(_05202_),
    .B(_05225_),
    .Y(_05226_));
 sky130_fd_sc_hd__nand2_2 _27236_ (.A(_05217_),
    .B(_05224_),
    .Y(_05227_));
 sky130_fd_sc_hd__nand3_2 _27237_ (.A(_05197_),
    .B(_05227_),
    .C(_05201_),
    .Y(_05228_));
 sky130_fd_sc_hd__nand3b_2 _27238_ (.A_N(_05165_),
    .B(_05226_),
    .C(_05228_),
    .Y(_05229_));
 sky130_fd_sc_hd__nand2_2 _27239_ (.A(_05202_),
    .B(_05227_),
    .Y(_05230_));
 sky130_fd_sc_hd__nand3_2 _27240_ (.A(_05225_),
    .B(_05197_),
    .C(_05201_),
    .Y(_05231_));
 sky130_fd_sc_hd__nand3_2 _27241_ (.A(_05230_),
    .B(_05165_),
    .C(_05231_),
    .Y(_05232_));
 sky130_fd_sc_hd__nor2_2 _27242_ (.A(_05103_),
    .B(_05147_),
    .Y(_05233_));
 sky130_fd_sc_hd__a31o_2 _27243_ (.A1(_05145_),
    .A2(_19395_),
    .A3(_19638_),
    .B1(_05233_),
    .X(_05234_));
 sky130_fd_sc_hd__a21o_2 _27244_ (.A1(_05229_),
    .A2(_05232_),
    .B1(_05234_),
    .X(_05235_));
 sky130_fd_sc_hd__a21boi_2 _27245_ (.A1(_05164_),
    .A2(_05165_),
    .B1_N(_05134_),
    .Y(_05236_));
 sky130_fd_sc_hd__o21ai_2 _27246_ (.A1(_05171_),
    .A2(_05236_),
    .B1(_05168_),
    .Y(_05237_));
 sky130_fd_sc_hd__nand3_2 _27247_ (.A(_05229_),
    .B(_05232_),
    .C(_05234_),
    .Y(_05238_));
 sky130_fd_sc_hd__nand3_2 _27248_ (.A(_05235_),
    .B(_05237_),
    .C(_05238_),
    .Y(_05239_));
 sky130_fd_sc_hd__inv_2 _27249_ (.A(_05239_),
    .Y(_05240_));
 sky130_fd_sc_hd__nand3_2 _27250_ (.A(_05172_),
    .B(_05137_),
    .C(_05173_),
    .Y(_05241_));
 sky130_fd_sc_hd__a21oi_2 _27251_ (.A1(_05235_),
    .A2(_05238_),
    .B1(_05237_),
    .Y(_05242_));
 sky130_fd_sc_hd__nor2_2 _27252_ (.A(_05241_),
    .B(_05242_),
    .Y(_05243_));
 sky130_fd_sc_hd__inv_2 _27253_ (.A(_19385_),
    .Y(_05244_));
 sky130_fd_sc_hd__nand2_2 _27254_ (.A(_05220_),
    .B(_05216_),
    .Y(_05245_));
 sky130_fd_sc_hd__a22oi_2 _27255_ (.A1(_05187_),
    .A2(_05105_),
    .B1(_05189_),
    .B2(_05119_),
    .Y(_05246_));
 sky130_fd_sc_hd__nand2_2 _27256_ (.A(_05180_),
    .B(_19635_),
    .Y(_05247_));
 sky130_fd_sc_hd__buf_1 _27257_ (.A(\pcpi_mul.rs1[2] ),
    .X(_05248_));
 sky130_fd_sc_hd__nand2_2 _27258_ (.A(_05155_),
    .B(_05248_),
    .Y(_05249_));
 sky130_fd_sc_hd__nor2_2 _27259_ (.A(_05247_),
    .B(_05249_),
    .Y(_05250_));
 sky130_fd_sc_hd__buf_1 _27260_ (.A(\pcpi_mul.rs1[6] ),
    .X(_05251_));
 sky130_fd_sc_hd__nand2_2 _27261_ (.A(_05157_),
    .B(_05251_),
    .Y(_05252_));
 sky130_fd_sc_hd__inv_2 _27262_ (.A(_05252_),
    .Y(_05253_));
 sky130_fd_sc_hd__o21ai_2 _27263_ (.A1(_05246_),
    .A2(_05250_),
    .B1(_05253_),
    .Y(_05254_));
 sky130_fd_sc_hd__a21oi_2 _27264_ (.A1(_05183_),
    .A2(_05185_),
    .B1(_05182_),
    .Y(_05255_));
 sky130_fd_sc_hd__buf_1 _27265_ (.A(_05100_),
    .X(_05256_));
 sky130_fd_sc_hd__nand2_2 _27266_ (.A(_05247_),
    .B(_05249_),
    .Y(_05257_));
 sky130_fd_sc_hd__o211ai_2 _27267_ (.A1(_05256_),
    .A2(_05199_),
    .B1(_05252_),
    .C1(_05257_),
    .Y(_05258_));
 sky130_fd_sc_hd__nand3_2 _27268_ (.A(_05254_),
    .B(_05255_),
    .C(_05258_),
    .Y(_05259_));
 sky130_fd_sc_hd__inv_2 _27269_ (.A(_19621_),
    .Y(_05260_));
 sky130_fd_sc_hd__buf_1 _27270_ (.A(_05260_),
    .X(_05261_));
 sky130_fd_sc_hd__o22ai_2 _27271_ (.A1(_04835_),
    .A2(_05261_),
    .B1(_05246_),
    .B2(_05250_),
    .Y(_05262_));
 sky130_fd_sc_hd__o211ai_2 _27272_ (.A1(_05256_),
    .A2(_05199_),
    .B1(_05257_),
    .C1(_05253_),
    .Y(_05263_));
 sky130_fd_sc_hd__o22ai_2 _27273_ (.A1(_04837_),
    .A2(_05199_),
    .B1(_05195_),
    .B2(_05191_),
    .Y(_05264_));
 sky130_fd_sc_hd__nand3_2 _27274_ (.A(_05262_),
    .B(_05263_),
    .C(_05264_),
    .Y(_05265_));
 sky130_fd_sc_hd__nand2_2 _27275_ (.A(_19624_),
    .B(_05211_),
    .Y(_05266_));
 sky130_fd_sc_hd__nor2_2 _27276_ (.A(_05102_),
    .B(_05266_),
    .Y(_05267_));
 sky130_fd_sc_hd__buf_1 _27277_ (.A(_19397_),
    .X(_05268_));
 sky130_fd_sc_hd__buf_1 _27278_ (.A(_05193_),
    .X(_05269_));
 sky130_fd_sc_hd__a22o_2 _27279_ (.A1(_05268_),
    .A2(_05222_),
    .B1(_05221_),
    .B2(_05269_),
    .X(_05270_));
 sky130_fd_sc_hd__buf_1 _27280_ (.A(_05146_),
    .X(_05271_));
 sky130_fd_sc_hd__nand2_2 _27281_ (.A(\pcpi_mul.rs2[3] ),
    .B(_05271_),
    .Y(_05272_));
 sky130_fd_sc_hd__nand3b_2 _27282_ (.A_N(_05267_),
    .B(_05270_),
    .C(_05272_),
    .Y(_05273_));
 sky130_fd_sc_hd__a22oi_2 _27283_ (.A1(_05209_),
    .A2(_05212_),
    .B1(_05210_),
    .B2(_05194_),
    .Y(_05274_));
 sky130_fd_sc_hd__buf_1 _27284_ (.A(_05267_),
    .X(_05275_));
 sky130_fd_sc_hd__inv_2 _27285_ (.A(_05272_),
    .Y(_05276_));
 sky130_fd_sc_hd__o21ai_2 _27286_ (.A1(_05274_),
    .A2(_05275_),
    .B1(_05276_),
    .Y(_05277_));
 sky130_fd_sc_hd__nand2_2 _27287_ (.A(_05273_),
    .B(_05277_),
    .Y(_05278_));
 sky130_fd_sc_hd__a21oi_2 _27288_ (.A1(_05259_),
    .A2(_05265_),
    .B1(_05278_),
    .Y(_05279_));
 sky130_fd_sc_hd__nor3_2 _27289_ (.A(_05274_),
    .B(_05276_),
    .C(_05275_),
    .Y(_05280_));
 sky130_fd_sc_hd__o21a_2 _27290_ (.A1(_05274_),
    .A2(_05275_),
    .B1(_05276_),
    .X(_05281_));
 sky130_fd_sc_hd__o211a_2 _27291_ (.A1(_05280_),
    .A2(_05281_),
    .B1(_05265_),
    .C1(_05259_),
    .X(_05282_));
 sky130_fd_sc_hd__o21a_2 _27292_ (.A1(_05191_),
    .A2(_05182_),
    .B1(_05195_),
    .X(_05283_));
 sky130_fd_sc_hd__nand2_2 _27293_ (.A(_05186_),
    .B(_05160_),
    .Y(_05284_));
 sky130_fd_sc_hd__o2bb2ai_2 _27294_ (.A1_N(_05227_),
    .A2_N(_05201_),
    .B1(_05283_),
    .B2(_05284_),
    .Y(_05285_));
 sky130_fd_sc_hd__o21bai_2 _27295_ (.A1(_05279_),
    .A2(_05282_),
    .B1_N(_05285_),
    .Y(_05286_));
 sky130_fd_sc_hd__nor3_2 _27296_ (.A(_05272_),
    .B(_05274_),
    .C(_05275_),
    .Y(_05287_));
 sky130_fd_sc_hd__o21a_2 _27297_ (.A1(_05274_),
    .A2(_05275_),
    .B1(_05272_),
    .X(_05288_));
 sky130_fd_sc_hd__o2bb2ai_2 _27298_ (.A1_N(_05265_),
    .A2_N(_05259_),
    .B1(_05287_),
    .B2(_05288_),
    .Y(_05289_));
 sky130_fd_sc_hd__nand3_2 _27299_ (.A(_05278_),
    .B(_05259_),
    .C(_05265_),
    .Y(_05290_));
 sky130_fd_sc_hd__nand3_2 _27300_ (.A(_05285_),
    .B(_05289_),
    .C(_05290_),
    .Y(_05291_));
 sky130_fd_sc_hd__a22oi_2 _27301_ (.A1(_05223_),
    .A2(_05245_),
    .B1(_05286_),
    .B2(_05291_),
    .Y(_05292_));
 sky130_fd_sc_hd__nand2_2 _27302_ (.A(_05245_),
    .B(_05223_),
    .Y(_05293_));
 sky130_fd_sc_hd__a21oi_2 _27303_ (.A1(_05289_),
    .A2(_05290_),
    .B1(_05285_),
    .Y(_05294_));
 sky130_fd_sc_hd__and3_2 _27304_ (.A(_05262_),
    .B(_05263_),
    .C(_05264_),
    .X(_05295_));
 sky130_fd_sc_hd__nand2_2 _27305_ (.A(_05278_),
    .B(_05259_),
    .Y(_05296_));
 sky130_fd_sc_hd__o211a_2 _27306_ (.A1(_05295_),
    .A2(_05296_),
    .B1(_05289_),
    .C1(_05285_),
    .X(_05297_));
 sky130_fd_sc_hd__nor3_2 _27307_ (.A(_05293_),
    .B(_05294_),
    .C(_05297_),
    .Y(_05298_));
 sky130_fd_sc_hd__o22ai_2 _27308_ (.A1(_05244_),
    .A2(_04840_),
    .B1(_05292_),
    .B2(_05298_),
    .Y(_05299_));
 sky130_fd_sc_hd__o21ai_2 _27309_ (.A1(_05294_),
    .A2(_05297_),
    .B1(_05293_),
    .Y(_05300_));
 sky130_fd_sc_hd__nand3b_2 _27310_ (.A_N(_05293_),
    .B(_05286_),
    .C(_05291_),
    .Y(_05301_));
 sky130_fd_sc_hd__nor2_2 _27311_ (.A(_05244_),
    .B(_04840_),
    .Y(_05302_));
 sky130_fd_sc_hd__nand3_2 _27312_ (.A(_05300_),
    .B(_05301_),
    .C(_05302_),
    .Y(_05303_));
 sky130_fd_sc_hd__nand2_2 _27313_ (.A(_05232_),
    .B(_05234_),
    .Y(_05304_));
 sky130_fd_sc_hd__nand2_2 _27314_ (.A(_05304_),
    .B(_05229_),
    .Y(_05305_));
 sky130_fd_sc_hd__a21oi_2 _27315_ (.A1(_05299_),
    .A2(_05303_),
    .B1(_05305_),
    .Y(_05306_));
 sky130_fd_sc_hd__nand2_2 _27316_ (.A(_05300_),
    .B(_05302_),
    .Y(_05307_));
 sky130_fd_sc_hd__o211a_2 _27317_ (.A1(_05298_),
    .A2(_05307_),
    .B1(_05305_),
    .C1(_05299_),
    .X(_05308_));
 sky130_fd_sc_hd__o22ai_2 _27318_ (.A1(_05240_),
    .A2(_05243_),
    .B1(_05306_),
    .B2(_05308_),
    .Y(_05309_));
 sky130_fd_sc_hd__a21o_2 _27319_ (.A1(_05299_),
    .A2(_05303_),
    .B1(_05305_),
    .X(_05310_));
 sky130_fd_sc_hd__a21o_2 _27320_ (.A1(_05241_),
    .A2(_05239_),
    .B1(_05242_),
    .X(_05311_));
 sky130_fd_sc_hd__nand3_2 _27321_ (.A(_05299_),
    .B(_05303_),
    .C(_05305_),
    .Y(_05312_));
 sky130_fd_sc_hd__nand3_2 _27322_ (.A(_05310_),
    .B(_05311_),
    .C(_05312_),
    .Y(_05313_));
 sky130_fd_sc_hd__nor2_2 _27323_ (.A(_05242_),
    .B(_05240_),
    .Y(_05314_));
 sky130_fd_sc_hd__nand3b_2 _27324_ (.A_N(_05140_),
    .B(_05314_),
    .C(_05175_),
    .Y(_05315_));
 sky130_fd_sc_hd__a21oi_2 _27325_ (.A1(_05309_),
    .A2(_05313_),
    .B1(_05315_),
    .Y(_05316_));
 sky130_fd_sc_hd__and3_2 _27326_ (.A(_05309_),
    .B(_05313_),
    .C(_05315_),
    .X(_05317_));
 sky130_fd_sc_hd__nor2_2 _27327_ (.A(_05316_),
    .B(_05317_),
    .Y(_02683_));
 sky130_fd_sc_hd__a22oi_2 _27328_ (.A1(_19388_),
    .A2(_05215_),
    .B1(_19391_),
    .B2(_19630_),
    .Y(_05318_));
 sky130_fd_sc_hd__inv_2 _27329_ (.A(_05146_),
    .Y(_05319_));
 sky130_fd_sc_hd__buf_1 _27330_ (.A(_05319_),
    .X(_05320_));
 sky130_fd_sc_hd__buf_1 _27331_ (.A(_19387_),
    .X(_05321_));
 sky130_fd_sc_hd__buf_1 _27332_ (.A(\pcpi_mul.rs2[4] ),
    .X(_05322_));
 sky130_fd_sc_hd__buf_1 _27333_ (.A(_19632_),
    .X(_05323_));
 sky130_fd_sc_hd__nand3_2 _27334_ (.A(_05321_),
    .B(_05322_),
    .C(_05323_),
    .Y(_05324_));
 sky130_fd_sc_hd__nor2_2 _27335_ (.A(_05320_),
    .B(_05324_),
    .Y(_05325_));
 sky130_fd_sc_hd__nand2_2 _27336_ (.A(_04834_),
    .B(_19618_),
    .Y(_05326_));
 sky130_fd_sc_hd__o21ai_2 _27337_ (.A1(_05318_),
    .A2(_05325_),
    .B1(_05326_),
    .Y(_05327_));
 sky130_fd_sc_hd__o22ai_2 _27338_ (.A1(_05101_),
    .A2(_05199_),
    .B1(_05252_),
    .B2(_05246_),
    .Y(_05328_));
 sky130_fd_sc_hd__inv_2 _27339_ (.A(_05326_),
    .Y(_05329_));
 sky130_fd_sc_hd__buf_1 _27340_ (.A(_19629_),
    .X(_05330_));
 sky130_fd_sc_hd__a22o_2 _27341_ (.A1(_19388_),
    .A2(_05215_),
    .B1(_19391_),
    .B2(_05330_),
    .X(_05331_));
 sky130_fd_sc_hd__o211ai_2 _27342_ (.A1(_05320_),
    .A2(_05324_),
    .B1(_05329_),
    .C1(_05331_),
    .Y(_05332_));
 sky130_fd_sc_hd__nand3_2 _27343_ (.A(_05327_),
    .B(_05328_),
    .C(_05332_),
    .Y(_05333_));
 sky130_fd_sc_hd__o21ai_2 _27344_ (.A1(_05318_),
    .A2(_05325_),
    .B1(_05329_),
    .Y(_05334_));
 sky130_fd_sc_hd__a21oi_2 _27345_ (.A1(_05253_),
    .A2(_05257_),
    .B1(_05250_),
    .Y(_05335_));
 sky130_fd_sc_hd__o211ai_2 _27346_ (.A1(_05320_),
    .A2(_05324_),
    .B1(_05326_),
    .C1(_05331_),
    .Y(_05336_));
 sky130_fd_sc_hd__nand3_2 _27347_ (.A(_05334_),
    .B(_05335_),
    .C(_05336_),
    .Y(_05337_));
 sky130_fd_sc_hd__buf_1 _27348_ (.A(_05211_),
    .X(_05338_));
 sky130_fd_sc_hd__nand2_2 _27349_ (.A(\pcpi_mul.rs2[3] ),
    .B(_05338_),
    .Y(_05339_));
 sky130_fd_sc_hd__buf_1 _27350_ (.A(_19624_),
    .X(_05340_));
 sky130_fd_sc_hd__buf_1 _27351_ (.A(_05340_),
    .X(_05341_));
 sky130_fd_sc_hd__buf_1 _27352_ (.A(\pcpi_mul.rs1[6] ),
    .X(_05342_));
 sky130_fd_sc_hd__buf_1 _27353_ (.A(_05342_),
    .X(_05343_));
 sky130_fd_sc_hd__a22oi_2 _27354_ (.A1(_05123_),
    .A2(_05341_),
    .B1(_05118_),
    .B2(_05343_),
    .Y(_05344_));
 sky130_fd_sc_hd__buf_1 _27355_ (.A(_19624_),
    .X(_05345_));
 sky130_fd_sc_hd__nand2_2 _27356_ (.A(_05122_),
    .B(_05345_),
    .Y(_05346_));
 sky130_fd_sc_hd__buf_1 _27357_ (.A(_19621_),
    .X(_05347_));
 sky130_fd_sc_hd__nand2_2 _27358_ (.A(_19400_),
    .B(_05347_),
    .Y(_05348_));
 sky130_fd_sc_hd__nor2_2 _27359_ (.A(_05346_),
    .B(_05348_),
    .Y(_05349_));
 sky130_fd_sc_hd__nor3_2 _27360_ (.A(_05339_),
    .B(_05344_),
    .C(_05349_),
    .Y(_05350_));
 sky130_fd_sc_hd__o21a_2 _27361_ (.A1(_05344_),
    .A2(_05349_),
    .B1(_05339_),
    .X(_05351_));
 sky130_fd_sc_hd__o2bb2ai_2 _27362_ (.A1_N(_05333_),
    .A2_N(_05337_),
    .B1(_05350_),
    .B2(_05351_),
    .Y(_05352_));
 sky130_fd_sc_hd__nand2_2 _27363_ (.A(_05346_),
    .B(_05348_),
    .Y(_05353_));
 sky130_fd_sc_hd__nand3b_2 _27364_ (.A_N(_05349_),
    .B(_05339_),
    .C(_05353_),
    .Y(_05354_));
 sky130_fd_sc_hd__inv_2 _27365_ (.A(_05339_),
    .Y(_05355_));
 sky130_fd_sc_hd__o21ai_2 _27366_ (.A1(_05344_),
    .A2(_05349_),
    .B1(_05355_),
    .Y(_05356_));
 sky130_fd_sc_hd__nand2_2 _27367_ (.A(_05354_),
    .B(_05356_),
    .Y(_05357_));
 sky130_fd_sc_hd__nand3_2 _27368_ (.A(_05357_),
    .B(_05337_),
    .C(_05333_),
    .Y(_05358_));
 sky130_fd_sc_hd__nand2_2 _27369_ (.A(_05296_),
    .B(_05265_),
    .Y(_05359_));
 sky130_fd_sc_hd__a21oi_2 _27370_ (.A1(_05352_),
    .A2(_05358_),
    .B1(_05359_),
    .Y(_05360_));
 sky130_fd_sc_hd__and3_2 _27371_ (.A(_05327_),
    .B(_05328_),
    .C(_05332_),
    .X(_05361_));
 sky130_fd_sc_hd__nand2_2 _27372_ (.A(_05357_),
    .B(_05337_),
    .Y(_05362_));
 sky130_fd_sc_hd__o211a_2 _27373_ (.A1(_05361_),
    .A2(_05362_),
    .B1(_05352_),
    .C1(_05359_),
    .X(_05363_));
 sky130_fd_sc_hd__nor2_2 _27374_ (.A(_05275_),
    .B(_05287_),
    .Y(_05364_));
 sky130_fd_sc_hd__o21ai_2 _27375_ (.A1(_05360_),
    .A2(_05363_),
    .B1(_05364_),
    .Y(_05365_));
 sky130_fd_sc_hd__a21o_2 _27376_ (.A1(_05352_),
    .A2(_05358_),
    .B1(_05359_),
    .X(_05366_));
 sky130_fd_sc_hd__nand3_2 _27377_ (.A(_05359_),
    .B(_05352_),
    .C(_05358_),
    .Y(_05367_));
 sky130_fd_sc_hd__inv_2 _27378_ (.A(_05364_),
    .Y(_05368_));
 sky130_fd_sc_hd__nand3_2 _27379_ (.A(_05366_),
    .B(_05367_),
    .C(_05368_),
    .Y(_05369_));
 sky130_fd_sc_hd__nand2_2 _27380_ (.A(_19384_),
    .B(_19641_),
    .Y(_05370_));
 sky130_fd_sc_hd__nand2_2 _27381_ (.A(_19386_),
    .B(_19637_),
    .Y(_05371_));
 sky130_fd_sc_hd__nor2_2 _27382_ (.A(_05370_),
    .B(_05371_),
    .Y(_05372_));
 sky130_fd_sc_hd__inv_2 _27383_ (.A(_05372_),
    .Y(_05373_));
 sky130_fd_sc_hd__nand2_2 _27384_ (.A(_05370_),
    .B(_05371_),
    .Y(_05374_));
 sky130_fd_sc_hd__nand2_2 _27385_ (.A(_05373_),
    .B(_05374_),
    .Y(_05375_));
 sky130_fd_sc_hd__inv_2 _27386_ (.A(_05375_),
    .Y(_05376_));
 sky130_fd_sc_hd__nand3_2 _27387_ (.A(_05365_),
    .B(_05369_),
    .C(_05376_),
    .Y(_05377_));
 sky130_fd_sc_hd__buf_1 _27388_ (.A(_05377_),
    .X(_05378_));
 sky130_fd_sc_hd__o21ai_2 _27389_ (.A1(_05360_),
    .A2(_05363_),
    .B1(_05368_),
    .Y(_05379_));
 sky130_fd_sc_hd__nand3_2 _27390_ (.A(_05366_),
    .B(_05367_),
    .C(_05364_),
    .Y(_05380_));
 sky130_fd_sc_hd__nand3_2 _27391_ (.A(_05379_),
    .B(_05375_),
    .C(_05380_),
    .Y(_05381_));
 sky130_fd_sc_hd__o2bb2ai_2 _27392_ (.A1_N(_05378_),
    .A2_N(_05381_),
    .B1(_05298_),
    .B2(_05307_),
    .Y(_05382_));
 sky130_fd_sc_hd__nand3b_2 _27393_ (.A_N(_05303_),
    .B(_05377_),
    .C(_05381_),
    .Y(_05383_));
 sky130_fd_sc_hd__nor2_2 _27394_ (.A(_05293_),
    .B(_05294_),
    .Y(_05384_));
 sky130_fd_sc_hd__nor2_2 _27395_ (.A(_05297_),
    .B(_05384_),
    .Y(_05385_));
 sky130_fd_sc_hd__inv_2 _27396_ (.A(_05385_),
    .Y(_05386_));
 sky130_fd_sc_hd__a21oi_2 _27397_ (.A1(_05382_),
    .A2(_05383_),
    .B1(_05386_),
    .Y(_05387_));
 sky130_fd_sc_hd__o211a_2 _27398_ (.A1(_05297_),
    .A2(_05384_),
    .B1(_05383_),
    .C1(_05382_),
    .X(_05388_));
 sky130_fd_sc_hd__nor2_2 _27399_ (.A(_05387_),
    .B(_05388_),
    .Y(_05389_));
 sky130_fd_sc_hd__a21oi_2 _27400_ (.A1(_05310_),
    .A2(_05240_),
    .B1(_05308_),
    .Y(_05390_));
 sky130_fd_sc_hd__and3_2 _27401_ (.A(_05310_),
    .B(_05312_),
    .C(_05243_),
    .X(_05391_));
 sky130_fd_sc_hd__a211oi_2 _27402_ (.A1(_05389_),
    .A2(_05390_),
    .B1(_05391_),
    .C1(_05316_),
    .Y(_05392_));
 sky130_fd_sc_hd__nor2_2 _27403_ (.A(_05239_),
    .B(_05306_),
    .Y(_05393_));
 sky130_fd_sc_hd__o22ai_2 _27404_ (.A1(_05308_),
    .A2(_05393_),
    .B1(_05387_),
    .B2(_05388_),
    .Y(_05394_));
 sky130_fd_sc_hd__nand2_2 _27405_ (.A(_05382_),
    .B(_05383_),
    .Y(_05395_));
 sky130_fd_sc_hd__nand2_2 _27406_ (.A(_05395_),
    .B(_05385_),
    .Y(_05396_));
 sky130_fd_sc_hd__nand3_2 _27407_ (.A(_05382_),
    .B(_05383_),
    .C(_05386_),
    .Y(_05397_));
 sky130_fd_sc_hd__nand3_2 _27408_ (.A(_05390_),
    .B(_05396_),
    .C(_05397_),
    .Y(_05398_));
 sky130_fd_sc_hd__o2bb2ai_2 _27409_ (.A1_N(_05398_),
    .A2_N(_05394_),
    .B1(_05391_),
    .B2(_05316_),
    .Y(_05399_));
 sky130_fd_sc_hd__a21boi_2 _27410_ (.A1(_05392_),
    .A2(_05394_),
    .B1_N(_05399_),
    .Y(_02684_));
 sky130_fd_sc_hd__buf_1 _27411_ (.A(_05388_),
    .X(_05400_));
 sky130_fd_sc_hd__nand2_2 _27412_ (.A(_05362_),
    .B(_05333_),
    .Y(_05401_));
 sky130_fd_sc_hd__buf_1 _27413_ (.A(_05180_),
    .X(_05402_));
 sky130_fd_sc_hd__buf_1 _27414_ (.A(_05189_),
    .X(_05403_));
 sky130_fd_sc_hd__a22oi_2 _27415_ (.A1(_05402_),
    .A2(_05204_),
    .B1(_05403_),
    .B2(_05207_),
    .Y(_05404_));
 sky130_fd_sc_hd__nand2_2 _27416_ (.A(_05189_),
    .B(_19627_),
    .Y(_05405_));
 sky130_fd_sc_hd__nand2_2 _27417_ (.A(_05187_),
    .B(_05218_),
    .Y(_05406_));
 sky130_fd_sc_hd__nor2_2 _27418_ (.A(_05405_),
    .B(_05406_),
    .Y(_05407_));
 sky130_fd_sc_hd__buf_1 _27419_ (.A(\pcpi_mul.rs1[8] ),
    .X(_05408_));
 sky130_fd_sc_hd__nand2_2 _27420_ (.A(_04834_),
    .B(_05408_),
    .Y(_05409_));
 sky130_fd_sc_hd__o21ai_2 _27421_ (.A1(_05404_),
    .A2(_05407_),
    .B1(_05409_),
    .Y(_05410_));
 sky130_fd_sc_hd__inv_2 _27422_ (.A(_05409_),
    .Y(_05411_));
 sky130_fd_sc_hd__nand2_2 _27423_ (.A(_05405_),
    .B(_05406_),
    .Y(_05412_));
 sky130_fd_sc_hd__nand3b_2 _27424_ (.A_N(_05407_),
    .B(_05411_),
    .C(_05412_),
    .Y(_05413_));
 sky130_fd_sc_hd__nor2_2 _27425_ (.A(_05329_),
    .B(_05325_),
    .Y(_05414_));
 sky130_fd_sc_hd__o2bb2ai_2 _27426_ (.A1_N(_05410_),
    .A2_N(_05413_),
    .B1(_05318_),
    .B2(_05414_),
    .Y(_05415_));
 sky130_fd_sc_hd__nor2_2 _27427_ (.A(_05326_),
    .B(_05318_),
    .Y(_05416_));
 sky130_fd_sc_hd__o211ai_2 _27428_ (.A1(_05325_),
    .A2(_05416_),
    .B1(_05410_),
    .C1(_05413_),
    .Y(_05417_));
 sky130_fd_sc_hd__nand2_2 _27429_ (.A(_05415_),
    .B(_05417_),
    .Y(_05418_));
 sky130_fd_sc_hd__buf_1 _27430_ (.A(\pcpi_mul.rs1[7] ),
    .X(_05419_));
 sky130_fd_sc_hd__buf_1 _27431_ (.A(_05419_),
    .X(_05420_));
 sky130_fd_sc_hd__buf_1 _27432_ (.A(_05420_),
    .X(_05421_));
 sky130_fd_sc_hd__buf_1 _27433_ (.A(_05251_),
    .X(_05422_));
 sky130_fd_sc_hd__nand2_2 _27434_ (.A(_05268_),
    .B(_05422_),
    .Y(_05423_));
 sky130_fd_sc_hd__a21o_2 _27435_ (.A1(_05205_),
    .A2(_05421_),
    .B1(_05423_),
    .X(_05424_));
 sky130_fd_sc_hd__buf_1 _27436_ (.A(_05251_),
    .X(_05425_));
 sky130_fd_sc_hd__buf_1 _27437_ (.A(_05419_),
    .X(_05426_));
 sky130_fd_sc_hd__nand2_2 _27438_ (.A(_05210_),
    .B(_05426_),
    .Y(_05427_));
 sky130_fd_sc_hd__a21o_2 _27439_ (.A1(_19398_),
    .A2(_05425_),
    .B1(_05427_),
    .X(_05428_));
 sky130_fd_sc_hd__nand2_2 _27440_ (.A(_05115_),
    .B(_19626_),
    .Y(_05429_));
 sky130_fd_sc_hd__a21oi_2 _27441_ (.A1(_05424_),
    .A2(_05428_),
    .B1(_05429_),
    .Y(_05430_));
 sky130_fd_sc_hd__and3_2 _27442_ (.A(_05424_),
    .B(_05428_),
    .C(_05429_),
    .X(_05431_));
 sky130_fd_sc_hd__nor2_2 _27443_ (.A(_05430_),
    .B(_05431_),
    .Y(_05432_));
 sky130_fd_sc_hd__nand2_2 _27444_ (.A(_05418_),
    .B(_05432_),
    .Y(_05433_));
 sky130_fd_sc_hd__nand3_2 _27445_ (.A(_05424_),
    .B(_05428_),
    .C(_05429_),
    .Y(_05434_));
 sky130_fd_sc_hd__or2b_2 _27446_ (.A(_05430_),
    .B_N(_05434_),
    .X(_05435_));
 sky130_fd_sc_hd__nand3_2 _27447_ (.A(_05435_),
    .B(_05415_),
    .C(_05417_),
    .Y(_05436_));
 sky130_fd_sc_hd__nand3b_2 _27448_ (.A_N(_05401_),
    .B(_05433_),
    .C(_05436_),
    .Y(_05437_));
 sky130_fd_sc_hd__nand2_2 _27449_ (.A(_05418_),
    .B(_05435_),
    .Y(_05438_));
 sky130_fd_sc_hd__nand3_2 _27450_ (.A(_05432_),
    .B(_05415_),
    .C(_05417_),
    .Y(_05439_));
 sky130_fd_sc_hd__nand3_2 _27451_ (.A(_05438_),
    .B(_05401_),
    .C(_05439_),
    .Y(_05440_));
 sky130_fd_sc_hd__nand2_2 _27452_ (.A(_05437_),
    .B(_05440_),
    .Y(_05441_));
 sky130_fd_sc_hd__a21oi_2 _27453_ (.A1(_05355_),
    .A2(_05353_),
    .B1(_05349_),
    .Y(_05442_));
 sky130_fd_sc_hd__nand2_2 _27454_ (.A(_05441_),
    .B(_05442_),
    .Y(_05443_));
 sky130_fd_sc_hd__nand3b_2 _27455_ (.A_N(_05442_),
    .B(_05437_),
    .C(_05440_),
    .Y(_05444_));
 sky130_fd_sc_hd__buf_1 _27456_ (.A(_19382_),
    .X(_05445_));
 sky130_fd_sc_hd__nand2_2 _27457_ (.A(_05445_),
    .B(_05190_),
    .Y(_05446_));
 sky130_fd_sc_hd__buf_1 _27458_ (.A(\pcpi_mul.rs2[8] ),
    .X(_05447_));
 sky130_fd_sc_hd__buf_1 _27459_ (.A(_05447_),
    .X(_05448_));
 sky130_fd_sc_hd__nand2_2 _27460_ (.A(_05448_),
    .B(_05188_),
    .Y(_05449_));
 sky130_fd_sc_hd__nor2_2 _27461_ (.A(_05446_),
    .B(_05449_),
    .Y(_05450_));
 sky130_fd_sc_hd__nand2_2 _27462_ (.A(_05446_),
    .B(_05449_),
    .Y(_05451_));
 sky130_fd_sc_hd__inv_2 _27463_ (.A(_05451_),
    .Y(_05452_));
 sky130_fd_sc_hd__nand2_2 _27464_ (.A(_19386_),
    .B(_05120_),
    .Y(_05453_));
 sky130_fd_sc_hd__o21bai_2 _27465_ (.A1(_05450_),
    .A2(_05452_),
    .B1_N(_05453_),
    .Y(_05454_));
 sky130_fd_sc_hd__inv_2 _27466_ (.A(_05450_),
    .Y(_05455_));
 sky130_fd_sc_hd__nand3_2 _27467_ (.A(_05455_),
    .B(_05453_),
    .C(_05451_),
    .Y(_05456_));
 sky130_fd_sc_hd__nand2_2 _27468_ (.A(_05454_),
    .B(_05456_),
    .Y(_05457_));
 sky130_fd_sc_hd__or2_2 _27469_ (.A(_05372_),
    .B(_05457_),
    .X(_05458_));
 sky130_fd_sc_hd__nand2_2 _27470_ (.A(_05457_),
    .B(_05372_),
    .Y(_05459_));
 sky130_fd_sc_hd__nand2_2 _27471_ (.A(_05458_),
    .B(_05459_),
    .Y(_05460_));
 sky130_fd_sc_hd__inv_2 _27472_ (.A(_05460_),
    .Y(_05461_));
 sky130_fd_sc_hd__a21oi_2 _27473_ (.A1(_05443_),
    .A2(_05444_),
    .B1(_05461_),
    .Y(_05462_));
 sky130_fd_sc_hd__and3_2 _27474_ (.A(_05443_),
    .B(_05444_),
    .C(_05461_),
    .X(_05463_));
 sky130_fd_sc_hd__o21ai_2 _27475_ (.A1(_05462_),
    .A2(_05463_),
    .B1(_05378_),
    .Y(_05464_));
 sky130_fd_sc_hd__a21o_2 _27476_ (.A1(_05443_),
    .A2(_05444_),
    .B1(_05461_),
    .X(_05465_));
 sky130_fd_sc_hd__inv_2 _27477_ (.A(_05377_),
    .Y(_05466_));
 sky130_fd_sc_hd__a21oi_2 _27478_ (.A1(_05441_),
    .A2(_05442_),
    .B1(_05460_),
    .Y(_05467_));
 sky130_fd_sc_hd__nand2_2 _27479_ (.A(_05467_),
    .B(_05444_),
    .Y(_05468_));
 sky130_fd_sc_hd__nand3_2 _27480_ (.A(_05465_),
    .B(_05466_),
    .C(_05468_),
    .Y(_05469_));
 sky130_fd_sc_hd__nand2_2 _27481_ (.A(_05464_),
    .B(_05469_),
    .Y(_05470_));
 sky130_fd_sc_hd__nor2_2 _27482_ (.A(_05364_),
    .B(_05360_),
    .Y(_05471_));
 sky130_fd_sc_hd__nand3b_2 _27483_ (.A_N(_05471_),
    .B(_05383_),
    .C(_05367_),
    .Y(_05472_));
 sky130_fd_sc_hd__inv_2 _27484_ (.A(_05303_),
    .Y(_05473_));
 sky130_fd_sc_hd__o2111ai_2 _27485_ (.A1(_05363_),
    .A2(_05471_),
    .B1(_05378_),
    .C1(_05381_),
    .D1(_05473_),
    .Y(_05474_));
 sky130_fd_sc_hd__nand2_2 _27486_ (.A(_05472_),
    .B(_05474_),
    .Y(_05475_));
 sky130_fd_sc_hd__nand2_2 _27487_ (.A(_05470_),
    .B(_05475_),
    .Y(_05476_));
 sky130_fd_sc_hd__nand2_2 _27488_ (.A(_05465_),
    .B(_05466_),
    .Y(_05477_));
 sky130_fd_sc_hd__o2111ai_2 _27489_ (.A1(_05463_),
    .A2(_05477_),
    .B1(_05474_),
    .C1(_05464_),
    .D1(_05472_),
    .Y(_05478_));
 sky130_fd_sc_hd__nand2_2 _27490_ (.A(_05396_),
    .B(_05308_),
    .Y(_05479_));
 sky130_fd_sc_hd__nand3_2 _27491_ (.A(_05476_),
    .B(_05478_),
    .C(_05479_),
    .Y(_05480_));
 sky130_fd_sc_hd__a21oi_2 _27492_ (.A1(_05395_),
    .A2(_05385_),
    .B1(_05312_),
    .Y(_05481_));
 sky130_fd_sc_hd__nand3_2 _27493_ (.A(_05475_),
    .B(_05464_),
    .C(_05469_),
    .Y(_05482_));
 sky130_fd_sc_hd__nand3_2 _27494_ (.A(_05470_),
    .B(_05474_),
    .C(_05472_),
    .Y(_05483_));
 sky130_fd_sc_hd__o211ai_2 _27495_ (.A1(_05400_),
    .A2(_05481_),
    .B1(_05482_),
    .C1(_05483_),
    .Y(_05484_));
 sky130_fd_sc_hd__o21ai_2 _27496_ (.A1(_05400_),
    .A2(_05480_),
    .B1(_05484_),
    .Y(_05485_));
 sky130_fd_sc_hd__nand3_2 _27497_ (.A(_05389_),
    .B(_05312_),
    .C(_05393_),
    .Y(_05486_));
 sky130_fd_sc_hd__nand2_2 _27498_ (.A(_05399_),
    .B(_05486_),
    .Y(_05487_));
 sky130_fd_sc_hd__xor2_2 _27499_ (.A(_05485_),
    .B(_05487_),
    .X(_02685_));
 sky130_fd_sc_hd__nand2_2 _27500_ (.A(_05483_),
    .B(_05482_),
    .Y(_05488_));
 sky130_fd_sc_hd__nor2_2 _27501_ (.A(_05400_),
    .B(_05479_),
    .Y(_05489_));
 sky130_fd_sc_hd__a22oi_2 _27502_ (.A1(_05488_),
    .A2(_05489_),
    .B1(_05487_),
    .B2(_05485_),
    .Y(_05490_));
 sky130_fd_sc_hd__nand2_2 _27503_ (.A(_05444_),
    .B(_05440_),
    .Y(_05491_));
 sky130_fd_sc_hd__inv_2 _27504_ (.A(_05491_),
    .Y(_05492_));
 sky130_fd_sc_hd__nand2_2 _27505_ (.A(_05469_),
    .B(_05492_),
    .Y(_05493_));
 sky130_fd_sc_hd__nor2_2 _27506_ (.A(_05378_),
    .B(_05492_),
    .Y(_05494_));
 sky130_fd_sc_hd__nand3_2 _27507_ (.A(_05494_),
    .B(_05468_),
    .C(_05465_),
    .Y(_05495_));
 sky130_fd_sc_hd__inv_2 _27508_ (.A(\pcpi_mul.rs2[9] ),
    .Y(_05496_));
 sky130_fd_sc_hd__buf_1 _27509_ (.A(_05496_),
    .X(_05497_));
 sky130_fd_sc_hd__buf_1 _27510_ (.A(_05497_),
    .X(_05498_));
 sky130_fd_sc_hd__nand2_2 _27511_ (.A(_05432_),
    .B(_05415_),
    .Y(_05499_));
 sky130_fd_sc_hd__nand2_2 _27512_ (.A(_05499_),
    .B(_05417_),
    .Y(_05500_));
 sky130_fd_sc_hd__buf_1 _27513_ (.A(_05260_),
    .X(_05501_));
 sky130_fd_sc_hd__buf_1 _27514_ (.A(\pcpi_mul.rs1[7] ),
    .X(_05502_));
 sky130_fd_sc_hd__nand2_2 _27515_ (.A(_05122_),
    .B(_05502_),
    .Y(_05503_));
 sky130_fd_sc_hd__a21o_2 _27516_ (.A1(_05221_),
    .A2(_19616_),
    .B1(_05503_),
    .X(_05504_));
 sky130_fd_sc_hd__buf_1 _27517_ (.A(_19618_),
    .X(_05505_));
 sky130_fd_sc_hd__buf_1 _27518_ (.A(\pcpi_mul.rs1[8] ),
    .X(_05506_));
 sky130_fd_sc_hd__nand2_2 _27519_ (.A(_19400_),
    .B(_05506_),
    .Y(_05507_));
 sky130_fd_sc_hd__a21o_2 _27520_ (.A1(_05203_),
    .A2(_05505_),
    .B1(_05507_),
    .X(_05508_));
 sky130_fd_sc_hd__o211a_2 _27521_ (.A1(_05149_),
    .A2(_05501_),
    .B1(_05504_),
    .C1(_05508_),
    .X(_05509_));
 sky130_fd_sc_hd__nand2_2 _27522_ (.A(_05115_),
    .B(_19623_),
    .Y(_05510_));
 sky130_fd_sc_hd__a21oi_2 _27523_ (.A1(_05504_),
    .A2(_05508_),
    .B1(_05510_),
    .Y(_05511_));
 sky130_fd_sc_hd__nand2_2 _27524_ (.A(_05321_),
    .B(_05206_),
    .Y(_05512_));
 sky130_fd_sc_hd__nand2_2 _27525_ (.A(_05322_),
    .B(_05184_),
    .Y(_05513_));
 sky130_fd_sc_hd__nor2_2 _27526_ (.A(_05512_),
    .B(_05513_),
    .Y(_05514_));
 sky130_fd_sc_hd__and2_2 _27527_ (.A(_05512_),
    .B(_05513_),
    .X(_05515_));
 sky130_fd_sc_hd__buf_1 _27528_ (.A(\pcpi_mul.rs1[9] ),
    .X(_05516_));
 sky130_fd_sc_hd__nand2_2 _27529_ (.A(_05157_),
    .B(_05516_),
    .Y(_05517_));
 sky130_fd_sc_hd__o21ai_2 _27530_ (.A1(_05514_),
    .A2(_05515_),
    .B1(_05517_),
    .Y(_05518_));
 sky130_fd_sc_hd__or2_2 _27531_ (.A(_05512_),
    .B(_05513_),
    .X(_05519_));
 sky130_fd_sc_hd__inv_2 _27532_ (.A(_05517_),
    .Y(_05520_));
 sky130_fd_sc_hd__nand2_2 _27533_ (.A(_05512_),
    .B(_05513_),
    .Y(_05521_));
 sky130_fd_sc_hd__nand3_2 _27534_ (.A(_05519_),
    .B(_05520_),
    .C(_05521_),
    .Y(_05522_));
 sky130_fd_sc_hd__a21o_2 _27535_ (.A1(_05411_),
    .A2(_05412_),
    .B1(_05407_),
    .X(_05523_));
 sky130_fd_sc_hd__nand3_2 _27536_ (.A(_05518_),
    .B(_05522_),
    .C(_05523_),
    .Y(_05524_));
 sky130_fd_sc_hd__o21ai_2 _27537_ (.A1(_05514_),
    .A2(_05515_),
    .B1(_05520_),
    .Y(_05525_));
 sky130_fd_sc_hd__nand3_2 _27538_ (.A(_05519_),
    .B(_05517_),
    .C(_05521_),
    .Y(_05526_));
 sky130_fd_sc_hd__a21oi_2 _27539_ (.A1(_05411_),
    .A2(_05412_),
    .B1(_05407_),
    .Y(_05527_));
 sky130_fd_sc_hd__nand3_2 _27540_ (.A(_05525_),
    .B(_05526_),
    .C(_05527_),
    .Y(_05528_));
 sky130_fd_sc_hd__nand2_2 _27541_ (.A(_05524_),
    .B(_05528_),
    .Y(_05529_));
 sky130_fd_sc_hd__o21ai_2 _27542_ (.A1(_05509_),
    .A2(_05511_),
    .B1(_05529_),
    .Y(_05530_));
 sky130_fd_sc_hd__nor2_2 _27543_ (.A(_05511_),
    .B(_05509_),
    .Y(_05531_));
 sky130_fd_sc_hd__nand3_2 _27544_ (.A(_05531_),
    .B(_05524_),
    .C(_05528_),
    .Y(_05532_));
 sky130_fd_sc_hd__nand3_2 _27545_ (.A(_05500_),
    .B(_05530_),
    .C(_05532_),
    .Y(_05533_));
 sky130_fd_sc_hd__a21boi_2 _27546_ (.A1(_05432_),
    .A2(_05415_),
    .B1_N(_05417_),
    .Y(_05534_));
 sky130_fd_sc_hd__nand3b_2 _27547_ (.A_N(_05531_),
    .B(_05524_),
    .C(_05528_),
    .Y(_05535_));
 sky130_fd_sc_hd__nand2_2 _27548_ (.A(_05529_),
    .B(_05531_),
    .Y(_05536_));
 sky130_fd_sc_hd__nand3_2 _27549_ (.A(_05534_),
    .B(_05535_),
    .C(_05536_),
    .Y(_05537_));
 sky130_fd_sc_hd__nand2_2 _27550_ (.A(_05533_),
    .B(_05537_),
    .Y(_05538_));
 sky130_fd_sc_hd__nor2_2 _27551_ (.A(_05423_),
    .B(_05427_),
    .Y(_05539_));
 sky130_fd_sc_hd__nor2_2 _27552_ (.A(_05539_),
    .B(_05430_),
    .Y(_05540_));
 sky130_fd_sc_hd__nand2_2 _27553_ (.A(_05538_),
    .B(_05540_),
    .Y(_05541_));
 sky130_fd_sc_hd__buf_1 _27554_ (.A(_05447_),
    .X(_05542_));
 sky130_fd_sc_hd__buf_1 _27555_ (.A(_05104_),
    .X(_05543_));
 sky130_fd_sc_hd__nand2_2 _27556_ (.A(_05542_),
    .B(_05543_),
    .Y(_05544_));
 sky130_fd_sc_hd__buf_1 _27557_ (.A(_19632_),
    .X(_05545_));
 sky130_fd_sc_hd__nand2_2 _27558_ (.A(_19383_),
    .B(_05545_),
    .Y(_05546_));
 sky130_fd_sc_hd__nor2_2 _27559_ (.A(_05544_),
    .B(_05546_),
    .Y(_05547_));
 sky130_fd_sc_hd__and2_2 _27560_ (.A(_05544_),
    .B(_05546_),
    .X(_05548_));
 sky130_fd_sc_hd__nand2_2 _27561_ (.A(_19385_),
    .B(_05218_),
    .Y(_05549_));
 sky130_fd_sc_hd__inv_2 _27562_ (.A(_05549_),
    .Y(_05550_));
 sky130_fd_sc_hd__o21ai_2 _27563_ (.A1(_05547_),
    .A2(_05548_),
    .B1(_05550_),
    .Y(_05551_));
 sky130_fd_sc_hd__nand2_2 _27564_ (.A(_05544_),
    .B(_05546_),
    .Y(_05552_));
 sky130_fd_sc_hd__nand3b_2 _27565_ (.A_N(_05547_),
    .B(_05549_),
    .C(_05552_),
    .Y(_05553_));
 sky130_fd_sc_hd__nor2_2 _27566_ (.A(_05453_),
    .B(_05452_),
    .Y(_05554_));
 sky130_fd_sc_hd__o2bb2ai_2 _27567_ (.A1_N(_05551_),
    .A2_N(_05553_),
    .B1(_05450_),
    .B2(_05554_),
    .Y(_05555_));
 sky130_fd_sc_hd__o2111ai_2 _27568_ (.A1(_05453_),
    .A2(_05452_),
    .B1(_05455_),
    .C1(_05553_),
    .D1(_05551_),
    .Y(_05556_));
 sky130_fd_sc_hd__nand2_2 _27569_ (.A(_05555_),
    .B(_05556_),
    .Y(_05557_));
 sky130_fd_sc_hd__nor2_2 _27570_ (.A(_05459_),
    .B(_05557_),
    .Y(_05558_));
 sky130_fd_sc_hd__nand2_2 _27571_ (.A(_05557_),
    .B(_05459_),
    .Y(_05559_));
 sky130_fd_sc_hd__and2b_2 _27572_ (.A_N(_05558_),
    .B(_05559_),
    .X(_05560_));
 sky130_fd_sc_hd__inv_2 _27573_ (.A(_05540_),
    .Y(_05561_));
 sky130_fd_sc_hd__nand3_2 _27574_ (.A(_05533_),
    .B(_05537_),
    .C(_05561_),
    .Y(_05562_));
 sky130_fd_sc_hd__nand3_2 _27575_ (.A(_05541_),
    .B(_05560_),
    .C(_05562_),
    .Y(_05563_));
 sky130_fd_sc_hd__o2bb2ai_2 _27576_ (.A1_N(_05533_),
    .A2_N(_05537_),
    .B1(_05539_),
    .B2(_05430_),
    .Y(_05564_));
 sky130_fd_sc_hd__or2_2 _27577_ (.A(_05459_),
    .B(_05557_),
    .X(_05565_));
 sky130_fd_sc_hd__nand2_2 _27578_ (.A(_05565_),
    .B(_05559_),
    .Y(_05566_));
 sky130_fd_sc_hd__nand3_2 _27579_ (.A(_05533_),
    .B(_05537_),
    .C(_05540_),
    .Y(_05567_));
 sky130_fd_sc_hd__nand3_2 _27580_ (.A(_05564_),
    .B(_05566_),
    .C(_05567_),
    .Y(_05568_));
 sky130_fd_sc_hd__a22oi_2 _27581_ (.A1(_05467_),
    .A2(_05444_),
    .B1(_05563_),
    .B2(_05568_),
    .Y(_05569_));
 sky130_fd_sc_hd__o2111a_2 _27582_ (.A1(_05442_),
    .A2(_05441_),
    .B1(_05467_),
    .C1(_05568_),
    .D1(_05563_),
    .X(_05570_));
 sky130_fd_sc_hd__o22ai_2 _27583_ (.A1(_05498_),
    .A2(_04840_),
    .B1(_05569_),
    .B2(_05570_),
    .Y(_05571_));
 sky130_fd_sc_hd__nand3_2 _27584_ (.A(_05463_),
    .B(_05563_),
    .C(_05568_),
    .Y(_05572_));
 sky130_fd_sc_hd__nand2_2 _27585_ (.A(_05563_),
    .B(_05568_),
    .Y(_05573_));
 sky130_fd_sc_hd__nand2_2 _27586_ (.A(_05573_),
    .B(_05468_),
    .Y(_05574_));
 sky130_fd_sc_hd__nor2_2 _27587_ (.A(_05498_),
    .B(_04840_),
    .Y(_05575_));
 sky130_fd_sc_hd__nand3_2 _27588_ (.A(_05572_),
    .B(_05574_),
    .C(_05575_),
    .Y(_05576_));
 sky130_fd_sc_hd__a22oi_2 _27589_ (.A1(_05493_),
    .A2(_05495_),
    .B1(_05571_),
    .B2(_05576_),
    .Y(_05577_));
 sky130_fd_sc_hd__nand3_2 _27590_ (.A(_05465_),
    .B(_05468_),
    .C(_05491_),
    .Y(_05578_));
 sky130_fd_sc_hd__o2111a_2 _27591_ (.A1(_05378_),
    .A2(_05578_),
    .B1(_05576_),
    .C1(_05493_),
    .D1(_05571_),
    .X(_05579_));
 sky130_fd_sc_hd__inv_2 _27592_ (.A(_05474_),
    .Y(_05580_));
 sky130_fd_sc_hd__a31o_2 _27593_ (.A1(_05464_),
    .A2(_05469_),
    .A3(_05472_),
    .B1(_05580_),
    .X(_05581_));
 sky130_fd_sc_hd__inv_2 _27594_ (.A(_05581_),
    .Y(_05582_));
 sky130_fd_sc_hd__o21ai_2 _27595_ (.A1(_05577_),
    .A2(_05579_),
    .B1(_05582_),
    .Y(_05583_));
 sky130_fd_sc_hd__a22o_2 _27596_ (.A1(_05495_),
    .A2(_05493_),
    .B1(_05571_),
    .B2(_05576_),
    .X(_05584_));
 sky130_fd_sc_hd__o2111ai_2 _27597_ (.A1(_05378_),
    .A2(_05578_),
    .B1(_05493_),
    .C1(_05576_),
    .D1(_05571_),
    .Y(_05585_));
 sky130_fd_sc_hd__nand3_2 _27598_ (.A(_05584_),
    .B(_05585_),
    .C(_05581_),
    .Y(_05586_));
 sky130_fd_sc_hd__a22oi_2 _27599_ (.A1(_05400_),
    .A2(_05488_),
    .B1(_05583_),
    .B2(_05586_),
    .Y(_05587_));
 sky130_fd_sc_hd__a31o_2 _27600_ (.A1(_05400_),
    .A2(_05488_),
    .A3(_05583_),
    .B1(_05587_),
    .X(_05588_));
 sky130_fd_sc_hd__xor2_2 _27601_ (.A(_05490_),
    .B(_05588_),
    .X(_02686_));
 sky130_fd_sc_hd__nand2_2 _27602_ (.A(_05488_),
    .B(_05400_),
    .Y(_05589_));
 sky130_fd_sc_hd__inv_2 _27603_ (.A(_05583_),
    .Y(_05590_));
 sky130_fd_sc_hd__o22ai_2 _27604_ (.A1(_05589_),
    .A2(_05590_),
    .B1(_05587_),
    .B2(_05490_),
    .Y(_05591_));
 sky130_fd_sc_hd__nand2_2 _27605_ (.A(_05531_),
    .B(_05528_),
    .Y(_05592_));
 sky130_fd_sc_hd__nand2_2 _27606_ (.A(_05592_),
    .B(_05524_),
    .Y(_05593_));
 sky130_fd_sc_hd__nand2_2 _27607_ (.A(_05321_),
    .B(_05340_),
    .Y(_05594_));
 sky130_fd_sc_hd__nand2_2 _27608_ (.A(_05155_),
    .B(_05342_),
    .Y(_05595_));
 sky130_fd_sc_hd__nor2_2 _27609_ (.A(_05594_),
    .B(_05595_),
    .Y(_05596_));
 sky130_fd_sc_hd__buf_1 _27610_ (.A(\pcpi_mul.rs1[10] ),
    .X(_05597_));
 sky130_fd_sc_hd__buf_1 _27611_ (.A(_05597_),
    .X(_05598_));
 sky130_fd_sc_hd__nand2_2 _27612_ (.A(_04834_),
    .B(_05598_),
    .Y(_05599_));
 sky130_fd_sc_hd__inv_2 _27613_ (.A(_05599_),
    .Y(_05600_));
 sky130_fd_sc_hd__nand2_2 _27614_ (.A(_05594_),
    .B(_05595_),
    .Y(_05601_));
 sky130_fd_sc_hd__nand2_2 _27615_ (.A(_05600_),
    .B(_05601_),
    .Y(_05602_));
 sky130_fd_sc_hd__a21o_2 _27616_ (.A1(_05520_),
    .A2(_05521_),
    .B1(_05514_),
    .X(_05603_));
 sky130_fd_sc_hd__and2_2 _27617_ (.A(_05594_),
    .B(_05595_),
    .X(_05604_));
 sky130_fd_sc_hd__o21ai_2 _27618_ (.A1(_05596_),
    .A2(_05604_),
    .B1(_05599_),
    .Y(_05605_));
 sky130_fd_sc_hd__o211ai_2 _27619_ (.A1(_05596_),
    .A2(_05602_),
    .B1(_05603_),
    .C1(_05605_),
    .Y(_05606_));
 sky130_fd_sc_hd__o21ai_2 _27620_ (.A1(_05596_),
    .A2(_05604_),
    .B1(_05600_),
    .Y(_05607_));
 sky130_fd_sc_hd__or2_2 _27621_ (.A(_05594_),
    .B(_05595_),
    .X(_05608_));
 sky130_fd_sc_hd__nand3_2 _27622_ (.A(_05608_),
    .B(_05599_),
    .C(_05601_),
    .Y(_05609_));
 sky130_fd_sc_hd__a21oi_2 _27623_ (.A1(_05520_),
    .A2(_05521_),
    .B1(_05514_),
    .Y(_05610_));
 sky130_fd_sc_hd__nand3_2 _27624_ (.A(_05607_),
    .B(_05609_),
    .C(_05610_),
    .Y(_05611_));
 sky130_fd_sc_hd__nand2_2 _27625_ (.A(_05606_),
    .B(_05611_),
    .Y(_05612_));
 sky130_fd_sc_hd__buf_1 _27626_ (.A(_19615_),
    .X(_05613_));
 sky130_fd_sc_hd__buf_1 _27627_ (.A(\pcpi_mul.rs1[9] ),
    .X(_05614_));
 sky130_fd_sc_hd__buf_1 _27628_ (.A(_05614_),
    .X(_05615_));
 sky130_fd_sc_hd__a22oi_2 _27629_ (.A1(_05203_),
    .A2(_05613_),
    .B1(_05143_),
    .B2(_05615_),
    .Y(_05616_));
 sky130_fd_sc_hd__nand2_2 _27630_ (.A(_19613_),
    .B(_05408_),
    .Y(_05617_));
 sky130_fd_sc_hd__nor2_2 _27631_ (.A(_05102_),
    .B(_05617_),
    .Y(_05618_));
 sky130_fd_sc_hd__nor2_2 _27632_ (.A(_05616_),
    .B(_05618_),
    .Y(_05619_));
 sky130_fd_sc_hd__nand2_2 _27633_ (.A(_19393_),
    .B(_05505_),
    .Y(_05620_));
 sky130_fd_sc_hd__nand2_2 _27634_ (.A(_05619_),
    .B(_05620_),
    .Y(_05621_));
 sky130_fd_sc_hd__inv_2 _27635_ (.A(_05620_),
    .Y(_05622_));
 sky130_fd_sc_hd__o21ai_2 _27636_ (.A1(_05616_),
    .A2(_05618_),
    .B1(_05622_),
    .Y(_05623_));
 sky130_fd_sc_hd__and2_2 _27637_ (.A(_05621_),
    .B(_05623_),
    .X(_05624_));
 sky130_fd_sc_hd__nand2_2 _27638_ (.A(_05612_),
    .B(_05624_),
    .Y(_05625_));
 sky130_fd_sc_hd__nand2_2 _27639_ (.A(_05621_),
    .B(_05623_),
    .Y(_05626_));
 sky130_fd_sc_hd__nand3_2 _27640_ (.A(_05606_),
    .B(_05611_),
    .C(_05626_),
    .Y(_05627_));
 sky130_fd_sc_hd__nand3_2 _27641_ (.A(_05593_),
    .B(_05625_),
    .C(_05627_),
    .Y(_05628_));
 sky130_fd_sc_hd__nand2_2 _27642_ (.A(_05612_),
    .B(_05626_),
    .Y(_05629_));
 sky130_fd_sc_hd__a21boi_2 _27643_ (.A1(_05531_),
    .A2(_05528_),
    .B1_N(_05524_),
    .Y(_05630_));
 sky130_fd_sc_hd__nand3_2 _27644_ (.A(_05624_),
    .B(_05606_),
    .C(_05611_),
    .Y(_05631_));
 sky130_fd_sc_hd__nand3_2 _27645_ (.A(_05629_),
    .B(_05630_),
    .C(_05631_),
    .Y(_05632_));
 sky130_fd_sc_hd__o21bai_2 _27646_ (.A1(_05503_),
    .A2(_05507_),
    .B1_N(_05511_),
    .Y(_05633_));
 sky130_fd_sc_hd__a21o_2 _27647_ (.A1(_05628_),
    .A2(_05632_),
    .B1(_05633_),
    .X(_05634_));
 sky130_fd_sc_hd__nand3_2 _27648_ (.A(_05628_),
    .B(_05632_),
    .C(_05633_),
    .Y(_05635_));
 sky130_fd_sc_hd__nand3_2 _27649_ (.A(_05556_),
    .B(_05457_),
    .C(_05372_),
    .Y(_05636_));
 sky130_fd_sc_hd__nand2_2 _27650_ (.A(_05636_),
    .B(_05555_),
    .Y(_05637_));
 sky130_fd_sc_hd__nand2_2 _27651_ (.A(_19386_),
    .B(_19628_),
    .Y(_05638_));
 sky130_fd_sc_hd__buf_1 _27652_ (.A(\pcpi_mul.rs2[8] ),
    .X(_05639_));
 sky130_fd_sc_hd__nand2_2 _27653_ (.A(_05639_),
    .B(_05323_),
    .Y(_05640_));
 sky130_fd_sc_hd__buf_1 _27654_ (.A(\pcpi_mul.rs2[7] ),
    .X(_05641_));
 sky130_fd_sc_hd__nand2_2 _27655_ (.A(_05641_),
    .B(_05271_),
    .Y(_05642_));
 sky130_fd_sc_hd__nor2_2 _27656_ (.A(_05640_),
    .B(_05642_),
    .Y(_05643_));
 sky130_fd_sc_hd__inv_2 _27657_ (.A(_05643_),
    .Y(_05644_));
 sky130_fd_sc_hd__nand2_2 _27658_ (.A(_05640_),
    .B(_05642_),
    .Y(_05645_));
 sky130_fd_sc_hd__nand3b_2 _27659_ (.A_N(_05638_),
    .B(_05644_),
    .C(_05645_),
    .Y(_05646_));
 sky130_fd_sc_hd__inv_2 _27660_ (.A(_05645_),
    .Y(_05647_));
 sky130_fd_sc_hd__o21ai_2 _27661_ (.A1(_05643_),
    .A2(_05647_),
    .B1(_05638_),
    .Y(_05648_));
 sky130_fd_sc_hd__nand2_2 _27662_ (.A(_05646_),
    .B(_05648_),
    .Y(_05649_));
 sky130_fd_sc_hd__a21o_2 _27663_ (.A1(_05550_),
    .A2(_05552_),
    .B1(_05547_),
    .X(_05650_));
 sky130_fd_sc_hd__inv_2 _27664_ (.A(_05650_),
    .Y(_05651_));
 sky130_fd_sc_hd__nand2_2 _27665_ (.A(_05649_),
    .B(_05651_),
    .Y(_05652_));
 sky130_fd_sc_hd__nand3_2 _27666_ (.A(_05646_),
    .B(_05648_),
    .C(_05650_),
    .Y(_05653_));
 sky130_fd_sc_hd__nand2_2 _27667_ (.A(_05652_),
    .B(_05653_),
    .Y(_05654_));
 sky130_fd_sc_hd__nand2_2 _27668_ (.A(_05637_),
    .B(_05654_),
    .Y(_05655_));
 sky130_fd_sc_hd__nor2_2 _27669_ (.A(_05450_),
    .B(_05554_),
    .Y(_05656_));
 sky130_fd_sc_hd__and2_2 _27670_ (.A(_05551_),
    .B(_05553_),
    .X(_05657_));
 sky130_fd_sc_hd__o2111ai_2 _27671_ (.A1(_05656_),
    .A2(_05657_),
    .B1(_05653_),
    .C1(_05652_),
    .D1(_05636_),
    .Y(_05658_));
 sky130_fd_sc_hd__nand2_2 _27672_ (.A(_05655_),
    .B(_05658_),
    .Y(_05659_));
 sky130_fd_sc_hd__a21o_2 _27673_ (.A1(_05634_),
    .A2(_05635_),
    .B1(_05659_),
    .X(_05660_));
 sky130_fd_sc_hd__a21oi_2 _27674_ (.A1(_05564_),
    .A2(_05567_),
    .B1(_05566_),
    .Y(_05661_));
 sky130_fd_sc_hd__nand3_2 _27675_ (.A(_05634_),
    .B(_05635_),
    .C(_05659_),
    .Y(_05662_));
 sky130_fd_sc_hd__nand3_2 _27676_ (.A(_05660_),
    .B(_05661_),
    .C(_05662_),
    .Y(_05663_));
 sky130_fd_sc_hd__buf_1 _27677_ (.A(_05663_),
    .X(_05664_));
 sky130_fd_sc_hd__a21oi_2 _27678_ (.A1(_05628_),
    .A2(_05632_),
    .B1(_05633_),
    .Y(_05665_));
 sky130_fd_sc_hd__nand2_2 _27679_ (.A(_05635_),
    .B(_05659_),
    .Y(_05666_));
 sky130_fd_sc_hd__nor2_2 _27680_ (.A(_05665_),
    .B(_05666_),
    .Y(_05667_));
 sky130_fd_sc_hd__a21oi_2 _27681_ (.A1(_05634_),
    .A2(_05635_),
    .B1(_05659_),
    .Y(_05668_));
 sky130_fd_sc_hd__o21ai_2 _27682_ (.A1(_05667_),
    .A2(_05668_),
    .B1(_05563_),
    .Y(_05669_));
 sky130_fd_sc_hd__buf_1 _27683_ (.A(_19372_),
    .X(_05670_));
 sky130_fd_sc_hd__nand2_2 _27684_ (.A(_05670_),
    .B(_19640_),
    .Y(_05671_));
 sky130_fd_sc_hd__buf_1 _27685_ (.A(\pcpi_mul.rs2[9] ),
    .X(_05672_));
 sky130_fd_sc_hd__buf_1 _27686_ (.A(_05672_),
    .X(_05673_));
 sky130_fd_sc_hd__nand2_2 _27687_ (.A(_05673_),
    .B(_19636_),
    .Y(_05674_));
 sky130_fd_sc_hd__nor2_2 _27688_ (.A(_05671_),
    .B(_05674_),
    .Y(_05675_));
 sky130_fd_sc_hd__nand2_2 _27689_ (.A(_05671_),
    .B(_05674_),
    .Y(_05676_));
 sky130_fd_sc_hd__inv_2 _27690_ (.A(_05676_),
    .Y(_05677_));
 sky130_fd_sc_hd__o2bb2ai_2 _27691_ (.A1_N(_05664_),
    .A2_N(_05669_),
    .B1(_05675_),
    .B2(_05677_),
    .Y(_05678_));
 sky130_fd_sc_hd__inv_2 _27692_ (.A(_05675_),
    .Y(_05679_));
 sky130_fd_sc_hd__nand2_2 _27693_ (.A(_05679_),
    .B(_05676_),
    .Y(_05680_));
 sky130_fd_sc_hd__inv_2 _27694_ (.A(_05680_),
    .Y(_05681_));
 sky130_fd_sc_hd__nand3_2 _27695_ (.A(_05669_),
    .B(_05664_),
    .C(_05681_),
    .Y(_05682_));
 sky130_fd_sc_hd__nand2_2 _27696_ (.A(_05574_),
    .B(_05575_),
    .Y(_05683_));
 sky130_fd_sc_hd__nor2_2 _27697_ (.A(_05570_),
    .B(_05683_),
    .Y(_05684_));
 sky130_fd_sc_hd__a21oi_2 _27698_ (.A1(_05678_),
    .A2(_05682_),
    .B1(_05684_),
    .Y(_05685_));
 sky130_fd_sc_hd__a21oi_2 _27699_ (.A1(_05669_),
    .A2(_05664_),
    .B1(_05681_),
    .Y(_05686_));
 sky130_fd_sc_hd__and3_2 _27700_ (.A(_05669_),
    .B(_05663_),
    .C(_05681_),
    .X(_05687_));
 sky130_fd_sc_hd__buf_1 _27701_ (.A(_05687_),
    .X(_05688_));
 sky130_fd_sc_hd__nor3_2 _27702_ (.A(_05576_),
    .B(_05686_),
    .C(_05688_),
    .Y(_05689_));
 sky130_fd_sc_hd__a21boi_2 _27703_ (.A1(_05561_),
    .A2(_05537_),
    .B1_N(_05533_),
    .Y(_05690_));
 sky130_fd_sc_hd__nor2_2 _27704_ (.A(_05690_),
    .B(_05572_),
    .Y(_05691_));
 sky130_fd_sc_hd__and2_2 _27705_ (.A(_05572_),
    .B(_05690_),
    .X(_05692_));
 sky130_fd_sc_hd__nor2_2 _27706_ (.A(_05691_),
    .B(_05692_),
    .Y(_05693_));
 sky130_fd_sc_hd__o21ai_2 _27707_ (.A1(_05685_),
    .A2(_05689_),
    .B1(_05693_),
    .Y(_05694_));
 sky130_fd_sc_hd__nand2_2 _27708_ (.A(_05585_),
    .B(_05495_),
    .Y(_05695_));
 sky130_fd_sc_hd__inv_2 _27709_ (.A(_05695_),
    .Y(_05696_));
 sky130_fd_sc_hd__o22ai_2 _27710_ (.A1(_05570_),
    .A2(_05683_),
    .B1(_05686_),
    .B2(_05688_),
    .Y(_05697_));
 sky130_fd_sc_hd__nand3_2 _27711_ (.A(_05684_),
    .B(_05682_),
    .C(_05678_),
    .Y(_05698_));
 sky130_fd_sc_hd__nand2_2 _27712_ (.A(_05572_),
    .B(_05690_),
    .Y(_05699_));
 sky130_fd_sc_hd__or2b_2 _27713_ (.A(_05691_),
    .B_N(_05699_),
    .X(_05700_));
 sky130_fd_sc_hd__nand3_2 _27714_ (.A(_05697_),
    .B(_05698_),
    .C(_05700_),
    .Y(_05701_));
 sky130_fd_sc_hd__nand3_2 _27715_ (.A(_05694_),
    .B(_05696_),
    .C(_05701_),
    .Y(_05702_));
 sky130_fd_sc_hd__inv_2 _27716_ (.A(_05586_),
    .Y(_05703_));
 sky130_fd_sc_hd__and2_2 _27717_ (.A(_05702_),
    .B(_05703_),
    .X(_05704_));
 sky130_fd_sc_hd__o22ai_2 _27718_ (.A1(_05692_),
    .A2(_05691_),
    .B1(_05685_),
    .B2(_05689_),
    .Y(_05705_));
 sky130_fd_sc_hd__nand3_2 _27719_ (.A(_05697_),
    .B(_05698_),
    .C(_05693_),
    .Y(_05706_));
 sky130_fd_sc_hd__nand3_2 _27720_ (.A(_05705_),
    .B(_05706_),
    .C(_05695_),
    .Y(_05707_));
 sky130_fd_sc_hd__nand2_2 _27721_ (.A(_05584_),
    .B(_05585_),
    .Y(_05708_));
 sky130_fd_sc_hd__o2bb2ai_2 _27722_ (.A1_N(_05707_),
    .A2_N(_05702_),
    .B1(_05582_),
    .B2(_05708_),
    .Y(_05709_));
 sky130_fd_sc_hd__and2b_2 _27723_ (.A_N(_05704_),
    .B(_05709_),
    .X(_05710_));
 sky130_fd_sc_hd__xor2_2 _27724_ (.A(_05591_),
    .B(_05710_),
    .X(_02629_));
 sky130_fd_sc_hd__a22oi_2 _27725_ (.A1(_05703_),
    .A2(_05702_),
    .B1(_05591_),
    .B2(_05709_),
    .Y(_05711_));
 sky130_fd_sc_hd__buf_1 _27726_ (.A(_05187_),
    .X(_05712_));
 sky130_fd_sc_hd__buf_1 _27727_ (.A(_05420_),
    .X(_05713_));
 sky130_fd_sc_hd__a22oi_2 _27728_ (.A1(_05712_),
    .A2(_05343_),
    .B1(_05403_),
    .B2(_05713_),
    .Y(_05714_));
 sky130_fd_sc_hd__and4_2 _27729_ (.A(_19387_),
    .B(_19390_),
    .C(_19618_),
    .D(_05251_),
    .X(_05715_));
 sky130_fd_sc_hd__buf_1 _27730_ (.A(_05715_),
    .X(_05716_));
 sky130_fd_sc_hd__buf_1 _27731_ (.A(_19605_),
    .X(_05717_));
 sky130_fd_sc_hd__nand2_2 _27732_ (.A(_05192_),
    .B(_05717_),
    .Y(_05718_));
 sky130_fd_sc_hd__inv_2 _27733_ (.A(_05718_),
    .Y(_05719_));
 sky130_fd_sc_hd__o21ai_2 _27734_ (.A1(_05714_),
    .A2(_05716_),
    .B1(_05719_),
    .Y(_05720_));
 sky130_fd_sc_hd__buf_1 _27735_ (.A(_05155_),
    .X(_05721_));
 sky130_fd_sc_hd__a22o_2 _27736_ (.A1(_05402_),
    .A2(_05343_),
    .B1(_05721_),
    .B2(_05421_),
    .X(_05722_));
 sky130_fd_sc_hd__nand3b_2 _27737_ (.A_N(_05716_),
    .B(_05718_),
    .C(_05722_),
    .Y(_05723_));
 sky130_fd_sc_hd__o2111ai_2 _27738_ (.A1(_05594_),
    .A2(_05595_),
    .B1(_05602_),
    .C1(_05720_),
    .D1(_05723_),
    .Y(_05724_));
 sky130_fd_sc_hd__nand2_2 _27739_ (.A(_05722_),
    .B(_05719_),
    .Y(_05725_));
 sky130_fd_sc_hd__o21ai_2 _27740_ (.A1(_05714_),
    .A2(_05716_),
    .B1(_05718_),
    .Y(_05726_));
 sky130_fd_sc_hd__nand2_2 _27741_ (.A(_05608_),
    .B(_05602_),
    .Y(_05727_));
 sky130_fd_sc_hd__o211ai_2 _27742_ (.A1(_05716_),
    .A2(_05725_),
    .B1(_05726_),
    .C1(_05727_),
    .Y(_05728_));
 sky130_fd_sc_hd__nand2_2 _27743_ (.A(_05724_),
    .B(_05728_),
    .Y(_05729_));
 sky130_fd_sc_hd__buf_1 _27744_ (.A(\pcpi_mul.rs1[8] ),
    .X(_05730_));
 sky130_fd_sc_hd__inv_2 _27745_ (.A(_05730_),
    .Y(_05731_));
 sky130_fd_sc_hd__buf_1 _27746_ (.A(_05731_),
    .X(_05732_));
 sky130_fd_sc_hd__buf_1 _27747_ (.A(_05597_),
    .X(_05733_));
 sky130_fd_sc_hd__buf_1 _27748_ (.A(_19612_),
    .X(_05734_));
 sky130_fd_sc_hd__nand2_2 _27749_ (.A(_05733_),
    .B(_05734_),
    .Y(_05735_));
 sky130_fd_sc_hd__buf_1 _27750_ (.A(_05122_),
    .X(_05736_));
 sky130_fd_sc_hd__buf_1 _27751_ (.A(_05516_),
    .X(_05737_));
 sky130_fd_sc_hd__buf_1 _27752_ (.A(_19608_),
    .X(_05738_));
 sky130_fd_sc_hd__a22o_2 _27753_ (.A1(_05736_),
    .A2(_05737_),
    .B1(_05118_),
    .B2(_05738_),
    .X(_05739_));
 sky130_fd_sc_hd__o21ai_2 _27754_ (.A1(_05103_),
    .A2(_05735_),
    .B1(_05739_),
    .Y(_05740_));
 sky130_fd_sc_hd__o21ai_2 _27755_ (.A1(_05151_),
    .A2(_05732_),
    .B1(_05740_),
    .Y(_05741_));
 sky130_fd_sc_hd__o2111ai_2 _27756_ (.A1(_05103_),
    .A2(_05735_),
    .B1(_05116_),
    .C1(_19617_),
    .D1(_05739_),
    .Y(_05742_));
 sky130_fd_sc_hd__nand2_2 _27757_ (.A(_05741_),
    .B(_05742_),
    .Y(_05743_));
 sky130_fd_sc_hd__nand2_2 _27758_ (.A(_05729_),
    .B(_05743_),
    .Y(_05744_));
 sky130_fd_sc_hd__nand2_2 _27759_ (.A(_05611_),
    .B(_05626_),
    .Y(_05745_));
 sky130_fd_sc_hd__nand2_2 _27760_ (.A(_05745_),
    .B(_05606_),
    .Y(_05746_));
 sky130_fd_sc_hd__and2_2 _27761_ (.A(_05741_),
    .B(_05742_),
    .X(_05747_));
 sky130_fd_sc_hd__nand3_2 _27762_ (.A(_05747_),
    .B(_05728_),
    .C(_05724_),
    .Y(_05748_));
 sky130_fd_sc_hd__nand3_2 _27763_ (.A(_05744_),
    .B(_05746_),
    .C(_05748_),
    .Y(_05749_));
 sky130_fd_sc_hd__nand2_2 _27764_ (.A(_05729_),
    .B(_05747_),
    .Y(_05750_));
 sky130_fd_sc_hd__a21boi_2 _27765_ (.A1(_05626_),
    .A2(_05611_),
    .B1_N(_05606_),
    .Y(_05751_));
 sky130_fd_sc_hd__nand3_2 _27766_ (.A(_05724_),
    .B(_05728_),
    .C(_05743_),
    .Y(_05752_));
 sky130_fd_sc_hd__nand3_2 _27767_ (.A(_05750_),
    .B(_05751_),
    .C(_05752_),
    .Y(_05753_));
 sky130_fd_sc_hd__nor2_2 _27768_ (.A(_05622_),
    .B(_05618_),
    .Y(_05754_));
 sky130_fd_sc_hd__o2bb2ai_2 _27769_ (.A1_N(_05749_),
    .A2_N(_05753_),
    .B1(_05616_),
    .B2(_05754_),
    .Y(_05755_));
 sky130_fd_sc_hd__nor2_2 _27770_ (.A(_05616_),
    .B(_05754_),
    .Y(_05756_));
 sky130_fd_sc_hd__nand3_2 _27771_ (.A(_05749_),
    .B(_05753_),
    .C(_05756_),
    .Y(_05757_));
 sky130_fd_sc_hd__buf_1 _27772_ (.A(_05447_),
    .X(_05758_));
 sky130_fd_sc_hd__nand2_2 _27773_ (.A(_05758_),
    .B(_05218_),
    .Y(_05759_));
 sky130_fd_sc_hd__buf_1 _27774_ (.A(\pcpi_mul.rs2[7] ),
    .X(_05760_));
 sky130_fd_sc_hd__nand2_2 _27775_ (.A(_05760_),
    .B(_19627_),
    .Y(_05761_));
 sky130_fd_sc_hd__nor2_2 _27776_ (.A(_05759_),
    .B(_05761_),
    .Y(_05762_));
 sky130_fd_sc_hd__buf_1 _27777_ (.A(\pcpi_mul.rs2[6] ),
    .X(_05763_));
 sky130_fd_sc_hd__buf_1 _27778_ (.A(_05763_),
    .X(_05764_));
 sky130_fd_sc_hd__buf_1 _27779_ (.A(_05193_),
    .X(_05765_));
 sky130_fd_sc_hd__nand2_2 _27780_ (.A(_05764_),
    .B(_05765_),
    .Y(_05766_));
 sky130_fd_sc_hd__inv_2 _27781_ (.A(_05766_),
    .Y(_05767_));
 sky130_fd_sc_hd__nand2_2 _27782_ (.A(_05759_),
    .B(_05761_),
    .Y(_05768_));
 sky130_fd_sc_hd__nand2_2 _27783_ (.A(_05767_),
    .B(_05768_),
    .Y(_05769_));
 sky130_fd_sc_hd__and2_2 _27784_ (.A(_05759_),
    .B(_05761_),
    .X(_05770_));
 sky130_fd_sc_hd__o21ai_2 _27785_ (.A1(_05762_),
    .A2(_05770_),
    .B1(_05766_),
    .Y(_05771_));
 sky130_fd_sc_hd__o211ai_2 _27786_ (.A1(_05762_),
    .A2(_05769_),
    .B1(_05675_),
    .C1(_05771_),
    .Y(_05772_));
 sky130_fd_sc_hd__o21ai_2 _27787_ (.A1(_05762_),
    .A2(_05770_),
    .B1(_05767_),
    .Y(_05773_));
 sky130_fd_sc_hd__nand3b_2 _27788_ (.A_N(_05762_),
    .B(_05768_),
    .C(_05766_),
    .Y(_05774_));
 sky130_fd_sc_hd__nand3_2 _27789_ (.A(_05773_),
    .B(_05774_),
    .C(_05679_),
    .Y(_05775_));
 sky130_fd_sc_hd__a31o_2 _27790_ (.A1(_05645_),
    .A2(_19386_),
    .A3(_19628_),
    .B1(_05643_),
    .X(_05776_));
 sky130_fd_sc_hd__a21oi_2 _27791_ (.A1(_05772_),
    .A2(_05775_),
    .B1(_05776_),
    .Y(_05777_));
 sky130_fd_sc_hd__nand2_2 _27792_ (.A(_05555_),
    .B(_05653_),
    .Y(_05778_));
 sky130_fd_sc_hd__nand2_2 _27793_ (.A(_05778_),
    .B(_05652_),
    .Y(_05779_));
 sky130_fd_sc_hd__nand3_2 _27794_ (.A(_05772_),
    .B(_05775_),
    .C(_05776_),
    .Y(_05780_));
 sky130_fd_sc_hd__nand2_2 _27795_ (.A(_05779_),
    .B(_05780_),
    .Y(_05781_));
 sky130_fd_sc_hd__inv_2 _27796_ (.A(_05653_),
    .Y(_05782_));
 sky130_fd_sc_hd__a21oi_2 _27797_ (.A1(_05649_),
    .A2(_05651_),
    .B1(_05555_),
    .Y(_05783_));
 sky130_fd_sc_hd__a21o_2 _27798_ (.A1(_05772_),
    .A2(_05775_),
    .B1(_05776_),
    .X(_05784_));
 sky130_fd_sc_hd__nand2_2 _27799_ (.A(_05784_),
    .B(_05780_),
    .Y(_05785_));
 sky130_fd_sc_hd__o21ai_2 _27800_ (.A1(_05782_),
    .A2(_05783_),
    .B1(_05785_),
    .Y(_05786_));
 sky130_fd_sc_hd__o21ai_2 _27801_ (.A1(_05777_),
    .A2(_05781_),
    .B1(_05786_),
    .Y(_05787_));
 sky130_fd_sc_hd__a21oi_2 _27802_ (.A1(_05755_),
    .A2(_05757_),
    .B1(_05787_),
    .Y(_05788_));
 sky130_fd_sc_hd__and3_2 _27803_ (.A(_05744_),
    .B(_05746_),
    .C(_05748_),
    .X(_05789_));
 sky130_fd_sc_hd__nand2_2 _27804_ (.A(_05753_),
    .B(_05756_),
    .Y(_05790_));
 sky130_fd_sc_hd__o211a_2 _27805_ (.A1(_05789_),
    .A2(_05790_),
    .B1(_05755_),
    .C1(_05787_),
    .X(_05791_));
 sky130_fd_sc_hd__o22a_2 _27806_ (.A1(_05565_),
    .A2(_05654_),
    .B1(_05665_),
    .B2(_05666_),
    .X(_05792_));
 sky130_fd_sc_hd__o21ai_2 _27807_ (.A1(_05788_),
    .A2(_05791_),
    .B1(_05792_),
    .Y(_05793_));
 sky130_fd_sc_hd__a21o_2 _27808_ (.A1(_05755_),
    .A2(_05757_),
    .B1(_05787_),
    .X(_05794_));
 sky130_fd_sc_hd__o22ai_2 _27809_ (.A1(_05565_),
    .A2(_05654_),
    .B1(_05665_),
    .B2(_05666_),
    .Y(_05795_));
 sky130_fd_sc_hd__nand3_2 _27810_ (.A(_05787_),
    .B(_05755_),
    .C(_05757_),
    .Y(_05796_));
 sky130_fd_sc_hd__nand3_2 _27811_ (.A(_05794_),
    .B(_05795_),
    .C(_05796_),
    .Y(_05797_));
 sky130_fd_sc_hd__nand2_2 _27812_ (.A(_05793_),
    .B(_05797_),
    .Y(_05798_));
 sky130_fd_sc_hd__nor2_2 _27813_ (.A(_05497_),
    .B(_05256_),
    .Y(_05799_));
 sky130_fd_sc_hd__buf_1 _27814_ (.A(\pcpi_mul.rs2[11] ),
    .X(_05800_));
 sky130_fd_sc_hd__buf_1 _27815_ (.A(_05800_),
    .X(_05801_));
 sky130_fd_sc_hd__buf_1 _27816_ (.A(\pcpi_mul.rs2[10] ),
    .X(_05802_));
 sky130_fd_sc_hd__buf_1 _27817_ (.A(_05802_),
    .X(_05803_));
 sky130_fd_sc_hd__buf_1 _27818_ (.A(_05104_),
    .X(_05804_));
 sky130_fd_sc_hd__buf_1 _27819_ (.A(_19639_),
    .X(_05805_));
 sky130_fd_sc_hd__and4_2 _27820_ (.A(_05801_),
    .B(_05803_),
    .C(_05804_),
    .D(_05805_),
    .X(_05806_));
 sky130_fd_sc_hd__buf_1 _27821_ (.A(_19370_),
    .X(_05807_));
 sky130_fd_sc_hd__buf_1 _27822_ (.A(_05802_),
    .X(_05808_));
 sky130_fd_sc_hd__a22o_2 _27823_ (.A1(_05807_),
    .A2(_05805_),
    .B1(_05808_),
    .B2(_05124_),
    .X(_05809_));
 sky130_fd_sc_hd__and2b_2 _27824_ (.A_N(_05806_),
    .B(_05809_),
    .X(_05810_));
 sky130_fd_sc_hd__xnor2_2 _27825_ (.A(_05799_),
    .B(_05810_),
    .Y(_05811_));
 sky130_fd_sc_hd__nand2_2 _27826_ (.A(_05798_),
    .B(_05811_),
    .Y(_05812_));
 sky130_fd_sc_hd__inv_2 _27827_ (.A(_05811_),
    .Y(_05813_));
 sky130_fd_sc_hd__nand3_2 _27828_ (.A(_05793_),
    .B(_05797_),
    .C(_05813_),
    .Y(_05814_));
 sky130_fd_sc_hd__nand3_2 _27829_ (.A(_05688_),
    .B(_05812_),
    .C(_05814_),
    .Y(_05815_));
 sky130_fd_sc_hd__nand2_2 _27830_ (.A(_05669_),
    .B(_05664_),
    .Y(_05816_));
 sky130_fd_sc_hd__a21oi_2 _27831_ (.A1(_05793_),
    .A2(_05797_),
    .B1(_05813_),
    .Y(_05817_));
 sky130_fd_sc_hd__nand2_2 _27832_ (.A(_05795_),
    .B(_05796_),
    .Y(_05818_));
 sky130_fd_sc_hd__o211a_2 _27833_ (.A1(_05788_),
    .A2(_05818_),
    .B1(_05813_),
    .C1(_05793_),
    .X(_05819_));
 sky130_fd_sc_hd__o22ai_2 _27834_ (.A1(_05680_),
    .A2(_05816_),
    .B1(_05817_),
    .B2(_05819_),
    .Y(_05820_));
 sky130_fd_sc_hd__a21boi_2 _27835_ (.A1(_05632_),
    .A2(_05633_),
    .B1_N(_05628_),
    .Y(_05821_));
 sky130_fd_sc_hd__nor2_2 _27836_ (.A(_05821_),
    .B(_05663_),
    .Y(_05822_));
 sky130_fd_sc_hd__nand2_2 _27837_ (.A(_05664_),
    .B(_05821_),
    .Y(_05823_));
 sky130_fd_sc_hd__inv_2 _27838_ (.A(_05823_),
    .Y(_05824_));
 sky130_fd_sc_hd__o2bb2ai_2 _27839_ (.A1_N(_05815_),
    .A2_N(_05820_),
    .B1(_05822_),
    .B2(_05824_),
    .Y(_05825_));
 sky130_fd_sc_hd__nand2_2 _27840_ (.A(_05684_),
    .B(_05678_),
    .Y(_05826_));
 sky130_fd_sc_hd__o22ai_2 _27841_ (.A1(_05688_),
    .A2(_05826_),
    .B1(_05700_),
    .B2(_05685_),
    .Y(_05827_));
 sky130_fd_sc_hd__nor2_2 _27842_ (.A(_05822_),
    .B(_05824_),
    .Y(_05828_));
 sky130_fd_sc_hd__nand3_2 _27843_ (.A(_05820_),
    .B(_05815_),
    .C(_05828_),
    .Y(_05829_));
 sky130_fd_sc_hd__nand3_2 _27844_ (.A(_05825_),
    .B(_05827_),
    .C(_05829_),
    .Y(_05830_));
 sky130_fd_sc_hd__inv_2 _27845_ (.A(_05663_),
    .Y(_05831_));
 sky130_fd_sc_hd__nor2_2 _27846_ (.A(_05821_),
    .B(_05831_),
    .Y(_05832_));
 sky130_fd_sc_hd__and2_2 _27847_ (.A(_05831_),
    .B(_05821_),
    .X(_05833_));
 sky130_fd_sc_hd__o2bb2ai_2 _27848_ (.A1_N(_05815_),
    .A2_N(_05820_),
    .B1(_05832_),
    .B2(_05833_),
    .Y(_05834_));
 sky130_fd_sc_hd__a21oi_2 _27849_ (.A1(_05697_),
    .A2(_05693_),
    .B1(_05689_),
    .Y(_05835_));
 sky130_fd_sc_hd__inv_2 _27850_ (.A(_05822_),
    .Y(_05836_));
 sky130_fd_sc_hd__nand2_2 _27851_ (.A(_05836_),
    .B(_05823_),
    .Y(_05837_));
 sky130_fd_sc_hd__nand3_2 _27852_ (.A(_05820_),
    .B(_05815_),
    .C(_05837_),
    .Y(_05838_));
 sky130_fd_sc_hd__nand3_2 _27853_ (.A(_05834_),
    .B(_05835_),
    .C(_05838_),
    .Y(_05839_));
 sky130_fd_sc_hd__o2bb2ai_2 _27854_ (.A1_N(_05830_),
    .A2_N(_05839_),
    .B1(_05572_),
    .B2(_05690_),
    .Y(_05840_));
 sky130_fd_sc_hd__nand2_2 _27855_ (.A(_05839_),
    .B(_05691_),
    .Y(_05841_));
 sky130_fd_sc_hd__inv_2 _27856_ (.A(_05707_),
    .Y(_05842_));
 sky130_fd_sc_hd__a21oi_2 _27857_ (.A1(_05840_),
    .A2(_05841_),
    .B1(_05842_),
    .Y(_05843_));
 sky130_fd_sc_hd__inv_2 _27858_ (.A(_05841_),
    .Y(_05844_));
 sky130_fd_sc_hd__nand2_2 _27859_ (.A(_05840_),
    .B(_05842_),
    .Y(_05845_));
 sky130_fd_sc_hd__nor2_2 _27860_ (.A(_05844_),
    .B(_05845_),
    .Y(_05846_));
 sky130_fd_sc_hd__or2_2 _27861_ (.A(_05843_),
    .B(_05846_),
    .X(_05847_));
 sky130_fd_sc_hd__nand2_2 _27862_ (.A(_05847_),
    .B(_05711_),
    .Y(_05848_));
 sky130_fd_sc_hd__o21a_2 _27863_ (.A1(_05711_),
    .A2(_05843_),
    .B1(_05848_),
    .X(_02630_));
 sky130_fd_sc_hd__inv_2 _27864_ (.A(\pcpi_mul.rs1[4] ),
    .Y(_05849_));
 sky130_fd_sc_hd__buf_1 _27865_ (.A(_05849_),
    .X(_05850_));
 sky130_fd_sc_hd__buf_1 _27866_ (.A(_05447_),
    .X(_05851_));
 sky130_fd_sc_hd__nand3_2 _27867_ (.A(_05851_),
    .B(_19383_),
    .C(_05194_),
    .Y(_05852_));
 sky130_fd_sc_hd__nor2_2 _27868_ (.A(_05850_),
    .B(_05852_),
    .Y(_05853_));
 sky130_fd_sc_hd__inv_2 _27869_ (.A(_05641_),
    .Y(_05854_));
 sky130_fd_sc_hd__inv_2 _27870_ (.A(\pcpi_mul.rs1[5] ),
    .Y(_05855_));
 sky130_fd_sc_hd__buf_1 _27871_ (.A(_05855_),
    .X(_05856_));
 sky130_fd_sc_hd__buf_1 _27872_ (.A(_19379_),
    .X(_05857_));
 sky130_fd_sc_hd__nand2_2 _27873_ (.A(_05857_),
    .B(_05338_),
    .Y(_05858_));
 sky130_fd_sc_hd__o21a_2 _27874_ (.A1(_05854_),
    .A2(_05856_),
    .B1(_05858_),
    .X(_05859_));
 sky130_fd_sc_hd__nand2_2 _27875_ (.A(_05764_),
    .B(_05425_),
    .Y(_05860_));
 sky130_fd_sc_hd__o21ai_2 _27876_ (.A1(_05853_),
    .A2(_05859_),
    .B1(_05860_),
    .Y(_05861_));
 sky130_fd_sc_hd__a21o_2 _27877_ (.A1(_05799_),
    .A2(_05809_),
    .B1(_05806_),
    .X(_05862_));
 sky130_fd_sc_hd__or2_2 _27878_ (.A(_05850_),
    .B(_05852_),
    .X(_05863_));
 sky130_fd_sc_hd__inv_2 _27879_ (.A(_05860_),
    .Y(_05864_));
 sky130_fd_sc_hd__buf_1 _27880_ (.A(_05856_),
    .X(_05865_));
 sky130_fd_sc_hd__o21ai_2 _27881_ (.A1(_05854_),
    .A2(_05865_),
    .B1(_05858_),
    .Y(_05866_));
 sky130_fd_sc_hd__nand3_2 _27882_ (.A(_05863_),
    .B(_05864_),
    .C(_05866_),
    .Y(_05867_));
 sky130_fd_sc_hd__nand3_2 _27883_ (.A(_05861_),
    .B(_05862_),
    .C(_05867_),
    .Y(_05868_));
 sky130_fd_sc_hd__o21ai_2 _27884_ (.A1(_05853_),
    .A2(_05859_),
    .B1(_05864_),
    .Y(_05869_));
 sky130_fd_sc_hd__a21oi_2 _27885_ (.A1(_05799_),
    .A2(_05809_),
    .B1(_05806_),
    .Y(_05870_));
 sky130_fd_sc_hd__nand3_2 _27886_ (.A(_05863_),
    .B(_05860_),
    .C(_05866_),
    .Y(_05871_));
 sky130_fd_sc_hd__nand3_2 _27887_ (.A(_05869_),
    .B(_05870_),
    .C(_05871_),
    .Y(_05872_));
 sky130_fd_sc_hd__nand2_2 _27888_ (.A(_05868_),
    .B(_05872_),
    .Y(_05873_));
 sky130_fd_sc_hd__a21oi_2 _27889_ (.A1(_05767_),
    .A2(_05768_),
    .B1(_05762_),
    .Y(_05874_));
 sky130_fd_sc_hd__nand2_2 _27890_ (.A(_05873_),
    .B(_05874_),
    .Y(_05875_));
 sky130_fd_sc_hd__inv_2 _27891_ (.A(_05874_),
    .Y(_05876_));
 sky130_fd_sc_hd__nand3_2 _27892_ (.A(_05868_),
    .B(_05872_),
    .C(_05876_),
    .Y(_05877_));
 sky130_fd_sc_hd__nand2_2 _27893_ (.A(_05875_),
    .B(_05877_),
    .Y(_05878_));
 sky130_fd_sc_hd__nand2_2 _27894_ (.A(_05775_),
    .B(_05776_),
    .Y(_05879_));
 sky130_fd_sc_hd__nand2_2 _27895_ (.A(_05879_),
    .B(_05772_),
    .Y(_05880_));
 sky130_fd_sc_hd__inv_2 _27896_ (.A(_05880_),
    .Y(_05881_));
 sky130_fd_sc_hd__nand2_2 _27897_ (.A(_05878_),
    .B(_05881_),
    .Y(_05882_));
 sky130_fd_sc_hd__nand2_2 _27898_ (.A(_05782_),
    .B(_05780_),
    .Y(_05883_));
 sky130_fd_sc_hd__nor2_2 _27899_ (.A(_05777_),
    .B(_05883_),
    .Y(_05884_));
 sky130_fd_sc_hd__nand3_2 _27900_ (.A(_05875_),
    .B(_05880_),
    .C(_05877_),
    .Y(_05885_));
 sky130_fd_sc_hd__nand3_2 _27901_ (.A(_05882_),
    .B(_05884_),
    .C(_05885_),
    .Y(_05886_));
 sky130_fd_sc_hd__a21oi_2 _27902_ (.A1(_05875_),
    .A2(_05877_),
    .B1(_05880_),
    .Y(_05887_));
 sky130_fd_sc_hd__and3_2 _27903_ (.A(_05875_),
    .B(_05880_),
    .C(_05877_),
    .X(_05888_));
 sky130_fd_sc_hd__o22ai_2 _27904_ (.A1(_05653_),
    .A2(_05785_),
    .B1(_05887_),
    .B2(_05888_),
    .Y(_05889_));
 sky130_fd_sc_hd__a21bo_2 _27905_ (.A1(_05747_),
    .A2(_05724_),
    .B1_N(_05728_),
    .X(_05890_));
 sky130_fd_sc_hd__buf_1 _27906_ (.A(_19390_),
    .X(_05891_));
 sky130_fd_sc_hd__buf_1 _27907_ (.A(_05891_),
    .X(_05892_));
 sky130_fd_sc_hd__buf_1 _27908_ (.A(_05408_),
    .X(_05893_));
 sky130_fd_sc_hd__a22oi_2 _27909_ (.A1(_05712_),
    .A2(_05713_),
    .B1(_05892_),
    .B2(_05893_),
    .Y(_05894_));
 sky130_fd_sc_hd__and4_2 _27910_ (.A(_19388_),
    .B(_19391_),
    .C(_19616_),
    .D(_19619_),
    .X(_05895_));
 sky130_fd_sc_hd__buf_1 _27911_ (.A(\pcpi_mul.rs1[12] ),
    .X(_05896_));
 sky130_fd_sc_hd__buf_1 _27912_ (.A(_05896_),
    .X(_05897_));
 sky130_fd_sc_hd__nand2_2 _27913_ (.A(_05192_),
    .B(_05897_),
    .Y(_05898_));
 sky130_fd_sc_hd__o21ai_2 _27914_ (.A1(_05894_),
    .A2(_05895_),
    .B1(_05898_),
    .Y(_05899_));
 sky130_fd_sc_hd__inv_2 _27915_ (.A(_05898_),
    .Y(_05900_));
 sky130_fd_sc_hd__a22o_2 _27916_ (.A1(_05402_),
    .A2(_05421_),
    .B1(_05721_),
    .B2(_05893_),
    .X(_05901_));
 sky130_fd_sc_hd__nand3b_2 _27917_ (.A_N(_05895_),
    .B(_05900_),
    .C(_05901_),
    .Y(_05902_));
 sky130_fd_sc_hd__nor2_2 _27918_ (.A(_05719_),
    .B(_05716_),
    .Y(_05903_));
 sky130_fd_sc_hd__o2bb2ai_2 _27919_ (.A1_N(_05899_),
    .A2_N(_05902_),
    .B1(_05714_),
    .B2(_05903_),
    .Y(_05904_));
 sky130_fd_sc_hd__a21o_2 _27920_ (.A1(_05722_),
    .A2(_05719_),
    .B1(_05716_),
    .X(_05905_));
 sky130_fd_sc_hd__nand3_2 _27921_ (.A(_05905_),
    .B(_05902_),
    .C(_05899_),
    .Y(_05906_));
 sky130_fd_sc_hd__nand2_2 _27922_ (.A(_05904_),
    .B(_05906_),
    .Y(_05907_));
 sky130_fd_sc_hd__nand2_2 _27923_ (.A(_05123_),
    .B(_05738_),
    .Y(_05908_));
 sky130_fd_sc_hd__buf_1 _27924_ (.A(_19400_),
    .X(_05909_));
 sky130_fd_sc_hd__buf_1 _27925_ (.A(\pcpi_mul.rs1[11] ),
    .X(_05910_));
 sky130_fd_sc_hd__buf_1 _27926_ (.A(_05910_),
    .X(_05911_));
 sky130_fd_sc_hd__nand2_2 _27927_ (.A(_05909_),
    .B(_05911_),
    .Y(_05912_));
 sky130_fd_sc_hd__nor2_2 _27928_ (.A(_05908_),
    .B(_05912_),
    .Y(_05913_));
 sky130_fd_sc_hd__and2_2 _27929_ (.A(_05908_),
    .B(_05912_),
    .X(_05914_));
 sky130_fd_sc_hd__nor2_2 _27930_ (.A(_05913_),
    .B(_05914_),
    .Y(_05915_));
 sky130_fd_sc_hd__nand3_2 _27931_ (.A(_05915_),
    .B(_19395_),
    .C(_19614_),
    .Y(_05916_));
 sky130_fd_sc_hd__nand2_2 _27932_ (.A(_19394_),
    .B(_19614_),
    .Y(_05917_));
 sky130_fd_sc_hd__o21ai_2 _27933_ (.A1(_05913_),
    .A2(_05914_),
    .B1(_05917_),
    .Y(_05918_));
 sky130_fd_sc_hd__nand2_2 _27934_ (.A(_05916_),
    .B(_05918_),
    .Y(_05919_));
 sky130_fd_sc_hd__nand2_2 _27935_ (.A(_05907_),
    .B(_05919_),
    .Y(_05920_));
 sky130_fd_sc_hd__nor3_2 _27936_ (.A(_05917_),
    .B(_05913_),
    .C(_05914_),
    .Y(_05921_));
 sky130_fd_sc_hd__and2b_2 _27937_ (.A_N(_05921_),
    .B(_05918_),
    .X(_05922_));
 sky130_fd_sc_hd__nand3_2 _27938_ (.A(_05922_),
    .B(_05904_),
    .C(_05906_),
    .Y(_05923_));
 sky130_fd_sc_hd__nand3_2 _27939_ (.A(_05890_),
    .B(_05920_),
    .C(_05923_),
    .Y(_05924_));
 sky130_fd_sc_hd__nand2_2 _27940_ (.A(_05907_),
    .B(_05922_),
    .Y(_05925_));
 sky130_fd_sc_hd__a21boi_2 _27941_ (.A1(_05747_),
    .A2(_05724_),
    .B1_N(_05728_),
    .Y(_05926_));
 sky130_fd_sc_hd__nand3_2 _27942_ (.A(_05919_),
    .B(_05904_),
    .C(_05906_),
    .Y(_05927_));
 sky130_fd_sc_hd__nand3_2 _27943_ (.A(_05925_),
    .B(_05926_),
    .C(_05927_),
    .Y(_05928_));
 sky130_fd_sc_hd__nor2_2 _27944_ (.A(_05103_),
    .B(_05735_),
    .Y(_05929_));
 sky130_fd_sc_hd__inv_2 _27945_ (.A(_05742_),
    .Y(_05930_));
 sky130_fd_sc_hd__nor2_2 _27946_ (.A(_05929_),
    .B(_05930_),
    .Y(_05931_));
 sky130_fd_sc_hd__inv_2 _27947_ (.A(_05931_),
    .Y(_05932_));
 sky130_fd_sc_hd__a21oi_2 _27948_ (.A1(_05924_),
    .A2(_05928_),
    .B1(_05932_),
    .Y(_05933_));
 sky130_fd_sc_hd__nand2_2 _27949_ (.A(_05924_),
    .B(_05928_),
    .Y(_05934_));
 sky130_fd_sc_hd__nor2_2 _27950_ (.A(_05931_),
    .B(_05934_),
    .Y(_05935_));
 sky130_fd_sc_hd__o2bb2ai_2 _27951_ (.A1_N(_05886_),
    .A2_N(_05889_),
    .B1(_05933_),
    .B2(_05935_),
    .Y(_05936_));
 sky130_fd_sc_hd__nand2_2 _27952_ (.A(_05783_),
    .B(_05653_),
    .Y(_05937_));
 sky130_fd_sc_hd__o21ai_2 _27953_ (.A1(_05785_),
    .A2(_05937_),
    .B1(_05796_),
    .Y(_05938_));
 sky130_fd_sc_hd__and3_2 _27954_ (.A(_05890_),
    .B(_05920_),
    .C(_05923_),
    .X(_05939_));
 sky130_fd_sc_hd__nand2_2 _27955_ (.A(_05928_),
    .B(_05932_),
    .Y(_05940_));
 sky130_fd_sc_hd__nand2_2 _27956_ (.A(_05934_),
    .B(_05931_),
    .Y(_05941_));
 sky130_fd_sc_hd__o2111ai_2 _27957_ (.A1(_05939_),
    .A2(_05940_),
    .B1(_05886_),
    .C1(_05941_),
    .D1(_05889_),
    .Y(_05942_));
 sky130_fd_sc_hd__nand3_2 _27958_ (.A(_05936_),
    .B(_05938_),
    .C(_05942_),
    .Y(_05943_));
 sky130_fd_sc_hd__a21oi_2 _27959_ (.A1(_05924_),
    .A2(_05928_),
    .B1(_05931_),
    .Y(_05944_));
 sky130_fd_sc_hd__nand3_2 _27960_ (.A(_05924_),
    .B(_05928_),
    .C(_05931_),
    .Y(_05945_));
 sky130_fd_sc_hd__inv_2 _27961_ (.A(_05945_),
    .Y(_05946_));
 sky130_fd_sc_hd__o2bb2ai_2 _27962_ (.A1_N(_05886_),
    .A2_N(_05889_),
    .B1(_05944_),
    .B2(_05946_),
    .Y(_05947_));
 sky130_fd_sc_hd__nor2_2 _27963_ (.A(_05785_),
    .B(_05937_),
    .Y(_05948_));
 sky130_fd_sc_hd__a31oi_2 _27964_ (.A1(_05787_),
    .A2(_05755_),
    .A3(_05757_),
    .B1(_05948_),
    .Y(_05949_));
 sky130_fd_sc_hd__nand2_2 _27965_ (.A(_05884_),
    .B(_05885_),
    .Y(_05950_));
 sky130_fd_sc_hd__nand2_2 _27966_ (.A(_05934_),
    .B(_05932_),
    .Y(_05951_));
 sky130_fd_sc_hd__o2111ai_2 _27967_ (.A1(_05887_),
    .A2(_05950_),
    .B1(_05945_),
    .C1(_05951_),
    .D1(_05889_),
    .Y(_05952_));
 sky130_fd_sc_hd__nand3_2 _27968_ (.A(_05947_),
    .B(_05949_),
    .C(_05952_),
    .Y(_05953_));
 sky130_fd_sc_hd__nor2_2 _27969_ (.A(_05497_),
    .B(_05320_),
    .Y(_05954_));
 sky130_fd_sc_hd__buf_1 _27970_ (.A(\pcpi_mul.rs2[11] ),
    .X(_05955_));
 sky130_fd_sc_hd__buf_1 _27971_ (.A(_05955_),
    .X(_05956_));
 sky130_fd_sc_hd__nand2_2 _27972_ (.A(_05956_),
    .B(_05543_),
    .Y(_05957_));
 sky130_fd_sc_hd__buf_1 _27973_ (.A(_19372_),
    .X(_05958_));
 sky130_fd_sc_hd__nand2_2 _27974_ (.A(_05958_),
    .B(_05119_),
    .Y(_05959_));
 sky130_fd_sc_hd__nor2_2 _27975_ (.A(_05957_),
    .B(_05959_),
    .Y(_05960_));
 sky130_fd_sc_hd__nand2_2 _27976_ (.A(_05957_),
    .B(_05959_),
    .Y(_05961_));
 sky130_fd_sc_hd__or3b_2 _27977_ (.A(_05954_),
    .B(_05960_),
    .C_N(_05961_),
    .X(_05962_));
 sky130_fd_sc_hd__nand2_2 _27978_ (.A(_19369_),
    .B(_19642_),
    .Y(_05963_));
 sky130_fd_sc_hd__inv_2 _27979_ (.A(_05963_),
    .Y(_05964_));
 sky130_fd_sc_hd__or2_2 _27980_ (.A(_05957_),
    .B(_05959_),
    .X(_05965_));
 sky130_fd_sc_hd__nand2_2 _27981_ (.A(_05965_),
    .B(_05961_),
    .Y(_05966_));
 sky130_fd_sc_hd__nand2_2 _27982_ (.A(_05966_),
    .B(_05954_),
    .Y(_05967_));
 sky130_fd_sc_hd__and3_2 _27983_ (.A(_05962_),
    .B(_05964_),
    .C(_05967_),
    .X(_05968_));
 sky130_fd_sc_hd__nor2_2 _27984_ (.A(_05954_),
    .B(_05966_),
    .Y(_05969_));
 sky130_fd_sc_hd__and2b_2 _27985_ (.A_N(_05969_),
    .B(_05967_),
    .X(_05970_));
 sky130_fd_sc_hd__nor2_2 _27986_ (.A(_05964_),
    .B(_05970_),
    .Y(_05971_));
 sky130_fd_sc_hd__or2_2 _27987_ (.A(_05968_),
    .B(_05971_),
    .X(_05972_));
 sky130_fd_sc_hd__a21o_2 _27988_ (.A1(_05943_),
    .A2(_05953_),
    .B1(_05972_),
    .X(_05973_));
 sky130_fd_sc_hd__nand3_2 _27989_ (.A(_05943_),
    .B(_05953_),
    .C(_05972_),
    .Y(_05974_));
 sky130_fd_sc_hd__nand3_2 _27990_ (.A(_05973_),
    .B(_05819_),
    .C(_05974_),
    .Y(_05975_));
 sky130_fd_sc_hd__a21oi_2 _27991_ (.A1(_05943_),
    .A2(_05953_),
    .B1(_05972_),
    .Y(_05976_));
 sky130_fd_sc_hd__o211a_2 _27992_ (.A1(_05968_),
    .A2(_05971_),
    .B1(_05953_),
    .C1(_05943_),
    .X(_05977_));
 sky130_fd_sc_hd__o22ai_2 _27993_ (.A1(_05811_),
    .A2(_05798_),
    .B1(_05976_),
    .B2(_05977_),
    .Y(_05978_));
 sky130_fd_sc_hd__and2_2 _27994_ (.A(_05790_),
    .B(_05749_),
    .X(_05979_));
 sky130_fd_sc_hd__inv_2 _27995_ (.A(_05797_),
    .Y(_05980_));
 sky130_fd_sc_hd__nor2_2 _27996_ (.A(_05979_),
    .B(_05980_),
    .Y(_05981_));
 sky130_fd_sc_hd__inv_2 _27997_ (.A(_05979_),
    .Y(_05982_));
 sky130_fd_sc_hd__nor2_2 _27998_ (.A(_05982_),
    .B(_05797_),
    .Y(_05983_));
 sky130_fd_sc_hd__o2bb2ai_2 _27999_ (.A1_N(_05975_),
    .A2_N(_05978_),
    .B1(_05981_),
    .B2(_05983_),
    .Y(_05984_));
 sky130_fd_sc_hd__a21boi_2 _28000_ (.A1(_05820_),
    .A2(_05828_),
    .B1_N(_05815_),
    .Y(_05985_));
 sky130_fd_sc_hd__nor2_2 _28001_ (.A(_05979_),
    .B(_05797_),
    .Y(_05986_));
 sky130_fd_sc_hd__nor2_2 _28002_ (.A(_05982_),
    .B(_05980_),
    .Y(_05987_));
 sky130_fd_sc_hd__nor2_2 _28003_ (.A(_05986_),
    .B(_05987_),
    .Y(_05988_));
 sky130_fd_sc_hd__nand3b_2 _28004_ (.A_N(_05988_),
    .B(_05978_),
    .C(_05975_),
    .Y(_05989_));
 sky130_fd_sc_hd__nand3_2 _28005_ (.A(_05984_),
    .B(_05985_),
    .C(_05989_),
    .Y(_05990_));
 sky130_fd_sc_hd__nand2_2 _28006_ (.A(_05990_),
    .B(_05822_),
    .Y(_05991_));
 sky130_fd_sc_hd__o2bb2ai_2 _28007_ (.A1_N(_05975_),
    .A2_N(_05978_),
    .B1(_05986_),
    .B2(_05987_),
    .Y(_05992_));
 sky130_fd_sc_hd__nand2_2 _28008_ (.A(_05688_),
    .B(_05812_),
    .Y(_05993_));
 sky130_fd_sc_hd__a21oi_2 _28009_ (.A1(_05812_),
    .A2(_05814_),
    .B1(_05688_),
    .Y(_05994_));
 sky130_fd_sc_hd__o22ai_2 _28010_ (.A1(_05819_),
    .A2(_05993_),
    .B1(_05837_),
    .B2(_05994_),
    .Y(_05995_));
 sky130_fd_sc_hd__nand3_2 _28011_ (.A(_05978_),
    .B(_05988_),
    .C(_05975_),
    .Y(_05996_));
 sky130_fd_sc_hd__nand3_2 _28012_ (.A(_05992_),
    .B(_05995_),
    .C(_05996_),
    .Y(_05997_));
 sky130_fd_sc_hd__nand2_2 _28013_ (.A(_05990_),
    .B(_05997_),
    .Y(_05998_));
 sky130_fd_sc_hd__a22oi_2 _28014_ (.A1(_05841_),
    .A2(_05830_),
    .B1(_05998_),
    .B2(_05836_),
    .Y(_05999_));
 sky130_fd_sc_hd__o2bb2ai_2 _28015_ (.A1_N(_05997_),
    .A2_N(_05990_),
    .B1(_05664_),
    .B2(_05821_),
    .Y(_06000_));
 sky130_fd_sc_hd__nand2_2 _28016_ (.A(_05841_),
    .B(_05830_),
    .Y(_06001_));
 sky130_fd_sc_hd__a21oi_2 _28017_ (.A1(_06000_),
    .A2(_05991_),
    .B1(_06001_),
    .Y(_06002_));
 sky130_fd_sc_hd__a21oi_2 _28018_ (.A1(_05991_),
    .A2(_05999_),
    .B1(_06002_),
    .Y(_06003_));
 sky130_fd_sc_hd__o22ai_2 _28019_ (.A1(_05844_),
    .A2(_05845_),
    .B1(_05843_),
    .B2(_05711_),
    .Y(_06004_));
 sky130_fd_sc_hd__xor2_2 _28020_ (.A(_06003_),
    .B(_06004_),
    .X(_02631_));
 sky130_fd_sc_hd__nand2_2 _28021_ (.A(_05978_),
    .B(_05988_),
    .Y(_06005_));
 sky130_fd_sc_hd__nand2_2 _28022_ (.A(_06005_),
    .B(_05975_),
    .Y(_06006_));
 sky130_fd_sc_hd__nand2_2 _28023_ (.A(_05942_),
    .B(_05886_),
    .Y(_06007_));
 sky130_fd_sc_hd__buf_1 _28024_ (.A(\pcpi_mul.rs2[8] ),
    .X(_06008_));
 sky130_fd_sc_hd__nand2_2 _28025_ (.A(_06008_),
    .B(_05340_),
    .Y(_06009_));
 sky130_fd_sc_hd__buf_1 _28026_ (.A(\pcpi_mul.rs2[7] ),
    .X(_06010_));
 sky130_fd_sc_hd__nand2_2 _28027_ (.A(_06010_),
    .B(_05251_),
    .Y(_06011_));
 sky130_fd_sc_hd__nor2_2 _28028_ (.A(_06009_),
    .B(_06011_),
    .Y(_06012_));
 sky130_fd_sc_hd__and2_2 _28029_ (.A(_06009_),
    .B(_06011_),
    .X(_06013_));
 sky130_fd_sc_hd__nand2_2 _28030_ (.A(_19385_),
    .B(_05420_),
    .Y(_06014_));
 sky130_fd_sc_hd__o21ai_2 _28031_ (.A1(_06012_),
    .A2(_06013_),
    .B1(_06014_),
    .Y(_06015_));
 sky130_fd_sc_hd__or2_2 _28032_ (.A(_06009_),
    .B(_06011_),
    .X(_06016_));
 sky130_fd_sc_hd__nand2_2 _28033_ (.A(_06009_),
    .B(_06011_),
    .Y(_06017_));
 sky130_fd_sc_hd__inv_2 _28034_ (.A(_06014_),
    .Y(_06018_));
 sky130_fd_sc_hd__nand3_2 _28035_ (.A(_06016_),
    .B(_06017_),
    .C(_06018_),
    .Y(_06019_));
 sky130_fd_sc_hd__buf_1 _28036_ (.A(_05673_),
    .X(_06020_));
 sky130_fd_sc_hd__a31o_2 _28037_ (.A1(_05961_),
    .A2(_06020_),
    .A3(_19631_),
    .B1(_05960_),
    .X(_06021_));
 sky130_fd_sc_hd__nand3_2 _28038_ (.A(_06015_),
    .B(_06019_),
    .C(_06021_),
    .Y(_06022_));
 sky130_fd_sc_hd__o21ai_2 _28039_ (.A1(_06012_),
    .A2(_06013_),
    .B1(_06018_),
    .Y(_06023_));
 sky130_fd_sc_hd__nand3_2 _28040_ (.A(_06016_),
    .B(_06017_),
    .C(_06014_),
    .Y(_06024_));
 sky130_fd_sc_hd__a21oi_2 _28041_ (.A1(_05954_),
    .A2(_05961_),
    .B1(_05960_),
    .Y(_06025_));
 sky130_fd_sc_hd__nand3_2 _28042_ (.A(_06023_),
    .B(_06024_),
    .C(_06025_),
    .Y(_06026_));
 sky130_fd_sc_hd__o21ai_2 _28043_ (.A1(_05860_),
    .A2(_05859_),
    .B1(_05863_),
    .Y(_06027_));
 sky130_fd_sc_hd__a21oi_2 _28044_ (.A1(_06022_),
    .A2(_06026_),
    .B1(_06027_),
    .Y(_06028_));
 sky130_fd_sc_hd__and3_2 _28045_ (.A(_06022_),
    .B(_06026_),
    .C(_06027_),
    .X(_06029_));
 sky130_fd_sc_hd__o22ai_2 _28046_ (.A1(_05963_),
    .A2(_05970_),
    .B1(_06028_),
    .B2(_06029_),
    .Y(_06030_));
 sky130_fd_sc_hd__a21o_2 _28047_ (.A1(_06022_),
    .A2(_06026_),
    .B1(_06027_),
    .X(_06031_));
 sky130_fd_sc_hd__a21oi_2 _28048_ (.A1(_05962_),
    .A2(_05967_),
    .B1(_05963_),
    .Y(_06032_));
 sky130_fd_sc_hd__nand3_2 _28049_ (.A(_06022_),
    .B(_06026_),
    .C(_06027_),
    .Y(_06033_));
 sky130_fd_sc_hd__nand3_2 _28050_ (.A(_06031_),
    .B(_06032_),
    .C(_06033_),
    .Y(_06034_));
 sky130_fd_sc_hd__inv_2 _28051_ (.A(_05872_),
    .Y(_06035_));
 sky130_fd_sc_hd__o21ai_2 _28052_ (.A1(_05874_),
    .A2(_06035_),
    .B1(_05868_),
    .Y(_06036_));
 sky130_fd_sc_hd__a21oi_2 _28053_ (.A1(_06030_),
    .A2(_06034_),
    .B1(_06036_),
    .Y(_06037_));
 sky130_fd_sc_hd__nand3_2 _28054_ (.A(_06030_),
    .B(_06034_),
    .C(_06036_),
    .Y(_06038_));
 sky130_fd_sc_hd__nand2_2 _28055_ (.A(_06038_),
    .B(_05888_),
    .Y(_06039_));
 sky130_fd_sc_hd__nor2_2 _28056_ (.A(_06037_),
    .B(_06039_),
    .Y(_06040_));
 sky130_fd_sc_hd__inv_2 _28057_ (.A(_05868_),
    .Y(_06041_));
 sky130_fd_sc_hd__nor2_2 _28058_ (.A(_05876_),
    .B(_06041_),
    .Y(_06042_));
 sky130_fd_sc_hd__a21oi_2 _28059_ (.A1(_06031_),
    .A2(_06033_),
    .B1(_06032_),
    .Y(_06043_));
 sky130_fd_sc_hd__inv_2 _28060_ (.A(_06022_),
    .Y(_06044_));
 sky130_fd_sc_hd__nand2_2 _28061_ (.A(_06026_),
    .B(_06027_),
    .Y(_06045_));
 sky130_fd_sc_hd__o211a_2 _28062_ (.A1(_06044_),
    .A2(_06045_),
    .B1(_06032_),
    .C1(_06031_),
    .X(_06046_));
 sky130_fd_sc_hd__o22ai_2 _28063_ (.A1(_06035_),
    .A2(_06042_),
    .B1(_06043_),
    .B2(_06046_),
    .Y(_06047_));
 sky130_fd_sc_hd__a21oi_2 _28064_ (.A1(_06047_),
    .A2(_06038_),
    .B1(_05888_),
    .Y(_06048_));
 sky130_fd_sc_hd__nor2_2 _28065_ (.A(_05913_),
    .B(_05921_),
    .Y(_06049_));
 sky130_fd_sc_hd__nor2_2 _28066_ (.A(_05898_),
    .B(_05894_),
    .Y(_06050_));
 sky130_fd_sc_hd__buf_1 _28067_ (.A(_05180_),
    .X(_06051_));
 sky130_fd_sc_hd__buf_1 _28068_ (.A(_05408_),
    .X(_06052_));
 sky130_fd_sc_hd__nand2_2 _28069_ (.A(_06051_),
    .B(_06052_),
    .Y(_06053_));
 sky130_fd_sc_hd__buf_1 _28070_ (.A(_05322_),
    .X(_06054_));
 sky130_fd_sc_hd__nand2_2 _28071_ (.A(_06054_),
    .B(_05615_),
    .Y(_06055_));
 sky130_fd_sc_hd__nor2_2 _28072_ (.A(_06053_),
    .B(_06055_),
    .Y(_06056_));
 sky130_fd_sc_hd__buf_1 _28073_ (.A(_05157_),
    .X(_06057_));
 sky130_fd_sc_hd__buf_1 _28074_ (.A(\pcpi_mul.rs1[13] ),
    .X(_06058_));
 sky130_fd_sc_hd__buf_1 _28075_ (.A(_06058_),
    .X(_06059_));
 sky130_fd_sc_hd__nand2_2 _28076_ (.A(_06057_),
    .B(_06059_),
    .Y(_06060_));
 sky130_fd_sc_hd__inv_2 _28077_ (.A(_06060_),
    .Y(_06061_));
 sky130_fd_sc_hd__nand2_2 _28078_ (.A(_06053_),
    .B(_06055_),
    .Y(_06062_));
 sky130_fd_sc_hd__nand2_2 _28079_ (.A(_06061_),
    .B(_06062_),
    .Y(_06063_));
 sky130_fd_sc_hd__and2_2 _28080_ (.A(_06053_),
    .B(_06055_),
    .X(_06064_));
 sky130_fd_sc_hd__o21ai_2 _28081_ (.A1(_06056_),
    .A2(_06064_),
    .B1(_06060_),
    .Y(_06065_));
 sky130_fd_sc_hd__o221ai_2 _28082_ (.A1(_05895_),
    .A2(_06050_),
    .B1(_06056_),
    .B2(_06063_),
    .C1(_06065_),
    .Y(_06066_));
 sky130_fd_sc_hd__o21ai_2 _28083_ (.A1(_06056_),
    .A2(_06064_),
    .B1(_06061_),
    .Y(_06067_));
 sky130_fd_sc_hd__nand3b_2 _28084_ (.A_N(_06056_),
    .B(_06062_),
    .C(_06060_),
    .Y(_06068_));
 sky130_fd_sc_hd__a21oi_2 _28085_ (.A1(_05901_),
    .A2(_05900_),
    .B1(_05895_),
    .Y(_06069_));
 sky130_fd_sc_hd__nand3_2 _28086_ (.A(_06067_),
    .B(_06068_),
    .C(_06069_),
    .Y(_06070_));
 sky130_fd_sc_hd__a22oi_2 _28087_ (.A1(_05141_),
    .A2(_19607_),
    .B1(_05144_),
    .B2(_19604_),
    .Y(_06071_));
 sky130_fd_sc_hd__buf_1 _28088_ (.A(_05122_),
    .X(_06072_));
 sky130_fd_sc_hd__buf_1 _28089_ (.A(_05897_),
    .X(_06073_));
 sky130_fd_sc_hd__buf_1 _28090_ (.A(_19606_),
    .X(_06074_));
 sky130_fd_sc_hd__and4_2 _28091_ (.A(_06072_),
    .B(_19401_),
    .C(_06073_),
    .D(_06074_),
    .X(_06075_));
 sky130_fd_sc_hd__nor2_2 _28092_ (.A(_06071_),
    .B(_06075_),
    .Y(_06076_));
 sky130_fd_sc_hd__nand2_2 _28093_ (.A(_19394_),
    .B(_19610_),
    .Y(_06077_));
 sky130_fd_sc_hd__nand2_2 _28094_ (.A(_06076_),
    .B(_06077_),
    .Y(_06078_));
 sky130_fd_sc_hd__o21bai_2 _28095_ (.A1(_06071_),
    .A2(_06075_),
    .B1_N(_06077_),
    .Y(_06079_));
 sky130_fd_sc_hd__nand2_2 _28096_ (.A(_06078_),
    .B(_06079_),
    .Y(_06080_));
 sky130_fd_sc_hd__a21o_2 _28097_ (.A1(_06066_),
    .A2(_06070_),
    .B1(_06080_),
    .X(_06081_));
 sky130_fd_sc_hd__nand3_2 _28098_ (.A(_06066_),
    .B(_06080_),
    .C(_06070_),
    .Y(_06082_));
 sky130_fd_sc_hd__a21oi_2 _28099_ (.A1(_05902_),
    .A2(_05899_),
    .B1(_05905_),
    .Y(_06083_));
 sky130_fd_sc_hd__o21ai_2 _28100_ (.A1(_06083_),
    .A2(_05919_),
    .B1(_05906_),
    .Y(_06084_));
 sky130_fd_sc_hd__a21oi_2 _28101_ (.A1(_06081_),
    .A2(_06082_),
    .B1(_06084_),
    .Y(_06085_));
 sky130_fd_sc_hd__nor2_2 _28102_ (.A(_06049_),
    .B(_06085_),
    .Y(_06086_));
 sky130_fd_sc_hd__nand3_2 _28103_ (.A(_06084_),
    .B(_06081_),
    .C(_06082_),
    .Y(_06087_));
 sky130_fd_sc_hd__and2_2 _28104_ (.A(_05919_),
    .B(_05906_),
    .X(_06088_));
 sky130_fd_sc_hd__o2bb2ai_2 _28105_ (.A1_N(_06081_),
    .A2_N(_06082_),
    .B1(_06083_),
    .B2(_06088_),
    .Y(_06089_));
 sky130_fd_sc_hd__inv_2 _28106_ (.A(_06049_),
    .Y(_06090_));
 sky130_fd_sc_hd__a21oi_2 _28107_ (.A1(_06089_),
    .A2(_06087_),
    .B1(_06090_),
    .Y(_06091_));
 sky130_fd_sc_hd__a21oi_2 _28108_ (.A1(_06086_),
    .A2(_06087_),
    .B1(_06091_),
    .Y(_06092_));
 sky130_fd_sc_hd__o21ai_2 _28109_ (.A1(_06040_),
    .A2(_06048_),
    .B1(_06092_),
    .Y(_06093_));
 sky130_fd_sc_hd__and3_2 _28110_ (.A(_06030_),
    .B(_06034_),
    .C(_06036_),
    .X(_06094_));
 sky130_fd_sc_hd__o22ai_2 _28111_ (.A1(_05881_),
    .A2(_05878_),
    .B1(_06037_),
    .B2(_06094_),
    .Y(_06095_));
 sky130_fd_sc_hd__nand3_2 _28112_ (.A(_06047_),
    .B(_05888_),
    .C(_06038_),
    .Y(_06096_));
 sky130_fd_sc_hd__a21o_2 _28113_ (.A1(_06089_),
    .A2(_06087_),
    .B1(_06090_),
    .X(_06097_));
 sky130_fd_sc_hd__nand3_2 _28114_ (.A(_06089_),
    .B(_06090_),
    .C(_06087_),
    .Y(_06098_));
 sky130_fd_sc_hd__nand2_2 _28115_ (.A(_06097_),
    .B(_06098_),
    .Y(_06099_));
 sky130_fd_sc_hd__nand3_2 _28116_ (.A(_06095_),
    .B(_06096_),
    .C(_06099_),
    .Y(_06100_));
 sky130_fd_sc_hd__nand3b_2 _28117_ (.A_N(_06007_),
    .B(_06093_),
    .C(_06100_),
    .Y(_06101_));
 sky130_fd_sc_hd__o21ai_2 _28118_ (.A1(_06040_),
    .A2(_06048_),
    .B1(_06099_),
    .Y(_06102_));
 sky130_fd_sc_hd__nand3_2 _28119_ (.A(_06095_),
    .B(_06096_),
    .C(_06092_),
    .Y(_06103_));
 sky130_fd_sc_hd__nand3_2 _28120_ (.A(_06102_),
    .B(_06103_),
    .C(_06007_),
    .Y(_06104_));
 sky130_fd_sc_hd__buf_1 _28121_ (.A(_05849_),
    .X(_06105_));
 sky130_fd_sc_hd__nor2_2 _28122_ (.A(_05497_),
    .B(_06105_),
    .Y(_06106_));
 sky130_fd_sc_hd__nand2_2 _28123_ (.A(_05956_),
    .B(_05119_),
    .Y(_06107_));
 sky130_fd_sc_hd__nand2_2 _28124_ (.A(_05958_),
    .B(_05218_),
    .Y(_06108_));
 sky130_fd_sc_hd__nor2_2 _28125_ (.A(_06107_),
    .B(_06108_),
    .Y(_06109_));
 sky130_fd_sc_hd__nand2_2 _28126_ (.A(_06107_),
    .B(_06108_),
    .Y(_06110_));
 sky130_fd_sc_hd__or3b_2 _28127_ (.A(_06106_),
    .B(_06109_),
    .C_N(_06110_),
    .X(_06111_));
 sky130_fd_sc_hd__or2_2 _28128_ (.A(_06107_),
    .B(_06108_),
    .X(_06112_));
 sky130_fd_sc_hd__inv_2 _28129_ (.A(_06106_),
    .Y(_06113_));
 sky130_fd_sc_hd__a21o_2 _28130_ (.A1(_06112_),
    .A2(_06110_),
    .B1(_06113_),
    .X(_06114_));
 sky130_fd_sc_hd__buf_1 _28131_ (.A(_19365_),
    .X(_06115_));
 sky130_fd_sc_hd__nand2_2 _28132_ (.A(_06115_),
    .B(_05805_),
    .Y(_06116_));
 sky130_fd_sc_hd__buf_1 _28133_ (.A(\pcpi_mul.rs2[12] ),
    .X(_06117_));
 sky130_fd_sc_hd__inv_2 _28134_ (.A(_06117_),
    .Y(_06118_));
 sky130_fd_sc_hd__buf_1 _28135_ (.A(_06118_),
    .X(_06119_));
 sky130_fd_sc_hd__or3_2 _28136_ (.A(_06116_),
    .B(_06119_),
    .C(_05106_),
    .X(_06120_));
 sky130_fd_sc_hd__buf_1 _28137_ (.A(_06118_),
    .X(_06121_));
 sky130_fd_sc_hd__o21ai_2 _28138_ (.A1(_06121_),
    .A2(_05106_),
    .B1(_06116_),
    .Y(_06122_));
 sky130_fd_sc_hd__nand2_2 _28139_ (.A(_06120_),
    .B(_06122_),
    .Y(_06123_));
 sky130_fd_sc_hd__a21oi_2 _28140_ (.A1(_06111_),
    .A2(_06114_),
    .B1(_06123_),
    .Y(_06124_));
 sky130_fd_sc_hd__and3_2 _28141_ (.A(_06111_),
    .B(_06123_),
    .C(_06114_),
    .X(_06125_));
 sky130_fd_sc_hd__or2_2 _28142_ (.A(_06124_),
    .B(_06125_),
    .X(_06126_));
 sky130_fd_sc_hd__inv_2 _28143_ (.A(_06126_),
    .Y(_06127_));
 sky130_fd_sc_hd__a21oi_2 _28144_ (.A1(_06101_),
    .A2(_06104_),
    .B1(_06127_),
    .Y(_06128_));
 sky130_fd_sc_hd__nand3_2 _28145_ (.A(_06101_),
    .B(_06104_),
    .C(_06127_),
    .Y(_06129_));
 sky130_fd_sc_hd__nand2_2 _28146_ (.A(_06129_),
    .B(_05977_),
    .Y(_06130_));
 sky130_fd_sc_hd__nor2_2 _28147_ (.A(_06128_),
    .B(_06130_),
    .Y(_06131_));
 sky130_fd_sc_hd__nand2_2 _28148_ (.A(_06101_),
    .B(_06104_),
    .Y(_06132_));
 sky130_fd_sc_hd__nand2_2 _28149_ (.A(_06132_),
    .B(_06126_),
    .Y(_06133_));
 sky130_fd_sc_hd__a21oi_2 _28150_ (.A1(_06133_),
    .A2(_06129_),
    .B1(_05977_),
    .Y(_06134_));
 sky130_fd_sc_hd__and2_2 _28151_ (.A(_05940_),
    .B(_05924_),
    .X(_06135_));
 sky130_fd_sc_hd__nor2_2 _28152_ (.A(_06135_),
    .B(_05943_),
    .Y(_06136_));
 sky130_fd_sc_hd__and2_2 _28153_ (.A(_05943_),
    .B(_06135_),
    .X(_06137_));
 sky130_fd_sc_hd__or2_2 _28154_ (.A(_06136_),
    .B(_06137_),
    .X(_06138_));
 sky130_fd_sc_hd__inv_2 _28155_ (.A(_06138_),
    .Y(_06139_));
 sky130_fd_sc_hd__o21ai_2 _28156_ (.A1(_06131_),
    .A2(_06134_),
    .B1(_06139_),
    .Y(_06140_));
 sky130_fd_sc_hd__a21o_2 _28157_ (.A1(_06133_),
    .A2(_06129_),
    .B1(_05977_),
    .X(_06141_));
 sky130_fd_sc_hd__a21o_2 _28158_ (.A1(_06126_),
    .A2(_06132_),
    .B1(_06130_),
    .X(_06142_));
 sky130_fd_sc_hd__nand3_2 _28159_ (.A(_06141_),
    .B(_06142_),
    .C(_06138_),
    .Y(_06143_));
 sky130_fd_sc_hd__nand3b_2 _28160_ (.A_N(_06006_),
    .B(_06140_),
    .C(_06143_),
    .Y(_06144_));
 sky130_fd_sc_hd__and2_2 _28161_ (.A(_06144_),
    .B(_05986_),
    .X(_06145_));
 sky130_fd_sc_hd__nand2_2 _28162_ (.A(_06141_),
    .B(_06139_),
    .Y(_06146_));
 sky130_fd_sc_hd__o21ai_2 _28163_ (.A1(_06131_),
    .A2(_06134_),
    .B1(_06138_),
    .Y(_06147_));
 sky130_fd_sc_hd__o211ai_2 _28164_ (.A1(_06131_),
    .A2(_06146_),
    .B1(_06006_),
    .C1(_06147_),
    .Y(_06148_));
 sky130_fd_sc_hd__a21oi_2 _28165_ (.A1(_06148_),
    .A2(_06144_),
    .B1(_05986_),
    .Y(_06149_));
 sky130_fd_sc_hd__nand2_2 _28166_ (.A(_05991_),
    .B(_05997_),
    .Y(_06150_));
 sky130_fd_sc_hd__o21bai_2 _28167_ (.A1(_06145_),
    .A2(_06149_),
    .B1_N(_06150_),
    .Y(_06151_));
 sky130_fd_sc_hd__a21o_2 _28168_ (.A1(_06148_),
    .A2(_06144_),
    .B1(_05986_),
    .X(_06152_));
 sky130_fd_sc_hd__nand2_2 _28169_ (.A(_06144_),
    .B(_05986_),
    .Y(_06153_));
 sky130_fd_sc_hd__nand3_2 _28170_ (.A(_06152_),
    .B(_06153_),
    .C(_06150_),
    .Y(_06154_));
 sky130_fd_sc_hd__nand2_2 _28171_ (.A(_06151_),
    .B(_06154_),
    .Y(_06155_));
 sky130_fd_sc_hd__a22oi_2 _28172_ (.A1(_05991_),
    .A2(_05999_),
    .B1(_06004_),
    .B2(_06003_),
    .Y(_06156_));
 sky130_fd_sc_hd__xor2_2 _28173_ (.A(_06155_),
    .B(_06156_),
    .X(_02632_));
 sky130_fd_sc_hd__a21oi_2 _28174_ (.A1(_06095_),
    .A2(_06092_),
    .B1(_06040_),
    .Y(_06157_));
 sky130_fd_sc_hd__nand2_2 _28175_ (.A(_06008_),
    .B(_05342_),
    .Y(_06158_));
 sky130_fd_sc_hd__nand2_2 _28176_ (.A(_06010_),
    .B(_05502_),
    .Y(_06159_));
 sky130_fd_sc_hd__nor2_2 _28177_ (.A(_06158_),
    .B(_06159_),
    .Y(_06160_));
 sky130_fd_sc_hd__and2_2 _28178_ (.A(_06158_),
    .B(_06159_),
    .X(_06161_));
 sky130_fd_sc_hd__buf_1 _28179_ (.A(\pcpi_mul.rs1[8] ),
    .X(_06162_));
 sky130_fd_sc_hd__nand2_2 _28180_ (.A(_19385_),
    .B(_06162_),
    .Y(_06163_));
 sky130_fd_sc_hd__o21ai_2 _28181_ (.A1(_06160_),
    .A2(_06161_),
    .B1(_06163_),
    .Y(_06164_));
 sky130_fd_sc_hd__a31o_2 _28182_ (.A1(_06110_),
    .A2(_06020_),
    .A3(_19628_),
    .B1(_06109_),
    .X(_06165_));
 sky130_fd_sc_hd__nand2_2 _28183_ (.A(_06158_),
    .B(_06159_),
    .Y(_06166_));
 sky130_fd_sc_hd__inv_2 _28184_ (.A(_06163_),
    .Y(_06167_));
 sky130_fd_sc_hd__nand3b_2 _28185_ (.A_N(_06160_),
    .B(_06166_),
    .C(_06167_),
    .Y(_06168_));
 sky130_fd_sc_hd__nand3_2 _28186_ (.A(_06164_),
    .B(_06165_),
    .C(_06168_),
    .Y(_06169_));
 sky130_fd_sc_hd__o21ai_2 _28187_ (.A1(_06160_),
    .A2(_06161_),
    .B1(_06167_),
    .Y(_06170_));
 sky130_fd_sc_hd__nand3b_2 _28188_ (.A_N(_06160_),
    .B(_06166_),
    .C(_06163_),
    .Y(_06171_));
 sky130_fd_sc_hd__a21oi_2 _28189_ (.A1(_06106_),
    .A2(_06110_),
    .B1(_06109_),
    .Y(_06172_));
 sky130_fd_sc_hd__nand3_2 _28190_ (.A(_06170_),
    .B(_06171_),
    .C(_06172_),
    .Y(_06173_));
 sky130_fd_sc_hd__nand2_2 _28191_ (.A(_06169_),
    .B(_06173_),
    .Y(_06174_));
 sky130_fd_sc_hd__a21oi_2 _28192_ (.A1(_06018_),
    .A2(_06017_),
    .B1(_06012_),
    .Y(_06175_));
 sky130_fd_sc_hd__nand2_2 _28193_ (.A(_06174_),
    .B(_06175_),
    .Y(_06176_));
 sky130_fd_sc_hd__inv_2 _28194_ (.A(_06175_),
    .Y(_06177_));
 sky130_fd_sc_hd__nand3_2 _28195_ (.A(_06169_),
    .B(_06173_),
    .C(_06177_),
    .Y(_06178_));
 sky130_fd_sc_hd__a21oi_2 _28196_ (.A1(_06176_),
    .A2(_06178_),
    .B1(_06124_),
    .Y(_06179_));
 sky130_fd_sc_hd__nand2_2 _28197_ (.A(_06173_),
    .B(_06177_),
    .Y(_06180_));
 sky130_fd_sc_hd__inv_2 _28198_ (.A(_06169_),
    .Y(_06181_));
 sky130_fd_sc_hd__o211a_2 _28199_ (.A1(_06180_),
    .A2(_06181_),
    .B1(_06124_),
    .C1(_06176_),
    .X(_06182_));
 sky130_fd_sc_hd__nand2_2 _28200_ (.A(_06045_),
    .B(_06022_),
    .Y(_06183_));
 sky130_fd_sc_hd__o21ai_2 _28201_ (.A1(_06179_),
    .A2(_06182_),
    .B1(_06183_),
    .Y(_06184_));
 sky130_fd_sc_hd__a21oi_2 _28202_ (.A1(_06030_),
    .A2(_06036_),
    .B1(_06046_),
    .Y(_06185_));
 sky130_fd_sc_hd__a21o_2 _28203_ (.A1(_06176_),
    .A2(_06178_),
    .B1(_06124_),
    .X(_06186_));
 sky130_fd_sc_hd__nand3_2 _28204_ (.A(_06176_),
    .B(_06124_),
    .C(_06178_),
    .Y(_06187_));
 sky130_fd_sc_hd__inv_2 _28205_ (.A(_06183_),
    .Y(_06188_));
 sky130_fd_sc_hd__nand3_2 _28206_ (.A(_06186_),
    .B(_06187_),
    .C(_06188_),
    .Y(_06189_));
 sky130_fd_sc_hd__nand3_2 _28207_ (.A(_06184_),
    .B(_06185_),
    .C(_06189_),
    .Y(_06190_));
 sky130_fd_sc_hd__a21oi_2 _28208_ (.A1(_05872_),
    .A2(_05876_),
    .B1(_06041_),
    .Y(_06191_));
 sky130_fd_sc_hd__o21ai_2 _28209_ (.A1(_06191_),
    .A2(_06043_),
    .B1(_06034_),
    .Y(_06192_));
 sky130_fd_sc_hd__inv_2 _28210_ (.A(_06026_),
    .Y(_06193_));
 sky130_fd_sc_hd__nor2_2 _28211_ (.A(_06027_),
    .B(_06044_),
    .Y(_06194_));
 sky130_fd_sc_hd__o22ai_2 _28212_ (.A1(_06193_),
    .A2(_06194_),
    .B1(_06179_),
    .B2(_06182_),
    .Y(_06195_));
 sky130_fd_sc_hd__nand3_2 _28213_ (.A(_06186_),
    .B(_06187_),
    .C(_06183_),
    .Y(_06196_));
 sky130_fd_sc_hd__nand3_2 _28214_ (.A(_06192_),
    .B(_06195_),
    .C(_06196_),
    .Y(_06197_));
 sky130_fd_sc_hd__nand2_2 _28215_ (.A(_06190_),
    .B(_06197_),
    .Y(_06198_));
 sky130_fd_sc_hd__buf_1 _28216_ (.A(_05180_),
    .X(_06199_));
 sky130_fd_sc_hd__nand2_2 _28217_ (.A(_06199_),
    .B(_05615_),
    .Y(_06200_));
 sky130_fd_sc_hd__buf_1 _28218_ (.A(_05155_),
    .X(_06201_));
 sky130_fd_sc_hd__nand2_2 _28219_ (.A(_06201_),
    .B(_19609_),
    .Y(_06202_));
 sky130_fd_sc_hd__nor2_2 _28220_ (.A(_06200_),
    .B(_06202_),
    .Y(_06203_));
 sky130_fd_sc_hd__and2_2 _28221_ (.A(_06200_),
    .B(_06202_),
    .X(_06204_));
 sky130_fd_sc_hd__buf_1 _28222_ (.A(\pcpi_mul.rs1[14] ),
    .X(_06205_));
 sky130_fd_sc_hd__buf_1 _28223_ (.A(_06205_),
    .X(_06206_));
 sky130_fd_sc_hd__nand2_2 _28224_ (.A(_06057_),
    .B(_06206_),
    .Y(_06207_));
 sky130_fd_sc_hd__inv_2 _28225_ (.A(_06207_),
    .Y(_06208_));
 sky130_fd_sc_hd__o21ai_2 _28226_ (.A1(_06203_),
    .A2(_06204_),
    .B1(_06208_),
    .Y(_06209_));
 sky130_fd_sc_hd__or2_2 _28227_ (.A(_06200_),
    .B(_06202_),
    .X(_06210_));
 sky130_fd_sc_hd__nand2_2 _28228_ (.A(_06200_),
    .B(_06202_),
    .Y(_06211_));
 sky130_fd_sc_hd__nand3_2 _28229_ (.A(_06210_),
    .B(_06211_),
    .C(_06207_),
    .Y(_06212_));
 sky130_fd_sc_hd__a21oi_2 _28230_ (.A1(_06061_),
    .A2(_06062_),
    .B1(_06056_),
    .Y(_06213_));
 sky130_fd_sc_hd__nand3_2 _28231_ (.A(_06209_),
    .B(_06212_),
    .C(_06213_),
    .Y(_06214_));
 sky130_fd_sc_hd__o21ai_2 _28232_ (.A1(_06203_),
    .A2(_06204_),
    .B1(_06207_),
    .Y(_06215_));
 sky130_fd_sc_hd__nand3_2 _28233_ (.A(_06210_),
    .B(_06211_),
    .C(_06208_),
    .Y(_06216_));
 sky130_fd_sc_hd__o21ai_2 _28234_ (.A1(_06053_),
    .A2(_06055_),
    .B1(_06063_),
    .Y(_06217_));
 sky130_fd_sc_hd__nand3_2 _28235_ (.A(_06215_),
    .B(_06216_),
    .C(_06217_),
    .Y(_06218_));
 sky130_fd_sc_hd__buf_1 _28236_ (.A(_05268_),
    .X(_06219_));
 sky130_fd_sc_hd__buf_1 _28237_ (.A(_05210_),
    .X(_06220_));
 sky130_fd_sc_hd__a22oi_2 _28238_ (.A1(_06219_),
    .A2(_06073_),
    .B1(_06220_),
    .B2(_19601_),
    .Y(_06221_));
 sky130_fd_sc_hd__buf_1 _28239_ (.A(_19600_),
    .X(_06222_));
 sky130_fd_sc_hd__and4_2 _28240_ (.A(_06219_),
    .B(_06220_),
    .C(_06222_),
    .D(_06073_),
    .X(_06223_));
 sky130_fd_sc_hd__inv_2 _28241_ (.A(_19605_),
    .Y(_06224_));
 sky130_fd_sc_hd__buf_1 _28242_ (.A(_06224_),
    .X(_06225_));
 sky130_fd_sc_hd__nor2_2 _28243_ (.A(_05150_),
    .B(_06225_),
    .Y(_06226_));
 sky130_fd_sc_hd__o21bai_2 _28244_ (.A1(_06221_),
    .A2(_06223_),
    .B1_N(_06226_),
    .Y(_06227_));
 sky130_fd_sc_hd__inv_2 _28245_ (.A(_06227_),
    .Y(_06228_));
 sky130_fd_sc_hd__inv_2 _28246_ (.A(_06221_),
    .Y(_06229_));
 sky130_fd_sc_hd__nand3b_2 _28247_ (.A_N(_06223_),
    .B(_06229_),
    .C(_06226_),
    .Y(_06230_));
 sky130_fd_sc_hd__inv_2 _28248_ (.A(_06230_),
    .Y(_06231_));
 sky130_fd_sc_hd__o2bb2ai_2 _28249_ (.A1_N(_06214_),
    .A2_N(_06218_),
    .B1(_06228_),
    .B2(_06231_),
    .Y(_06232_));
 sky130_fd_sc_hd__nand2_2 _28250_ (.A(_06230_),
    .B(_06227_),
    .Y(_06233_));
 sky130_fd_sc_hd__nand3b_2 _28251_ (.A_N(_06233_),
    .B(_06218_),
    .C(_06214_),
    .Y(_06234_));
 sky130_fd_sc_hd__nand2_2 _28252_ (.A(_06232_),
    .B(_06234_),
    .Y(_06235_));
 sky130_fd_sc_hd__a21boi_2 _28253_ (.A1(_06070_),
    .A2(_06080_),
    .B1_N(_06066_),
    .Y(_06236_));
 sky130_fd_sc_hd__nand2_2 _28254_ (.A(_06235_),
    .B(_06236_),
    .Y(_06237_));
 sky130_fd_sc_hd__nand2_2 _28255_ (.A(_06082_),
    .B(_06066_),
    .Y(_06238_));
 sky130_fd_sc_hd__nand3_2 _28256_ (.A(_06238_),
    .B(_06232_),
    .C(_06234_),
    .Y(_06239_));
 sky130_fd_sc_hd__a31o_2 _28257_ (.A1(_06076_),
    .A2(_19395_),
    .A3(_19610_),
    .B1(_06075_),
    .X(_06240_));
 sky130_fd_sc_hd__a21oi_2 _28258_ (.A1(_06237_),
    .A2(_06239_),
    .B1(_06240_),
    .Y(_06241_));
 sky130_fd_sc_hd__a21oi_2 _28259_ (.A1(_06232_),
    .A2(_06234_),
    .B1(_06238_),
    .Y(_06242_));
 sky130_fd_sc_hd__nand2_2 _28260_ (.A(_06239_),
    .B(_06240_),
    .Y(_06243_));
 sky130_fd_sc_hd__nor2_2 _28261_ (.A(_06242_),
    .B(_06243_),
    .Y(_06244_));
 sky130_fd_sc_hd__nor2_2 _28262_ (.A(_06241_),
    .B(_06244_),
    .Y(_06245_));
 sky130_fd_sc_hd__nand2_2 _28263_ (.A(_06198_),
    .B(_06245_),
    .Y(_06246_));
 sky130_fd_sc_hd__a21o_2 _28264_ (.A1(_06237_),
    .A2(_06239_),
    .B1(_06240_),
    .X(_06247_));
 sky130_fd_sc_hd__o21ai_2 _28265_ (.A1(_06242_),
    .A2(_06243_),
    .B1(_06247_),
    .Y(_06248_));
 sky130_fd_sc_hd__nand3_2 _28266_ (.A(_06248_),
    .B(_06190_),
    .C(_06197_),
    .Y(_06249_));
 sky130_fd_sc_hd__nand3_2 _28267_ (.A(_06157_),
    .B(_06246_),
    .C(_06249_),
    .Y(_06250_));
 sky130_fd_sc_hd__o22ai_2 _28268_ (.A1(_06037_),
    .A2(_06039_),
    .B1(_06099_),
    .B2(_06048_),
    .Y(_06251_));
 sky130_fd_sc_hd__o2bb2ai_2 _28269_ (.A1_N(_06190_),
    .A2_N(_06197_),
    .B1(_06241_),
    .B2(_06244_),
    .Y(_06252_));
 sky130_fd_sc_hd__nand3_2 _28270_ (.A(_06245_),
    .B(_06190_),
    .C(_06197_),
    .Y(_06253_));
 sky130_fd_sc_hd__nand3_2 _28271_ (.A(_06251_),
    .B(_06252_),
    .C(_06253_),
    .Y(_06254_));
 sky130_fd_sc_hd__nand2_2 _28272_ (.A(_06250_),
    .B(_06254_),
    .Y(_06255_));
 sky130_fd_sc_hd__buf_1 _28273_ (.A(_05955_),
    .X(_06256_));
 sky130_fd_sc_hd__nand2_2 _28274_ (.A(_06256_),
    .B(_19630_),
    .Y(_06257_));
 sky130_fd_sc_hd__buf_1 _28275_ (.A(_19372_),
    .X(_06258_));
 sky130_fd_sc_hd__nand2_2 _28276_ (.A(_06258_),
    .B(_05212_),
    .Y(_06259_));
 sky130_fd_sc_hd__nor2_2 _28277_ (.A(_06257_),
    .B(_06259_),
    .Y(_06260_));
 sky130_fd_sc_hd__nand2_2 _28278_ (.A(_06257_),
    .B(_06259_),
    .Y(_06261_));
 sky130_fd_sc_hd__inv_2 _28279_ (.A(_06261_),
    .Y(_06262_));
 sky130_fd_sc_hd__nand2_2 _28280_ (.A(_05673_),
    .B(_05194_),
    .Y(_06263_));
 sky130_fd_sc_hd__inv_2 _28281_ (.A(_06263_),
    .Y(_06264_));
 sky130_fd_sc_hd__o21ai_2 _28282_ (.A1(_06260_),
    .A2(_06262_),
    .B1(_06264_),
    .Y(_06265_));
 sky130_fd_sc_hd__nand3b_2 _28283_ (.A_N(_06260_),
    .B(_06263_),
    .C(_06261_),
    .Y(_06266_));
 sky130_fd_sc_hd__nand2_2 _28284_ (.A(_06265_),
    .B(_06266_),
    .Y(_06267_));
 sky130_fd_sc_hd__nor2_2 _28285_ (.A(_06121_),
    .B(_05101_),
    .Y(_06268_));
 sky130_fd_sc_hd__buf_1 _28286_ (.A(\pcpi_mul.rs2[14] ),
    .X(_06269_));
 sky130_fd_sc_hd__buf_1 _28287_ (.A(_06269_),
    .X(_06270_));
 sky130_fd_sc_hd__buf_1 _28288_ (.A(_06270_),
    .X(_06271_));
 sky130_fd_sc_hd__buf_1 _28289_ (.A(\pcpi_mul.rs2[13] ),
    .X(_06272_));
 sky130_fd_sc_hd__buf_1 _28290_ (.A(_06272_),
    .X(_06273_));
 sky130_fd_sc_hd__a22oi_2 _28291_ (.A1(_06271_),
    .A2(_05805_),
    .B1(_06273_),
    .B2(_05124_),
    .Y(_06274_));
 sky130_fd_sc_hd__buf_1 _28292_ (.A(\pcpi_mul.rs2[13] ),
    .X(_06275_));
 sky130_fd_sc_hd__buf_1 _28293_ (.A(_06275_),
    .X(_06276_));
 sky130_fd_sc_hd__nand2_2 _28294_ (.A(_06276_),
    .B(_05804_),
    .Y(_06277_));
 sky130_fd_sc_hd__buf_1 _28295_ (.A(_19362_),
    .X(_06278_));
 sky130_fd_sc_hd__nand2_2 _28296_ (.A(_06278_),
    .B(_19640_),
    .Y(_06279_));
 sky130_fd_sc_hd__nor2_2 _28297_ (.A(_06277_),
    .B(_06279_),
    .Y(_06280_));
 sky130_fd_sc_hd__nor2_2 _28298_ (.A(_06274_),
    .B(_06280_),
    .Y(_06281_));
 sky130_fd_sc_hd__nor2_2 _28299_ (.A(_06268_),
    .B(_06281_),
    .Y(_06282_));
 sky130_fd_sc_hd__a21o_2 _28300_ (.A1(_06268_),
    .A2(_06281_),
    .B1(_06120_),
    .X(_06283_));
 sky130_fd_sc_hd__o21ai_2 _28301_ (.A1(_06121_),
    .A2(_05101_),
    .B1(_06281_),
    .Y(_06284_));
 sky130_fd_sc_hd__o21ai_2 _28302_ (.A1(_06274_),
    .A2(_06280_),
    .B1(_06268_),
    .Y(_06285_));
 sky130_fd_sc_hd__nand3_2 _28303_ (.A(_06284_),
    .B(_06120_),
    .C(_06285_),
    .Y(_06286_));
 sky130_fd_sc_hd__o21ai_2 _28304_ (.A1(_06282_),
    .A2(_06283_),
    .B1(_06286_),
    .Y(_06287_));
 sky130_fd_sc_hd__nor2_2 _28305_ (.A(_06267_),
    .B(_06287_),
    .Y(_06288_));
 sky130_fd_sc_hd__and2_2 _28306_ (.A(_06287_),
    .B(_06267_),
    .X(_06289_));
 sky130_fd_sc_hd__nor2_2 _28307_ (.A(_06288_),
    .B(_06289_),
    .Y(_06290_));
 sky130_fd_sc_hd__a21oi_2 _28308_ (.A1(_06255_),
    .A2(_06290_),
    .B1(_06129_),
    .Y(_06291_));
 sky130_fd_sc_hd__buf_1 _28309_ (.A(_06254_),
    .X(_06292_));
 sky130_fd_sc_hd__inv_2 _28310_ (.A(_06290_),
    .Y(_06293_));
 sky130_fd_sc_hd__nand3_2 _28311_ (.A(_06250_),
    .B(_06292_),
    .C(_06293_),
    .Y(_06294_));
 sky130_fd_sc_hd__nand2_2 _28312_ (.A(_06291_),
    .B(_06294_),
    .Y(_06295_));
 sky130_fd_sc_hd__a21oi_2 _28313_ (.A1(_06250_),
    .A2(_06292_),
    .B1(_06293_),
    .Y(_06296_));
 sky130_fd_sc_hd__o211a_2 _28314_ (.A1(_06288_),
    .A2(_06289_),
    .B1(_06254_),
    .C1(_06250_),
    .X(_06297_));
 sky130_fd_sc_hd__o22ai_2 _28315_ (.A1(_06126_),
    .A2(_06132_),
    .B1(_06296_),
    .B2(_06297_),
    .Y(_06298_));
 sky130_fd_sc_hd__and2_2 _28316_ (.A(_06098_),
    .B(_06087_),
    .X(_06299_));
 sky130_fd_sc_hd__nor2_2 _28317_ (.A(_06299_),
    .B(_06104_),
    .Y(_06300_));
 sky130_fd_sc_hd__and2_2 _28318_ (.A(_06104_),
    .B(_06299_),
    .X(_06301_));
 sky130_fd_sc_hd__nor2_2 _28319_ (.A(_06300_),
    .B(_06301_),
    .Y(_06302_));
 sky130_fd_sc_hd__a21o_2 _28320_ (.A1(_06295_),
    .A2(_06298_),
    .B1(_06302_),
    .X(_06303_));
 sky130_fd_sc_hd__nand3_2 _28321_ (.A(_06295_),
    .B(_06298_),
    .C(_06302_),
    .Y(_06304_));
 sky130_fd_sc_hd__nand2_2 _28322_ (.A(_06146_),
    .B(_06142_),
    .Y(_06305_));
 sky130_fd_sc_hd__a21o_2 _28323_ (.A1(_06303_),
    .A2(_06304_),
    .B1(_06305_),
    .X(_06306_));
 sky130_fd_sc_hd__nand3_2 _28324_ (.A(_06305_),
    .B(_06303_),
    .C(_06304_),
    .Y(_06307_));
 sky130_fd_sc_hd__a21o_2 _28325_ (.A1(_06306_),
    .A2(_06307_),
    .B1(_06136_),
    .X(_06308_));
 sky130_fd_sc_hd__nand2_2 _28326_ (.A(_06153_),
    .B(_06148_),
    .Y(_06309_));
 sky130_fd_sc_hd__and2_2 _28327_ (.A(_06308_),
    .B(_06309_),
    .X(_06310_));
 sky130_fd_sc_hd__nand2_2 _28328_ (.A(_06306_),
    .B(_06136_),
    .Y(_06311_));
 sky130_fd_sc_hd__a21oi_2 _28329_ (.A1(_06308_),
    .A2(_06311_),
    .B1(_06309_),
    .Y(_06312_));
 sky130_fd_sc_hd__a21oi_2 _28330_ (.A1(_06310_),
    .A2(_06311_),
    .B1(_06312_),
    .Y(_06313_));
 sky130_fd_sc_hd__nand2_2 _28331_ (.A(_06152_),
    .B(_06150_),
    .Y(_06314_));
 sky130_fd_sc_hd__o22ai_2 _28332_ (.A1(_06145_),
    .A2(_06314_),
    .B1(_06155_),
    .B2(_06156_),
    .Y(_06315_));
 sky130_fd_sc_hd__or2_2 _28333_ (.A(_06313_),
    .B(_06315_),
    .X(_06316_));
 sky130_fd_sc_hd__nand2_2 _28334_ (.A(_06315_),
    .B(_06313_),
    .Y(_06317_));
 sky130_fd_sc_hd__and2_2 _28335_ (.A(_06316_),
    .B(_06317_),
    .X(_02633_));
 sky130_fd_sc_hd__nand2_2 _28336_ (.A(_06311_),
    .B(_06307_),
    .Y(_06318_));
 sky130_fd_sc_hd__o21a_2 _28337_ (.A1(_06242_),
    .A2(_06243_),
    .B1(_06239_),
    .X(_06319_));
 sky130_fd_sc_hd__and2b_2 _28338_ (.A_N(_06319_),
    .B(_06292_),
    .X(_06320_));
 sky130_fd_sc_hd__and2b_2 _28339_ (.A_N(_06292_),
    .B(_06319_),
    .X(_06321_));
 sky130_fd_sc_hd__a21boi_2 _28340_ (.A1(_06245_),
    .A2(_06190_),
    .B1_N(_06197_),
    .Y(_06322_));
 sky130_fd_sc_hd__nand2_2 _28341_ (.A(_05758_),
    .B(_05420_),
    .Y(_06323_));
 sky130_fd_sc_hd__nand2_2 _28342_ (.A(_05760_),
    .B(_05506_),
    .Y(_06324_));
 sky130_fd_sc_hd__nor2_2 _28343_ (.A(_06323_),
    .B(_06324_),
    .Y(_06325_));
 sky130_fd_sc_hd__nand2_2 _28344_ (.A(_06323_),
    .B(_06324_),
    .Y(_06326_));
 sky130_fd_sc_hd__buf_1 _28345_ (.A(_19612_),
    .X(_06327_));
 sky130_fd_sc_hd__nand2_2 _28346_ (.A(_19385_),
    .B(_06327_),
    .Y(_06328_));
 sky130_fd_sc_hd__inv_2 _28347_ (.A(_06328_),
    .Y(_06329_));
 sky130_fd_sc_hd__nand3b_2 _28348_ (.A_N(_06325_),
    .B(_06326_),
    .C(_06329_),
    .Y(_06330_));
 sky130_fd_sc_hd__a21o_2 _28349_ (.A1(_06264_),
    .A2(_06261_),
    .B1(_06260_),
    .X(_06331_));
 sky130_fd_sc_hd__inv_2 _28350_ (.A(_05419_),
    .Y(_06332_));
 sky130_fd_sc_hd__buf_1 _28351_ (.A(_06332_),
    .X(_06333_));
 sky130_fd_sc_hd__buf_1 _28352_ (.A(\pcpi_mul.rs2[7] ),
    .X(_06334_));
 sky130_fd_sc_hd__nand3_2 _28353_ (.A(_19379_),
    .B(_06334_),
    .C(_19615_),
    .Y(_06335_));
 sky130_fd_sc_hd__o21ai_2 _28354_ (.A1(_06333_),
    .A2(_06335_),
    .B1(_06326_),
    .Y(_06336_));
 sky130_fd_sc_hd__nand2_2 _28355_ (.A(_06336_),
    .B(_06328_),
    .Y(_06337_));
 sky130_fd_sc_hd__nand3_2 _28356_ (.A(_06330_),
    .B(_06331_),
    .C(_06337_),
    .Y(_06338_));
 sky130_fd_sc_hd__nand3b_2 _28357_ (.A_N(_06325_),
    .B(_06326_),
    .C(_06328_),
    .Y(_06339_));
 sky130_fd_sc_hd__a21oi_2 _28358_ (.A1(_06264_),
    .A2(_06261_),
    .B1(_06260_),
    .Y(_06340_));
 sky130_fd_sc_hd__nand2_2 _28359_ (.A(_06336_),
    .B(_06329_),
    .Y(_06341_));
 sky130_fd_sc_hd__nand3_2 _28360_ (.A(_06339_),
    .B(_06340_),
    .C(_06341_),
    .Y(_06342_));
 sky130_fd_sc_hd__a21o_2 _28361_ (.A1(_06167_),
    .A2(_06166_),
    .B1(_06160_),
    .X(_06343_));
 sky130_fd_sc_hd__a21o_2 _28362_ (.A1(_06338_),
    .A2(_06342_),
    .B1(_06343_),
    .X(_06344_));
 sky130_fd_sc_hd__nand3_2 _28363_ (.A(_06338_),
    .B(_06342_),
    .C(_06343_),
    .Y(_06345_));
 sky130_fd_sc_hd__o2bb2ai_2 _28364_ (.A1_N(_06286_),
    .A2_N(_06267_),
    .B1(_06282_),
    .B2(_06283_),
    .Y(_06346_));
 sky130_fd_sc_hd__a21oi_2 _28365_ (.A1(_06344_),
    .A2(_06345_),
    .B1(_06346_),
    .Y(_06347_));
 sky130_fd_sc_hd__inv_2 _28366_ (.A(_06338_),
    .Y(_06348_));
 sky130_fd_sc_hd__nand2_2 _28367_ (.A(_06342_),
    .B(_06343_),
    .Y(_06349_));
 sky130_fd_sc_hd__o211a_2 _28368_ (.A1(_06348_),
    .A2(_06349_),
    .B1(_06344_),
    .C1(_06346_),
    .X(_06350_));
 sky130_fd_sc_hd__nand2_2 _28369_ (.A(_06180_),
    .B(_06169_),
    .Y(_06351_));
 sky130_fd_sc_hd__inv_2 _28370_ (.A(_06351_),
    .Y(_06352_));
 sky130_fd_sc_hd__o21ai_2 _28371_ (.A1(_06347_),
    .A2(_06350_),
    .B1(_06352_),
    .Y(_06353_));
 sky130_fd_sc_hd__o21ai_2 _28372_ (.A1(_06188_),
    .A2(_06179_),
    .B1(_06187_),
    .Y(_06354_));
 sky130_fd_sc_hd__a21o_2 _28373_ (.A1(_06344_),
    .A2(_06345_),
    .B1(_06346_),
    .X(_06355_));
 sky130_fd_sc_hd__nand3_2 _28374_ (.A(_06346_),
    .B(_06344_),
    .C(_06345_),
    .Y(_06356_));
 sky130_fd_sc_hd__nand3_2 _28375_ (.A(_06355_),
    .B(_06351_),
    .C(_06356_),
    .Y(_06357_));
 sky130_fd_sc_hd__nand3_2 _28376_ (.A(_06353_),
    .B(_06354_),
    .C(_06357_),
    .Y(_06358_));
 sky130_fd_sc_hd__and2_2 _28377_ (.A(_06173_),
    .B(_06177_),
    .X(_06359_));
 sky130_fd_sc_hd__o22ai_2 _28378_ (.A1(_06181_),
    .A2(_06359_),
    .B1(_06347_),
    .B2(_06350_),
    .Y(_06360_));
 sky130_fd_sc_hd__nand2_2 _28379_ (.A(_06187_),
    .B(_06188_),
    .Y(_06361_));
 sky130_fd_sc_hd__nand2_2 _28380_ (.A(_06361_),
    .B(_06186_),
    .Y(_06362_));
 sky130_fd_sc_hd__nand3_2 _28381_ (.A(_06355_),
    .B(_06352_),
    .C(_06356_),
    .Y(_06363_));
 sky130_fd_sc_hd__nand3_2 _28382_ (.A(_06360_),
    .B(_06362_),
    .C(_06363_),
    .Y(_06364_));
 sky130_fd_sc_hd__nand2_2 _28383_ (.A(_06358_),
    .B(_06364_),
    .Y(_06365_));
 sky130_fd_sc_hd__and3_2 _28384_ (.A(_06209_),
    .B(_06212_),
    .C(_06213_),
    .X(_06366_));
 sky130_fd_sc_hd__o21ai_2 _28385_ (.A1(_06233_),
    .A2(_06366_),
    .B1(_06218_),
    .Y(_06367_));
 sky130_fd_sc_hd__nand2_2 _28386_ (.A(_19388_),
    .B(_05733_),
    .Y(_06368_));
 sky130_fd_sc_hd__buf_1 _28387_ (.A(\pcpi_mul.rs1[11] ),
    .X(_06369_));
 sky130_fd_sc_hd__nand2_2 _28388_ (.A(_05891_),
    .B(_06369_),
    .Y(_06370_));
 sky130_fd_sc_hd__nor2_2 _28389_ (.A(_06368_),
    .B(_06370_),
    .Y(_06371_));
 sky130_fd_sc_hd__buf_1 _28390_ (.A(\pcpi_mul.rs1[15] ),
    .X(_06372_));
 sky130_fd_sc_hd__buf_1 _28391_ (.A(_06372_),
    .X(_06373_));
 sky130_fd_sc_hd__nand2_2 _28392_ (.A(_19403_),
    .B(_06373_),
    .Y(_06374_));
 sky130_fd_sc_hd__inv_2 _28393_ (.A(_06374_),
    .Y(_06375_));
 sky130_fd_sc_hd__nand2_2 _28394_ (.A(_06368_),
    .B(_06370_),
    .Y(_06376_));
 sky130_fd_sc_hd__nand2_2 _28395_ (.A(_06375_),
    .B(_06376_),
    .Y(_06377_));
 sky130_fd_sc_hd__a21o_2 _28396_ (.A1(_06208_),
    .A2(_06211_),
    .B1(_06203_),
    .X(_06378_));
 sky130_fd_sc_hd__and2_2 _28397_ (.A(_06368_),
    .B(_06370_),
    .X(_06379_));
 sky130_fd_sc_hd__o21ai_2 _28398_ (.A1(_06371_),
    .A2(_06379_),
    .B1(_06374_),
    .Y(_06380_));
 sky130_fd_sc_hd__o211ai_2 _28399_ (.A1(_06371_),
    .A2(_06377_),
    .B1(_06378_),
    .C1(_06380_),
    .Y(_06381_));
 sky130_fd_sc_hd__o21ai_2 _28400_ (.A1(_06371_),
    .A2(_06379_),
    .B1(_06375_),
    .Y(_06382_));
 sky130_fd_sc_hd__or2_2 _28401_ (.A(_06368_),
    .B(_06370_),
    .X(_06383_));
 sky130_fd_sc_hd__nand3_2 _28402_ (.A(_06383_),
    .B(_06376_),
    .C(_06374_),
    .Y(_06384_));
 sky130_fd_sc_hd__a21oi_2 _28403_ (.A1(_06208_),
    .A2(_06211_),
    .B1(_06203_),
    .Y(_06385_));
 sky130_fd_sc_hd__nand3_2 _28404_ (.A(_06382_),
    .B(_06384_),
    .C(_06385_),
    .Y(_06386_));
 sky130_fd_sc_hd__buf_1 _28405_ (.A(\pcpi_mul.rs1[14] ),
    .X(_06387_));
 sky130_fd_sc_hd__buf_1 _28406_ (.A(_06387_),
    .X(_06388_));
 sky130_fd_sc_hd__and4_2 _28407_ (.A(_06072_),
    .B(_19401_),
    .C(_06388_),
    .D(_06222_),
    .X(_06389_));
 sky130_fd_sc_hd__inv_2 _28408_ (.A(\pcpi_mul.rs1[12] ),
    .Y(_06390_));
 sky130_fd_sc_hd__buf_1 _28409_ (.A(_06390_),
    .X(_06391_));
 sky130_fd_sc_hd__nor2_2 _28410_ (.A(_05150_),
    .B(_06391_),
    .Y(_06392_));
 sky130_fd_sc_hd__inv_2 _28411_ (.A(_06392_),
    .Y(_06393_));
 sky130_fd_sc_hd__inv_2 _28412_ (.A(_05205_),
    .Y(_06394_));
 sky130_fd_sc_hd__inv_2 _28413_ (.A(_06205_),
    .Y(_06395_));
 sky130_fd_sc_hd__buf_1 _28414_ (.A(_06395_),
    .X(_06396_));
 sky130_fd_sc_hd__buf_1 _28415_ (.A(_06396_),
    .X(_06397_));
 sky130_fd_sc_hd__nand2_2 _28416_ (.A(_05141_),
    .B(_06222_),
    .Y(_06398_));
 sky130_fd_sc_hd__o21ai_2 _28417_ (.A1(_06394_),
    .A2(_06397_),
    .B1(_06398_),
    .Y(_06399_));
 sky130_fd_sc_hd__nand3b_2 _28418_ (.A_N(_06389_),
    .B(_06393_),
    .C(_06399_),
    .Y(_06400_));
 sky130_fd_sc_hd__buf_1 _28419_ (.A(_06395_),
    .X(_06401_));
 sky130_fd_sc_hd__o21a_2 _28420_ (.A1(_06394_),
    .A2(_06401_),
    .B1(_06398_),
    .X(_06402_));
 sky130_fd_sc_hd__o21ai_2 _28421_ (.A1(_06389_),
    .A2(_06402_),
    .B1(_06392_),
    .Y(_06403_));
 sky130_fd_sc_hd__nand2_2 _28422_ (.A(_06400_),
    .B(_06403_),
    .Y(_06404_));
 sky130_fd_sc_hd__a21o_2 _28423_ (.A1(_06381_),
    .A2(_06386_),
    .B1(_06404_),
    .X(_06405_));
 sky130_fd_sc_hd__nand3_2 _28424_ (.A(_06404_),
    .B(_06381_),
    .C(_06386_),
    .Y(_06406_));
 sky130_fd_sc_hd__nand3_2 _28425_ (.A(_06367_),
    .B(_06405_),
    .C(_06406_),
    .Y(_06407_));
 sky130_fd_sc_hd__nor2_2 _28426_ (.A(_06223_),
    .B(_06231_),
    .Y(_06408_));
 sky130_fd_sc_hd__a21oi_2 _28427_ (.A1(_06405_),
    .A2(_06406_),
    .B1(_06367_),
    .Y(_06409_));
 sky130_fd_sc_hd__nor2_2 _28428_ (.A(_06408_),
    .B(_06409_),
    .Y(_06410_));
 sky130_fd_sc_hd__and2_2 _28429_ (.A(_06218_),
    .B(_06233_),
    .X(_06411_));
 sky130_fd_sc_hd__o2bb2ai_2 _28430_ (.A1_N(_06405_),
    .A2_N(_06406_),
    .B1(_06366_),
    .B2(_06411_),
    .Y(_06412_));
 sky130_fd_sc_hd__inv_2 _28431_ (.A(_06408_),
    .Y(_06413_));
 sky130_fd_sc_hd__a21oi_2 _28432_ (.A1(_06412_),
    .A2(_06407_),
    .B1(_06413_),
    .Y(_06414_));
 sky130_fd_sc_hd__a21oi_2 _28433_ (.A1(_06407_),
    .A2(_06410_),
    .B1(_06414_),
    .Y(_06415_));
 sky130_fd_sc_hd__nand2_2 _28434_ (.A(_06365_),
    .B(_06415_),
    .Y(_06416_));
 sky130_fd_sc_hd__and3_2 _28435_ (.A(_06412_),
    .B(_06413_),
    .C(_06407_),
    .X(_06417_));
 sky130_fd_sc_hd__o211ai_2 _28436_ (.A1(_06414_),
    .A2(_06417_),
    .B1(_06364_),
    .C1(_06358_),
    .Y(_06418_));
 sky130_fd_sc_hd__nand3_2 _28437_ (.A(_06322_),
    .B(_06416_),
    .C(_06418_),
    .Y(_06419_));
 sky130_fd_sc_hd__inv_2 _28438_ (.A(_06196_),
    .Y(_06420_));
 sky130_fd_sc_hd__nand2_2 _28439_ (.A(_06192_),
    .B(_06195_),
    .Y(_06421_));
 sky130_fd_sc_hd__a21oi_2 _28440_ (.A1(_06195_),
    .A2(_06196_),
    .B1(_06192_),
    .Y(_06422_));
 sky130_fd_sc_hd__o22ai_2 _28441_ (.A1(_06420_),
    .A2(_06421_),
    .B1(_06248_),
    .B2(_06422_),
    .Y(_06423_));
 sky130_fd_sc_hd__o2bb2ai_2 _28442_ (.A1_N(_06364_),
    .A2_N(_06358_),
    .B1(_06414_),
    .B2(_06417_),
    .Y(_06424_));
 sky130_fd_sc_hd__nand3_2 _28443_ (.A(_06415_),
    .B(_06364_),
    .C(_06358_),
    .Y(_06425_));
 sky130_fd_sc_hd__nand3_2 _28444_ (.A(_06423_),
    .B(_06424_),
    .C(_06425_),
    .Y(_06426_));
 sky130_fd_sc_hd__buf_1 _28445_ (.A(_06426_),
    .X(_06427_));
 sky130_fd_sc_hd__nand2_2 _28446_ (.A(_06419_),
    .B(_06427_),
    .Y(_06428_));
 sky130_fd_sc_hd__nand2_2 _28447_ (.A(_19360_),
    .B(_19642_),
    .Y(_06429_));
 sky130_fd_sc_hd__buf_1 _28448_ (.A(\pcpi_mul.rs2[11] ),
    .X(_06430_));
 sky130_fd_sc_hd__nand2_2 _28449_ (.A(_06430_),
    .B(_05158_),
    .Y(_06431_));
 sky130_fd_sc_hd__buf_1 _28450_ (.A(\pcpi_mul.rs2[10] ),
    .X(_06432_));
 sky130_fd_sc_hd__buf_1 _28451_ (.A(_06432_),
    .X(_06433_));
 sky130_fd_sc_hd__nand3b_2 _28452_ (.A_N(_06431_),
    .B(_06433_),
    .C(_05341_),
    .Y(_06434_));
 sky130_fd_sc_hd__nand2_2 _28453_ (.A(_19373_),
    .B(_05194_),
    .Y(_06435_));
 sky130_fd_sc_hd__nand2_2 _28454_ (.A(_06431_),
    .B(_06435_),
    .Y(_06436_));
 sky130_fd_sc_hd__nand2_2 _28455_ (.A(_05673_),
    .B(_05422_),
    .Y(_06437_));
 sky130_fd_sc_hd__a21o_2 _28456_ (.A1(_06434_),
    .A2(_06436_),
    .B1(_06437_),
    .X(_06438_));
 sky130_fd_sc_hd__nand3_2 _28457_ (.A(_06434_),
    .B(_06436_),
    .C(_06437_),
    .Y(_06439_));
 sky130_fd_sc_hd__nand2_2 _28458_ (.A(_06438_),
    .B(_06439_),
    .Y(_06440_));
 sky130_fd_sc_hd__buf_1 _28459_ (.A(_06269_),
    .X(_06441_));
 sky130_fd_sc_hd__nand2_2 _28460_ (.A(_06441_),
    .B(_05543_),
    .Y(_06442_));
 sky130_fd_sc_hd__buf_1 _28461_ (.A(\pcpi_mul.rs2[13] ),
    .X(_06443_));
 sky130_fd_sc_hd__nand2_2 _28462_ (.A(_06443_),
    .B(_05545_),
    .Y(_06444_));
 sky130_fd_sc_hd__nor2_2 _28463_ (.A(_06442_),
    .B(_06444_),
    .Y(_06445_));
 sky130_fd_sc_hd__buf_1 _28464_ (.A(_06117_),
    .X(_06446_));
 sky130_fd_sc_hd__buf_1 _28465_ (.A(_05146_),
    .X(_06447_));
 sky130_fd_sc_hd__nand2_2 _28466_ (.A(_06446_),
    .B(_06447_),
    .Y(_06448_));
 sky130_fd_sc_hd__inv_2 _28467_ (.A(_06448_),
    .Y(_06449_));
 sky130_fd_sc_hd__nand2_2 _28468_ (.A(_06442_),
    .B(_06444_),
    .Y(_06450_));
 sky130_fd_sc_hd__nand2_2 _28469_ (.A(_06449_),
    .B(_06450_),
    .Y(_06451_));
 sky130_fd_sc_hd__nand2_2 _28470_ (.A(_06277_),
    .B(_06279_),
    .Y(_06452_));
 sky130_fd_sc_hd__a31o_2 _28471_ (.A1(_06452_),
    .A2(_19369_),
    .A3(_19634_),
    .B1(_06280_),
    .X(_06453_));
 sky130_fd_sc_hd__and2_2 _28472_ (.A(_06442_),
    .B(_06444_),
    .X(_06454_));
 sky130_fd_sc_hd__o21ai_2 _28473_ (.A1(_06445_),
    .A2(_06454_),
    .B1(_06448_),
    .Y(_06455_));
 sky130_fd_sc_hd__o211ai_2 _28474_ (.A1(_06445_),
    .A2(_06451_),
    .B1(_06453_),
    .C1(_06455_),
    .Y(_06456_));
 sky130_fd_sc_hd__o21ai_2 _28475_ (.A1(_06445_),
    .A2(_06454_),
    .B1(_06449_),
    .Y(_06457_));
 sky130_fd_sc_hd__nand3b_2 _28476_ (.A_N(_06445_),
    .B(_06450_),
    .C(_06448_),
    .Y(_06458_));
 sky130_fd_sc_hd__a21oi_2 _28477_ (.A1(_06268_),
    .A2(_06452_),
    .B1(_06280_),
    .Y(_06459_));
 sky130_fd_sc_hd__nand3_2 _28478_ (.A(_06457_),
    .B(_06458_),
    .C(_06459_),
    .Y(_06460_));
 sky130_fd_sc_hd__nand2_2 _28479_ (.A(_06456_),
    .B(_06460_),
    .Y(_06461_));
 sky130_fd_sc_hd__xor2_2 _28480_ (.A(_06440_),
    .B(_06461_),
    .X(_06462_));
 sky130_fd_sc_hd__nor2_2 _28481_ (.A(_06429_),
    .B(_06462_),
    .Y(_06463_));
 sky130_fd_sc_hd__and2_2 _28482_ (.A(_06462_),
    .B(_06429_),
    .X(_06464_));
 sky130_fd_sc_hd__nor2_2 _28483_ (.A(_06463_),
    .B(_06464_),
    .Y(_06465_));
 sky130_fd_sc_hd__inv_2 _28484_ (.A(_06465_),
    .Y(_06466_));
 sky130_fd_sc_hd__nand2_2 _28485_ (.A(_06428_),
    .B(_06466_),
    .Y(_06467_));
 sky130_fd_sc_hd__nand3_2 _28486_ (.A(_06419_),
    .B(_06427_),
    .C(_06465_),
    .Y(_06468_));
 sky130_fd_sc_hd__a21oi_2 _28487_ (.A1(_06467_),
    .A2(_06468_),
    .B1(_06297_),
    .Y(_06469_));
 sky130_fd_sc_hd__a21oi_2 _28488_ (.A1(_06419_),
    .A2(_06427_),
    .B1(_06465_),
    .Y(_06470_));
 sky130_fd_sc_hd__and3_2 _28489_ (.A(_06419_),
    .B(_06426_),
    .C(_06465_),
    .X(_06471_));
 sky130_fd_sc_hd__nor3_2 _28490_ (.A(_06294_),
    .B(_06470_),
    .C(_06471_),
    .Y(_06472_));
 sky130_fd_sc_hd__o22ai_2 _28491_ (.A1(_06320_),
    .A2(_06321_),
    .B1(_06469_),
    .B2(_06472_),
    .Y(_06473_));
 sky130_fd_sc_hd__o22ai_2 _28492_ (.A1(_06255_),
    .A2(_06290_),
    .B1(_06470_),
    .B2(_06471_),
    .Y(_06474_));
 sky130_fd_sc_hd__nand3_2 _28493_ (.A(_06297_),
    .B(_06467_),
    .C(_06468_),
    .Y(_06475_));
 sky130_fd_sc_hd__nor2_2 _28494_ (.A(_06320_),
    .B(_06321_),
    .Y(_06476_));
 sky130_fd_sc_hd__nand3_2 _28495_ (.A(_06474_),
    .B(_06475_),
    .C(_06476_),
    .Y(_06477_));
 sky130_fd_sc_hd__nand2_2 _28496_ (.A(_06473_),
    .B(_06477_),
    .Y(_06478_));
 sky130_fd_sc_hd__a22o_2 _28497_ (.A1(_06294_),
    .A2(_06291_),
    .B1(_06298_),
    .B2(_06302_),
    .X(_06479_));
 sky130_fd_sc_hd__nand2_2 _28498_ (.A(_06478_),
    .B(_06479_),
    .Y(_06480_));
 sky130_fd_sc_hd__a22oi_2 _28499_ (.A1(_06294_),
    .A2(_06291_),
    .B1(_06298_),
    .B2(_06302_),
    .Y(_06481_));
 sky130_fd_sc_hd__nand3_2 _28500_ (.A(_06473_),
    .B(_06481_),
    .C(_06477_),
    .Y(_06482_));
 sky130_fd_sc_hd__a21o_2 _28501_ (.A1(_06480_),
    .A2(_06482_),
    .B1(_06300_),
    .X(_06483_));
 sky130_fd_sc_hd__nand2_2 _28502_ (.A(_06482_),
    .B(_06300_),
    .Y(_06484_));
 sky130_fd_sc_hd__and2_2 _28503_ (.A(_06483_),
    .B(_06484_),
    .X(_06485_));
 sky130_fd_sc_hd__or2_2 _28504_ (.A(_06318_),
    .B(_06485_),
    .X(_06486_));
 sky130_fd_sc_hd__nand2_2 _28505_ (.A(_06310_),
    .B(_06311_),
    .Y(_06487_));
 sky130_fd_sc_hd__nand2_2 _28506_ (.A(_06317_),
    .B(_06487_),
    .Y(_06488_));
 sky130_fd_sc_hd__nand2_2 _28507_ (.A(_06485_),
    .B(_06318_),
    .Y(_06489_));
 sky130_fd_sc_hd__nand3_2 _28508_ (.A(_06317_),
    .B(_06487_),
    .C(_06489_),
    .Y(_06490_));
 sky130_fd_sc_hd__nand2_2 _28509_ (.A(_06490_),
    .B(_06486_),
    .Y(_06491_));
 sky130_fd_sc_hd__o21a_2 _28510_ (.A1(_06486_),
    .A2(_06488_),
    .B1(_06491_),
    .X(_02634_));
 sky130_fd_sc_hd__buf_1 _28511_ (.A(_19612_),
    .X(_06492_));
 sky130_fd_sc_hd__a22oi_2 _28512_ (.A1(_05542_),
    .A2(_06162_),
    .B1(_19383_),
    .B2(_06492_),
    .Y(_06493_));
 sky130_fd_sc_hd__inv_2 _28513_ (.A(_05516_),
    .Y(_06494_));
 sky130_fd_sc_hd__nor2_2 _28514_ (.A(_06494_),
    .B(_06335_),
    .Y(_06495_));
 sky130_fd_sc_hd__buf_1 _28515_ (.A(\pcpi_mul.rs2[6] ),
    .X(_06496_));
 sky130_fd_sc_hd__buf_1 _28516_ (.A(_05597_),
    .X(_06497_));
 sky130_fd_sc_hd__nand2_2 _28517_ (.A(_06496_),
    .B(_06497_),
    .Y(_06498_));
 sky130_fd_sc_hd__o21ai_2 _28518_ (.A1(_06493_),
    .A2(_06495_),
    .B1(_06498_),
    .Y(_06499_));
 sky130_fd_sc_hd__buf_1 _28519_ (.A(_06430_),
    .X(_06500_));
 sky130_fd_sc_hd__buf_1 _28520_ (.A(_05158_),
    .X(_06501_));
 sky130_fd_sc_hd__buf_1 _28521_ (.A(_05193_),
    .X(_06502_));
 sky130_fd_sc_hd__a22oi_2 _28522_ (.A1(_06500_),
    .A2(_06501_),
    .B1(_06433_),
    .B2(_06502_),
    .Y(_06503_));
 sky130_fd_sc_hd__o21ai_2 _28523_ (.A1(_06437_),
    .A2(_06503_),
    .B1(_06434_),
    .Y(_06504_));
 sky130_fd_sc_hd__buf_1 _28524_ (.A(_06494_),
    .X(_06505_));
 sky130_fd_sc_hd__inv_2 _28525_ (.A(_06498_),
    .Y(_06506_));
 sky130_fd_sc_hd__buf_1 _28526_ (.A(\pcpi_mul.rs1[8] ),
    .X(_06507_));
 sky130_fd_sc_hd__buf_1 _28527_ (.A(_19382_),
    .X(_06508_));
 sky130_fd_sc_hd__a22o_2 _28528_ (.A1(_05851_),
    .A2(_06507_),
    .B1(_06508_),
    .B2(_05734_),
    .X(_06509_));
 sky130_fd_sc_hd__o211ai_2 _28529_ (.A1(_06505_),
    .A2(_06335_),
    .B1(_06506_),
    .C1(_06509_),
    .Y(_06510_));
 sky130_fd_sc_hd__nand3_2 _28530_ (.A(_06499_),
    .B(_06504_),
    .C(_06510_),
    .Y(_06511_));
 sky130_fd_sc_hd__o21ai_2 _28531_ (.A1(_06493_),
    .A2(_06495_),
    .B1(_06506_),
    .Y(_06512_));
 sky130_fd_sc_hd__o21ai_2 _28532_ (.A1(_06431_),
    .A2(_06435_),
    .B1(_06437_),
    .Y(_06513_));
 sky130_fd_sc_hd__nand2_2 _28533_ (.A(_06513_),
    .B(_06436_),
    .Y(_06514_));
 sky130_fd_sc_hd__o211ai_2 _28534_ (.A1(_06505_),
    .A2(_06335_),
    .B1(_06498_),
    .C1(_06509_),
    .Y(_06515_));
 sky130_fd_sc_hd__nand3_2 _28535_ (.A(_06512_),
    .B(_06514_),
    .C(_06515_),
    .Y(_06516_));
 sky130_fd_sc_hd__inv_2 _28536_ (.A(_06326_),
    .Y(_06517_));
 sky130_fd_sc_hd__nor2_2 _28537_ (.A(_06329_),
    .B(_06325_),
    .Y(_06518_));
 sky130_fd_sc_hd__nor2_2 _28538_ (.A(_06517_),
    .B(_06518_),
    .Y(_06519_));
 sky130_fd_sc_hd__nand3_2 _28539_ (.A(_06511_),
    .B(_06516_),
    .C(_06519_),
    .Y(_06520_));
 sky130_fd_sc_hd__o2bb2ai_2 _28540_ (.A1_N(_06511_),
    .A2_N(_06516_),
    .B1(_06517_),
    .B2(_06518_),
    .Y(_06521_));
 sky130_fd_sc_hd__nand2_2 _28541_ (.A(_06440_),
    .B(_06460_),
    .Y(_06522_));
 sky130_fd_sc_hd__nand2_2 _28542_ (.A(_06522_),
    .B(_06456_),
    .Y(_06523_));
 sky130_fd_sc_hd__a21oi_2 _28543_ (.A1(_06520_),
    .A2(_06521_),
    .B1(_06523_),
    .Y(_06524_));
 sky130_fd_sc_hd__a21boi_2 _28544_ (.A1(_06460_),
    .A2(_06440_),
    .B1_N(_06456_),
    .Y(_06525_));
 sky130_fd_sc_hd__nand2_2 _28545_ (.A(_06521_),
    .B(_06520_),
    .Y(_06526_));
 sky130_fd_sc_hd__nor2_2 _28546_ (.A(_06525_),
    .B(_06526_),
    .Y(_06527_));
 sky130_fd_sc_hd__and2_2 _28547_ (.A(_06349_),
    .B(_06338_),
    .X(_06528_));
 sky130_fd_sc_hd__o21ai_2 _28548_ (.A1(_06524_),
    .A2(_06527_),
    .B1(_06528_),
    .Y(_06529_));
 sky130_fd_sc_hd__a21oi_2 _28549_ (.A1(_06526_),
    .A2(_06525_),
    .B1(_06528_),
    .Y(_06530_));
 sky130_fd_sc_hd__nand3_2 _28550_ (.A(_06523_),
    .B(_06520_),
    .C(_06521_),
    .Y(_06531_));
 sky130_fd_sc_hd__nand2_2 _28551_ (.A(_06530_),
    .B(_06531_),
    .Y(_06532_));
 sky130_fd_sc_hd__o21ai_2 _28552_ (.A1(_06352_),
    .A2(_06347_),
    .B1(_06356_),
    .Y(_06533_));
 sky130_fd_sc_hd__a21oi_2 _28553_ (.A1(_06529_),
    .A2(_06532_),
    .B1(_06533_),
    .Y(_06534_));
 sky130_fd_sc_hd__a21o_2 _28554_ (.A1(_06526_),
    .A2(_06525_),
    .B1(_06528_),
    .X(_06535_));
 sky130_fd_sc_hd__o211a_2 _28555_ (.A1(_06527_),
    .A2(_06535_),
    .B1(_06533_),
    .C1(_06529_),
    .X(_06536_));
 sky130_fd_sc_hd__a22oi_2 _28556_ (.A1(_05712_),
    .A2(_06074_),
    .B1(_05892_),
    .B2(_19603_),
    .Y(_06537_));
 sky130_fd_sc_hd__buf_1 _28557_ (.A(_19602_),
    .X(_06538_));
 sky130_fd_sc_hd__buf_1 _28558_ (.A(\pcpi_mul.rs1[11] ),
    .X(_06539_));
 sky130_fd_sc_hd__buf_1 _28559_ (.A(_06539_),
    .X(_06540_));
 sky130_fd_sc_hd__and4_2 _28560_ (.A(_06051_),
    .B(_06201_),
    .C(_06538_),
    .D(_06540_),
    .X(_06541_));
 sky130_fd_sc_hd__buf_1 _28561_ (.A(\pcpi_mul.rs1[16] ),
    .X(_06542_));
 sky130_fd_sc_hd__nand2_2 _28562_ (.A(_19403_),
    .B(_06542_),
    .Y(_06543_));
 sky130_fd_sc_hd__inv_2 _28563_ (.A(_06543_),
    .Y(_06544_));
 sky130_fd_sc_hd__o21ai_2 _28564_ (.A1(_06537_),
    .A2(_06541_),
    .B1(_06544_),
    .Y(_06545_));
 sky130_fd_sc_hd__nand2_2 _28565_ (.A(_06051_),
    .B(_05911_),
    .Y(_06546_));
 sky130_fd_sc_hd__nand3b_2 _28566_ (.A_N(_06546_),
    .B(_19392_),
    .C(_06073_),
    .Y(_06547_));
 sky130_fd_sc_hd__a22o_2 _28567_ (.A1(_05402_),
    .A2(_05911_),
    .B1(_05721_),
    .B2(_19603_),
    .X(_06548_));
 sky130_fd_sc_hd__nand3_2 _28568_ (.A(_06547_),
    .B(_06543_),
    .C(_06548_),
    .Y(_06549_));
 sky130_fd_sc_hd__a21oi_2 _28569_ (.A1(_06375_),
    .A2(_06376_),
    .B1(_06371_),
    .Y(_06550_));
 sky130_fd_sc_hd__a21o_2 _28570_ (.A1(_06545_),
    .A2(_06549_),
    .B1(_06550_),
    .X(_06551_));
 sky130_fd_sc_hd__o21ai_2 _28571_ (.A1(_06537_),
    .A2(_06541_),
    .B1(_06543_),
    .Y(_06552_));
 sky130_fd_sc_hd__nand3_2 _28572_ (.A(_06547_),
    .B(_06544_),
    .C(_06548_),
    .Y(_06553_));
 sky130_fd_sc_hd__nand2_2 _28573_ (.A(_06383_),
    .B(_06377_),
    .Y(_06554_));
 sky130_fd_sc_hd__a21o_2 _28574_ (.A1(_06552_),
    .A2(_06553_),
    .B1(_06554_),
    .X(_06555_));
 sky130_fd_sc_hd__nand2_2 _28575_ (.A(_06551_),
    .B(_06555_),
    .Y(_06556_));
 sky130_fd_sc_hd__buf_1 _28576_ (.A(_19593_),
    .X(_06557_));
 sky130_fd_sc_hd__nand2_2 _28577_ (.A(_05268_),
    .B(_06206_),
    .Y(_06558_));
 sky130_fd_sc_hd__a21o_2 _28578_ (.A1(_05909_),
    .A2(_06557_),
    .B1(_06558_),
    .X(_06559_));
 sky130_fd_sc_hd__buf_1 _28579_ (.A(_06372_),
    .X(_06560_));
 sky130_fd_sc_hd__nand2_2 _28580_ (.A(_05221_),
    .B(_06560_),
    .Y(_06561_));
 sky130_fd_sc_hd__a21o_2 _28581_ (.A1(_05736_),
    .A2(_19597_),
    .B1(_06561_),
    .X(_06562_));
 sky130_fd_sc_hd__nand2_2 _28582_ (.A(_05115_),
    .B(_06222_),
    .Y(_06563_));
 sky130_fd_sc_hd__a21o_2 _28583_ (.A1(_06559_),
    .A2(_06562_),
    .B1(_06563_),
    .X(_06564_));
 sky130_fd_sc_hd__nand3_2 _28584_ (.A(_06559_),
    .B(_06562_),
    .C(_06563_),
    .Y(_06565_));
 sky130_fd_sc_hd__nand2_2 _28585_ (.A(_06564_),
    .B(_06565_),
    .Y(_06566_));
 sky130_fd_sc_hd__inv_2 _28586_ (.A(_06566_),
    .Y(_06567_));
 sky130_fd_sc_hd__nand2_2 _28587_ (.A(_06556_),
    .B(_06567_),
    .Y(_06568_));
 sky130_fd_sc_hd__nand3_2 _28588_ (.A(_06551_),
    .B(_06555_),
    .C(_06566_),
    .Y(_06569_));
 sky130_fd_sc_hd__a21boi_2 _28589_ (.A1(_06404_),
    .A2(_06386_),
    .B1_N(_06381_),
    .Y(_06570_));
 sky130_fd_sc_hd__nand3_2 _28590_ (.A(_06568_),
    .B(_06569_),
    .C(_06570_),
    .Y(_06571_));
 sky130_fd_sc_hd__nor3_2 _28591_ (.A(_06393_),
    .B(_06389_),
    .C(_06402_),
    .Y(_06572_));
 sky130_fd_sc_hd__nor2_2 _28592_ (.A(_06389_),
    .B(_06572_),
    .Y(_06573_));
 sky130_fd_sc_hd__inv_2 _28593_ (.A(_06573_),
    .Y(_06574_));
 sky130_fd_sc_hd__and2_2 _28594_ (.A(_06571_),
    .B(_06574_),
    .X(_06575_));
 sky130_fd_sc_hd__nand2_2 _28595_ (.A(_06556_),
    .B(_06566_),
    .Y(_06576_));
 sky130_fd_sc_hd__nand3_2 _28596_ (.A(_06567_),
    .B(_06551_),
    .C(_06555_),
    .Y(_06577_));
 sky130_fd_sc_hd__nand3b_2 _28597_ (.A_N(_06570_),
    .B(_06576_),
    .C(_06577_),
    .Y(_06578_));
 sky130_fd_sc_hd__a21oi_2 _28598_ (.A1(_06578_),
    .A2(_06571_),
    .B1(_06574_),
    .Y(_06579_));
 sky130_fd_sc_hd__a21oi_2 _28599_ (.A1(_06575_),
    .A2(_06578_),
    .B1(_06579_),
    .Y(_06580_));
 sky130_fd_sc_hd__o21ai_2 _28600_ (.A1(_06534_),
    .A2(_06536_),
    .B1(_06580_),
    .Y(_06581_));
 sky130_fd_sc_hd__a21boi_2 _28601_ (.A1(_06415_),
    .A2(_06364_),
    .B1_N(_06358_),
    .Y(_06582_));
 sky130_fd_sc_hd__a21o_2 _28602_ (.A1(_06575_),
    .A2(_06578_),
    .B1(_06579_),
    .X(_06583_));
 sky130_fd_sc_hd__a21o_2 _28603_ (.A1(_06529_),
    .A2(_06532_),
    .B1(_06533_),
    .X(_06584_));
 sky130_fd_sc_hd__nand3_2 _28604_ (.A(_06529_),
    .B(_06533_),
    .C(_06532_),
    .Y(_06585_));
 sky130_fd_sc_hd__nand3_2 _28605_ (.A(_06583_),
    .B(_06584_),
    .C(_06585_),
    .Y(_06586_));
 sky130_fd_sc_hd__nand3_2 _28606_ (.A(_06581_),
    .B(_06582_),
    .C(_06586_),
    .Y(_06587_));
 sky130_fd_sc_hd__nand2_2 _28607_ (.A(_06578_),
    .B(_06571_),
    .Y(_06588_));
 sky130_fd_sc_hd__nor2_2 _28608_ (.A(_06573_),
    .B(_06588_),
    .Y(_06589_));
 sky130_fd_sc_hd__o22ai_2 _28609_ (.A1(_06589_),
    .A2(_06579_),
    .B1(_06534_),
    .B2(_06536_),
    .Y(_06590_));
 sky130_fd_sc_hd__a21o_2 _28610_ (.A1(_06412_),
    .A2(_06407_),
    .B1(_06413_),
    .X(_06591_));
 sky130_fd_sc_hd__nand2_2 _28611_ (.A(_06410_),
    .B(_06407_),
    .Y(_06592_));
 sky130_fd_sc_hd__nand3_2 _28612_ (.A(_06364_),
    .B(_06591_),
    .C(_06592_),
    .Y(_06593_));
 sky130_fd_sc_hd__nand2_2 _28613_ (.A(_06593_),
    .B(_06358_),
    .Y(_06594_));
 sky130_fd_sc_hd__nand3_2 _28614_ (.A(_06584_),
    .B(_06580_),
    .C(_06585_),
    .Y(_06595_));
 sky130_fd_sc_hd__nand3_2 _28615_ (.A(_06590_),
    .B(_06594_),
    .C(_06595_),
    .Y(_06596_));
 sky130_fd_sc_hd__buf_1 _28616_ (.A(_06596_),
    .X(_06597_));
 sky130_fd_sc_hd__buf_1 _28617_ (.A(_05188_),
    .X(_06598_));
 sky130_fd_sc_hd__nand2_2 _28618_ (.A(_19358_),
    .B(_06598_),
    .Y(_06599_));
 sky130_fd_sc_hd__nand2_2 _28619_ (.A(_19360_),
    .B(_05124_),
    .Y(_06600_));
 sky130_fd_sc_hd__nor2_2 _28620_ (.A(_06599_),
    .B(_06600_),
    .Y(_06601_));
 sky130_fd_sc_hd__inv_2 _28621_ (.A(_06601_),
    .Y(_06602_));
 sky130_fd_sc_hd__nand2_2 _28622_ (.A(_06599_),
    .B(_06600_),
    .Y(_06603_));
 sky130_fd_sc_hd__nand2_2 _28623_ (.A(_06602_),
    .B(_06603_),
    .Y(_06604_));
 sky130_fd_sc_hd__buf_1 _28624_ (.A(_06432_),
    .X(_06605_));
 sky130_fd_sc_hd__buf_1 _28625_ (.A(_19621_),
    .X(_06606_));
 sky130_fd_sc_hd__a22oi_2 _28626_ (.A1(_06500_),
    .A2(_05269_),
    .B1(_06605_),
    .B2(_06606_),
    .Y(_06607_));
 sky130_fd_sc_hd__nand2_2 _28627_ (.A(_05800_),
    .B(_05184_),
    .Y(_06608_));
 sky130_fd_sc_hd__buf_1 _28628_ (.A(_19621_),
    .X(_06609_));
 sky130_fd_sc_hd__nand2_2 _28629_ (.A(_05802_),
    .B(_06609_),
    .Y(_06610_));
 sky130_fd_sc_hd__nor2_2 _28630_ (.A(_06608_),
    .B(_06610_),
    .Y(_06611_));
 sky130_fd_sc_hd__and2_2 _28631_ (.A(_19375_),
    .B(_05502_),
    .X(_06612_));
 sky130_fd_sc_hd__o21ai_2 _28632_ (.A1(_06607_),
    .A2(_06611_),
    .B1(_06612_),
    .Y(_06613_));
 sky130_fd_sc_hd__buf_1 _28633_ (.A(_05342_),
    .X(_06614_));
 sky130_fd_sc_hd__nand3_2 _28634_ (.A(_06500_),
    .B(_06605_),
    .C(_06614_),
    .Y(_06615_));
 sky130_fd_sc_hd__buf_1 _28635_ (.A(_05672_),
    .X(_06616_));
 sky130_fd_sc_hd__buf_1 _28636_ (.A(_05502_),
    .X(_06617_));
 sky130_fd_sc_hd__nand2_2 _28637_ (.A(_06616_),
    .B(_06617_),
    .Y(_06618_));
 sky130_fd_sc_hd__nand2_2 _28638_ (.A(_06608_),
    .B(_06610_),
    .Y(_06619_));
 sky130_fd_sc_hd__o211ai_2 _28639_ (.A1(_05865_),
    .A2(_06615_),
    .B1(_06618_),
    .C1(_06619_),
    .Y(_06620_));
 sky130_fd_sc_hd__nand2_2 _28640_ (.A(_06613_),
    .B(_06620_),
    .Y(_06621_));
 sky130_fd_sc_hd__buf_1 _28641_ (.A(_06447_),
    .X(_06622_));
 sky130_fd_sc_hd__a22oi_2 _28642_ (.A1(_06271_),
    .A2(_05120_),
    .B1(_06273_),
    .B2(_06622_),
    .Y(_06623_));
 sky130_fd_sc_hd__buf_1 _28643_ (.A(\pcpi_mul.rs2[14] ),
    .X(_06624_));
 sky130_fd_sc_hd__nand2_2 _28644_ (.A(_06624_),
    .B(_05119_),
    .Y(_06625_));
 sky130_fd_sc_hd__nand2_2 _28645_ (.A(_06443_),
    .B(_05213_),
    .Y(_06626_));
 sky130_fd_sc_hd__nor2_2 _28646_ (.A(_06625_),
    .B(_06626_),
    .Y(_06627_));
 sky130_fd_sc_hd__buf_1 _28647_ (.A(_19367_),
    .X(_06628_));
 sky130_fd_sc_hd__buf_1 _28648_ (.A(_05211_),
    .X(_06629_));
 sky130_fd_sc_hd__nand2_2 _28649_ (.A(_06628_),
    .B(_06629_),
    .Y(_06630_));
 sky130_fd_sc_hd__o21bai_2 _28650_ (.A1(_06623_),
    .A2(_06627_),
    .B1_N(_06630_),
    .Y(_06631_));
 sky130_fd_sc_hd__nand3b_2 _28651_ (.A_N(_06625_),
    .B(_06273_),
    .C(_06622_),
    .Y(_06632_));
 sky130_fd_sc_hd__nand2_2 _28652_ (.A(_06625_),
    .B(_06626_),
    .Y(_06633_));
 sky130_fd_sc_hd__nand3_2 _28653_ (.A(_06632_),
    .B(_06633_),
    .C(_06630_),
    .Y(_06634_));
 sky130_fd_sc_hd__a21oi_2 _28654_ (.A1(_06449_),
    .A2(_06450_),
    .B1(_06445_),
    .Y(_06635_));
 sky130_fd_sc_hd__a21o_2 _28655_ (.A1(_06631_),
    .A2(_06634_),
    .B1(_06635_),
    .X(_06636_));
 sky130_fd_sc_hd__nand3_2 _28656_ (.A(_06631_),
    .B(_06634_),
    .C(_06635_),
    .Y(_06637_));
 sky130_fd_sc_hd__nand2_2 _28657_ (.A(_06636_),
    .B(_06637_),
    .Y(_06638_));
 sky130_fd_sc_hd__xor2_2 _28658_ (.A(_06621_),
    .B(_06638_),
    .X(_06639_));
 sky130_fd_sc_hd__nor2_2 _28659_ (.A(_06604_),
    .B(_06639_),
    .Y(_06640_));
 sky130_fd_sc_hd__nand2_2 _28660_ (.A(_06639_),
    .B(_06604_),
    .Y(_06641_));
 sky130_fd_sc_hd__nand2_2 _28661_ (.A(_06463_),
    .B(_06641_),
    .Y(_06642_));
 sky130_fd_sc_hd__nor2_2 _28662_ (.A(_06640_),
    .B(_06642_),
    .Y(_06643_));
 sky130_fd_sc_hd__inv_2 _28663_ (.A(_06640_),
    .Y(_06644_));
 sky130_fd_sc_hd__a21oi_2 _28664_ (.A1(_06644_),
    .A2(_06641_),
    .B1(_06463_),
    .Y(_06645_));
 sky130_fd_sc_hd__nor2_2 _28665_ (.A(_06643_),
    .B(_06645_),
    .Y(_06646_));
 sky130_fd_sc_hd__a21oi_2 _28666_ (.A1(_06587_),
    .A2(_06597_),
    .B1(_06646_),
    .Y(_06647_));
 sky130_fd_sc_hd__a21boi_2 _28667_ (.A1(_06644_),
    .A2(_06641_),
    .B1_N(_06463_),
    .Y(_06648_));
 sky130_fd_sc_hd__o211a_2 _28668_ (.A1(_06429_),
    .A2(_06462_),
    .B1(_06641_),
    .C1(_06644_),
    .X(_06649_));
 sky130_fd_sc_hd__o211a_2 _28669_ (.A1(_06648_),
    .A2(_06649_),
    .B1(_06597_),
    .C1(_06587_),
    .X(_06650_));
 sky130_fd_sc_hd__o22ai_2 _28670_ (.A1(_06466_),
    .A2(_06428_),
    .B1(_06647_),
    .B2(_06650_),
    .Y(_06651_));
 sky130_fd_sc_hd__a21o_2 _28671_ (.A1(_06587_),
    .A2(_06597_),
    .B1(_06646_),
    .X(_06652_));
 sky130_fd_sc_hd__nand3_2 _28672_ (.A(_06587_),
    .B(_06596_),
    .C(_06646_),
    .Y(_06653_));
 sky130_fd_sc_hd__nand3_2 _28673_ (.A(_06652_),
    .B(_06471_),
    .C(_06653_),
    .Y(_06654_));
 sky130_fd_sc_hd__nand2_2 _28674_ (.A(_06651_),
    .B(_06654_),
    .Y(_06655_));
 sky130_fd_sc_hd__and3_2 _28675_ (.A(_06367_),
    .B(_06405_),
    .C(_06406_),
    .X(_06656_));
 sky130_fd_sc_hd__o21a_2 _28676_ (.A1(_06656_),
    .A2(_06417_),
    .B1(_06427_),
    .X(_06657_));
 sky130_fd_sc_hd__nor2_2 _28677_ (.A(_06656_),
    .B(_06410_),
    .Y(_06658_));
 sky130_fd_sc_hd__and2b_2 _28678_ (.A_N(_06426_),
    .B(_06658_),
    .X(_06659_));
 sky130_fd_sc_hd__nor2_2 _28679_ (.A(_06657_),
    .B(_06659_),
    .Y(_06660_));
 sky130_fd_sc_hd__nand2_2 _28680_ (.A(_06655_),
    .B(_06660_),
    .Y(_06661_));
 sky130_fd_sc_hd__o21ai_2 _28681_ (.A1(_06476_),
    .A2(_06469_),
    .B1(_06475_),
    .Y(_06662_));
 sky130_fd_sc_hd__nand3b_2 _28682_ (.A_N(_06660_),
    .B(_06654_),
    .C(_06651_),
    .Y(_06663_));
 sky130_fd_sc_hd__nand3_2 _28683_ (.A(_06661_),
    .B(_06662_),
    .C(_06663_),
    .Y(_06664_));
 sky130_fd_sc_hd__o2bb2ai_2 _28684_ (.A1_N(_06654_),
    .A2_N(_06651_),
    .B1(_06657_),
    .B2(_06659_),
    .Y(_06665_));
 sky130_fd_sc_hd__nor2_2 _28685_ (.A(_06319_),
    .B(_06292_),
    .Y(_06666_));
 sky130_fd_sc_hd__and2_2 _28686_ (.A(_06292_),
    .B(_06319_),
    .X(_06667_));
 sky130_fd_sc_hd__nor2_2 _28687_ (.A(_06666_),
    .B(_06667_),
    .Y(_06668_));
 sky130_fd_sc_hd__a21oi_2 _28688_ (.A1(_06474_),
    .A2(_06668_),
    .B1(_06472_),
    .Y(_06669_));
 sky130_fd_sc_hd__nand3_2 _28689_ (.A(_06651_),
    .B(_06654_),
    .C(_06660_),
    .Y(_06670_));
 sky130_fd_sc_hd__nand3_2 _28690_ (.A(_06665_),
    .B(_06669_),
    .C(_06670_),
    .Y(_06671_));
 sky130_fd_sc_hd__a21oi_2 _28691_ (.A1(_06664_),
    .A2(_06671_),
    .B1(_06666_),
    .Y(_06672_));
 sky130_fd_sc_hd__and3_2 _28692_ (.A(_06664_),
    .B(_06671_),
    .C(_06666_),
    .X(_06673_));
 sky130_fd_sc_hd__nand2_2 _28693_ (.A(_06484_),
    .B(_06480_),
    .Y(_06674_));
 sky130_fd_sc_hd__o21bai_2 _28694_ (.A1(_06672_),
    .A2(_06673_),
    .B1_N(_06674_),
    .Y(_06675_));
 sky130_fd_sc_hd__nand3_2 _28695_ (.A(_06664_),
    .B(_06671_),
    .C(_06666_),
    .Y(_06676_));
 sky130_fd_sc_hd__nand3b_2 _28696_ (.A_N(_06672_),
    .B(_06676_),
    .C(_06674_),
    .Y(_06677_));
 sky130_fd_sc_hd__nand2_2 _28697_ (.A(_06675_),
    .B(_06677_),
    .Y(_06678_));
 sky130_fd_sc_hd__or2_2 _28698_ (.A(_06678_),
    .B(_06491_),
    .X(_06679_));
 sky130_fd_sc_hd__nand2_2 _28699_ (.A(_06491_),
    .B(_06678_),
    .Y(_06680_));
 sky130_fd_sc_hd__and2_2 _28700_ (.A(_06679_),
    .B(_06680_),
    .X(_02635_));
 sky130_fd_sc_hd__and2b_2 _28701_ (.A_N(_06575_),
    .B(_06578_),
    .X(_06681_));
 sky130_fd_sc_hd__nor2_2 _28702_ (.A(_06681_),
    .B(_06597_),
    .Y(_06682_));
 sky130_fd_sc_hd__and2_2 _28703_ (.A(_06597_),
    .B(_06681_),
    .X(_06683_));
 sky130_fd_sc_hd__nand2_2 _28704_ (.A(_06526_),
    .B(_06525_),
    .Y(_06684_));
 sky130_fd_sc_hd__nand2_2 _28705_ (.A(_06531_),
    .B(_06528_),
    .Y(_06685_));
 sky130_fd_sc_hd__inv_2 _28706_ (.A(_06516_),
    .Y(_06686_));
 sky130_fd_sc_hd__o21a_2 _28707_ (.A1(_06517_),
    .A2(_06518_),
    .B1(_06511_),
    .X(_06687_));
 sky130_fd_sc_hd__buf_1 _28708_ (.A(_06224_),
    .X(_06688_));
 sky130_fd_sc_hd__a22oi_2 _28709_ (.A1(_05639_),
    .A2(_19613_),
    .B1(_05760_),
    .B2(_05598_),
    .Y(_06689_));
 sky130_fd_sc_hd__nand2_2 _28710_ (.A(_06008_),
    .B(_05614_),
    .Y(_06690_));
 sky130_fd_sc_hd__nand2_2 _28711_ (.A(_06010_),
    .B(_06497_),
    .Y(_06691_));
 sky130_fd_sc_hd__nor2_2 _28712_ (.A(_06690_),
    .B(_06691_),
    .Y(_06692_));
 sky130_fd_sc_hd__o22ai_2 _28713_ (.A1(_05244_),
    .A2(_06688_),
    .B1(_06689_),
    .B2(_06692_),
    .Y(_06693_));
 sky130_fd_sc_hd__inv_2 _28714_ (.A(_05597_),
    .Y(_06694_));
 sky130_fd_sc_hd__nand3_2 _28715_ (.A(_05851_),
    .B(_06508_),
    .C(_05734_),
    .Y(_06695_));
 sky130_fd_sc_hd__nand2_2 _28716_ (.A(_06690_),
    .B(_06691_),
    .Y(_06696_));
 sky130_fd_sc_hd__nand2_2 _28717_ (.A(_06496_),
    .B(_06539_),
    .Y(_06697_));
 sky130_fd_sc_hd__inv_2 _28718_ (.A(_06697_),
    .Y(_06698_));
 sky130_fd_sc_hd__o211ai_2 _28719_ (.A1(_06694_),
    .A2(_06695_),
    .B1(_06696_),
    .C1(_06698_),
    .Y(_06699_));
 sky130_fd_sc_hd__o22ai_2 _28720_ (.A1(_05856_),
    .A2(_06615_),
    .B1(_06618_),
    .B2(_06607_),
    .Y(_06700_));
 sky130_fd_sc_hd__nand3_2 _28721_ (.A(_06693_),
    .B(_06699_),
    .C(_06700_),
    .Y(_06701_));
 sky130_fd_sc_hd__buf_1 _28722_ (.A(_06701_),
    .X(_06702_));
 sky130_fd_sc_hd__o21ai_2 _28723_ (.A1(_06689_),
    .A2(_06692_),
    .B1(_06698_),
    .Y(_06703_));
 sky130_fd_sc_hd__a21oi_2 _28724_ (.A1(_06619_),
    .A2(_06612_),
    .B1(_06611_),
    .Y(_06704_));
 sky130_fd_sc_hd__o211ai_2 _28725_ (.A1(_06694_),
    .A2(_06695_),
    .B1(_06697_),
    .C1(_06696_),
    .Y(_06705_));
 sky130_fd_sc_hd__nand3_2 _28726_ (.A(_06703_),
    .B(_06704_),
    .C(_06705_),
    .Y(_06706_));
 sky130_fd_sc_hd__nor2_2 _28727_ (.A(_06506_),
    .B(_06495_),
    .Y(_06707_));
 sky130_fd_sc_hd__o2bb2ai_2 _28728_ (.A1_N(_06702_),
    .A2_N(_06706_),
    .B1(_06493_),
    .B2(_06707_),
    .Y(_06708_));
 sky130_fd_sc_hd__a21oi_2 _28729_ (.A1(_06509_),
    .A2(_06506_),
    .B1(_06495_),
    .Y(_06709_));
 sky130_fd_sc_hd__nand3b_2 _28730_ (.A_N(_06709_),
    .B(_06706_),
    .C(_06701_),
    .Y(_06710_));
 sky130_fd_sc_hd__nand2_2 _28731_ (.A(_06637_),
    .B(_06621_),
    .Y(_06711_));
 sky130_fd_sc_hd__nand2_2 _28732_ (.A(_06711_),
    .B(_06636_),
    .Y(_06712_));
 sky130_fd_sc_hd__a21oi_2 _28733_ (.A1(_06708_),
    .A2(_06710_),
    .B1(_06712_),
    .Y(_06713_));
 sky130_fd_sc_hd__a31oi_2 _28734_ (.A1(_06703_),
    .A2(_06704_),
    .A3(_06705_),
    .B1(_06709_),
    .Y(_06714_));
 sky130_fd_sc_hd__a2bb2oi_2 _28735_ (.A1_N(_06493_),
    .A2_N(_06707_),
    .B1(_06702_),
    .B2(_06706_),
    .Y(_06715_));
 sky130_fd_sc_hd__a221oi_2 _28736_ (.A1(_06714_),
    .A2(_06702_),
    .B1(_06711_),
    .B2(_06636_),
    .C1(_06715_),
    .Y(_06716_));
 sky130_fd_sc_hd__o22ai_2 _28737_ (.A1(_06686_),
    .A2(_06687_),
    .B1(_06713_),
    .B2(_06716_),
    .Y(_06717_));
 sky130_fd_sc_hd__a21o_2 _28738_ (.A1(_06708_),
    .A2(_06710_),
    .B1(_06712_),
    .X(_06718_));
 sky130_fd_sc_hd__nand3_2 _28739_ (.A(_06712_),
    .B(_06710_),
    .C(_06708_),
    .Y(_06719_));
 sky130_fd_sc_hd__nand2_2 _28740_ (.A(_06520_),
    .B(_06511_),
    .Y(_06720_));
 sky130_fd_sc_hd__nand3_2 _28741_ (.A(_06718_),
    .B(_06719_),
    .C(_06720_),
    .Y(_06721_));
 sky130_fd_sc_hd__a22oi_2 _28742_ (.A1(_06684_),
    .A2(_06685_),
    .B1(_06717_),
    .B2(_06721_),
    .Y(_06722_));
 sky130_fd_sc_hd__o211a_2 _28743_ (.A1(_06527_),
    .A2(_06530_),
    .B1(_06721_),
    .C1(_06717_),
    .X(_06723_));
 sky130_fd_sc_hd__buf_1 _28744_ (.A(_19599_),
    .X(_06724_));
 sky130_fd_sc_hd__a22oi_2 _28745_ (.A1(_19388_),
    .A2(_05897_),
    .B1(_06201_),
    .B2(_06724_),
    .Y(_06725_));
 sky130_fd_sc_hd__buf_1 _28746_ (.A(_19602_),
    .X(_06726_));
 sky130_fd_sc_hd__and4_2 _28747_ (.A(_06051_),
    .B(_06054_),
    .C(_06724_),
    .D(_06726_),
    .X(_06727_));
 sky130_fd_sc_hd__buf_1 _28748_ (.A(_19587_),
    .X(_06728_));
 sky130_fd_sc_hd__nand2_2 _28749_ (.A(_06057_),
    .B(_06728_),
    .Y(_06729_));
 sky130_fd_sc_hd__o21ai_2 _28750_ (.A1(_06725_),
    .A2(_06727_),
    .B1(_06729_),
    .Y(_06730_));
 sky130_fd_sc_hd__buf_1 _28751_ (.A(_19387_),
    .X(_06731_));
 sky130_fd_sc_hd__buf_1 _28752_ (.A(\pcpi_mul.rs1[12] ),
    .X(_06732_));
 sky130_fd_sc_hd__nand2_2 _28753_ (.A(_06731_),
    .B(_06732_),
    .Y(_06733_));
 sky130_fd_sc_hd__nand3b_2 _28754_ (.A_N(_06733_),
    .B(_06054_),
    .C(_06059_),
    .Y(_06734_));
 sky130_fd_sc_hd__buf_1 _28755_ (.A(_05187_),
    .X(_06735_));
 sky130_fd_sc_hd__buf_1 _28756_ (.A(_06058_),
    .X(_06736_));
 sky130_fd_sc_hd__a22o_2 _28757_ (.A1(_06735_),
    .A2(_19603_),
    .B1(_05403_),
    .B2(_06736_),
    .X(_06737_));
 sky130_fd_sc_hd__inv_2 _28758_ (.A(_06729_),
    .Y(_06738_));
 sky130_fd_sc_hd__nand3_2 _28759_ (.A(_06734_),
    .B(_06737_),
    .C(_06738_),
    .Y(_06739_));
 sky130_fd_sc_hd__o21ai_2 _28760_ (.A1(_06543_),
    .A2(_06537_),
    .B1(_06547_),
    .Y(_06740_));
 sky130_fd_sc_hd__nand3_2 _28761_ (.A(_06730_),
    .B(_06739_),
    .C(_06740_),
    .Y(_06741_));
 sky130_fd_sc_hd__o21ai_2 _28762_ (.A1(_06725_),
    .A2(_06727_),
    .B1(_06738_),
    .Y(_06742_));
 sky130_fd_sc_hd__a21oi_2 _28763_ (.A1(_06548_),
    .A2(_06544_),
    .B1(_06541_),
    .Y(_06743_));
 sky130_fd_sc_hd__nand3_2 _28764_ (.A(_06734_),
    .B(_06737_),
    .C(_06729_),
    .Y(_06744_));
 sky130_fd_sc_hd__nand3_2 _28765_ (.A(_06742_),
    .B(_06743_),
    .C(_06744_),
    .Y(_06745_));
 sky130_fd_sc_hd__nand2_2 _28766_ (.A(_05205_),
    .B(_19590_),
    .Y(_06746_));
 sky130_fd_sc_hd__nand3_2 _28767_ (.A(_06746_),
    .B(_05123_),
    .C(_06557_),
    .Y(_06747_));
 sky130_fd_sc_hd__buf_1 _28768_ (.A(_06372_),
    .X(_06748_));
 sky130_fd_sc_hd__nand2_2 _28769_ (.A(_19398_),
    .B(_06748_),
    .Y(_06749_));
 sky130_fd_sc_hd__buf_1 _28770_ (.A(_06542_),
    .X(_06750_));
 sky130_fd_sc_hd__nand3_2 _28771_ (.A(_06749_),
    .B(_05118_),
    .C(_06750_),
    .Y(_06751_));
 sky130_fd_sc_hd__nand2_2 _28772_ (.A(_05115_),
    .B(_06388_),
    .Y(_06752_));
 sky130_fd_sc_hd__and3_2 _28773_ (.A(_06747_),
    .B(_06751_),
    .C(_06752_),
    .X(_06753_));
 sky130_fd_sc_hd__a21oi_2 _28774_ (.A1(_06747_),
    .A2(_06751_),
    .B1(_06752_),
    .Y(_06754_));
 sky130_fd_sc_hd__o2bb2ai_2 _28775_ (.A1_N(_06741_),
    .A2_N(_06745_),
    .B1(_06753_),
    .B2(_06754_),
    .Y(_06755_));
 sky130_fd_sc_hd__nor2_2 _28776_ (.A(_06754_),
    .B(_06753_),
    .Y(_06756_));
 sky130_fd_sc_hd__nand3_2 _28777_ (.A(_06756_),
    .B(_06745_),
    .C(_06741_),
    .Y(_06757_));
 sky130_fd_sc_hd__nand2_2 _28778_ (.A(_06755_),
    .B(_06757_),
    .Y(_06758_));
 sky130_fd_sc_hd__a21oi_2 _28779_ (.A1(_06552_),
    .A2(_06553_),
    .B1(_06554_),
    .Y(_06759_));
 sky130_fd_sc_hd__o21a_2 _28780_ (.A1(_06759_),
    .A2(_06566_),
    .B1(_06551_),
    .X(_06760_));
 sky130_fd_sc_hd__nand2_2 _28781_ (.A(_06758_),
    .B(_06760_),
    .Y(_06761_));
 sky130_fd_sc_hd__o21ai_2 _28782_ (.A1(_06759_),
    .A2(_06566_),
    .B1(_06551_),
    .Y(_06762_));
 sky130_fd_sc_hd__nand3_2 _28783_ (.A(_06762_),
    .B(_06755_),
    .C(_06757_),
    .Y(_06763_));
 sky130_fd_sc_hd__nor2_2 _28784_ (.A(_06558_),
    .B(_06561_),
    .Y(_06764_));
 sky130_fd_sc_hd__inv_2 _28785_ (.A(_06564_),
    .Y(_06765_));
 sky130_fd_sc_hd__nor2_2 _28786_ (.A(_06764_),
    .B(_06765_),
    .Y(_06766_));
 sky130_fd_sc_hd__inv_2 _28787_ (.A(_06766_),
    .Y(_06767_));
 sky130_fd_sc_hd__a21oi_2 _28788_ (.A1(_06761_),
    .A2(_06763_),
    .B1(_06767_),
    .Y(_06768_));
 sky130_fd_sc_hd__o211a_2 _28789_ (.A1(_06764_),
    .A2(_06765_),
    .B1(_06763_),
    .C1(_06761_),
    .X(_06769_));
 sky130_fd_sc_hd__nor2_2 _28790_ (.A(_06768_),
    .B(_06769_),
    .Y(_06770_));
 sky130_fd_sc_hd__o21ai_2 _28791_ (.A1(_06722_),
    .A2(_06723_),
    .B1(_06770_),
    .Y(_06771_));
 sky130_fd_sc_hd__nand3_2 _28792_ (.A(_06644_),
    .B(_06463_),
    .C(_06641_),
    .Y(_06772_));
 sky130_fd_sc_hd__o21ai_2 _28793_ (.A1(_06528_),
    .A2(_06524_),
    .B1(_06531_),
    .Y(_06773_));
 sky130_fd_sc_hd__a21o_2 _28794_ (.A1(_06717_),
    .A2(_06721_),
    .B1(_06773_),
    .X(_06774_));
 sky130_fd_sc_hd__nand3_2 _28795_ (.A(_06773_),
    .B(_06717_),
    .C(_06721_),
    .Y(_06775_));
 sky130_fd_sc_hd__a21o_2 _28796_ (.A1(_06761_),
    .A2(_06763_),
    .B1(_06767_),
    .X(_06776_));
 sky130_fd_sc_hd__nand3_2 _28797_ (.A(_06761_),
    .B(_06763_),
    .C(_06767_),
    .Y(_06777_));
 sky130_fd_sc_hd__nand2_2 _28798_ (.A(_06776_),
    .B(_06777_),
    .Y(_06778_));
 sky130_fd_sc_hd__nand3_2 _28799_ (.A(_06774_),
    .B(_06775_),
    .C(_06778_),
    .Y(_06779_));
 sky130_fd_sc_hd__nand3_2 _28800_ (.A(_06771_),
    .B(_06772_),
    .C(_06779_),
    .Y(_06780_));
 sky130_fd_sc_hd__o22ai_2 _28801_ (.A1(_06769_),
    .A2(_06768_),
    .B1(_06722_),
    .B2(_06723_),
    .Y(_06781_));
 sky130_fd_sc_hd__nand3_2 _28802_ (.A(_06774_),
    .B(_06770_),
    .C(_06775_),
    .Y(_06782_));
 sky130_fd_sc_hd__nand3_2 _28803_ (.A(_06781_),
    .B(_06643_),
    .C(_06782_),
    .Y(_06783_));
 sky130_fd_sc_hd__buf_1 _28804_ (.A(_06783_),
    .X(_06784_));
 sky130_fd_sc_hd__nor2_2 _28805_ (.A(_06580_),
    .B(_06536_),
    .Y(_06785_));
 sky130_fd_sc_hd__o2bb2ai_2 _28806_ (.A1_N(_06780_),
    .A2_N(_06784_),
    .B1(_06534_),
    .B2(_06785_),
    .Y(_06786_));
 sky130_fd_sc_hd__o21ai_2 _28807_ (.A1(_06534_),
    .A2(_06583_),
    .B1(_06585_),
    .Y(_06787_));
 sky130_fd_sc_hd__nand3_2 _28808_ (.A(_06780_),
    .B(_06783_),
    .C(_06787_),
    .Y(_06788_));
 sky130_fd_sc_hd__buf_1 _28809_ (.A(_06788_),
    .X(_06789_));
 sky130_fd_sc_hd__buf_1 _28810_ (.A(_06270_),
    .X(_06790_));
 sky130_fd_sc_hd__a22oi_2 _28811_ (.A1(_06790_),
    .A2(_06622_),
    .B1(_06115_),
    .B2(_19628_),
    .Y(_06791_));
 sky130_fd_sc_hd__buf_1 _28812_ (.A(_05146_),
    .X(_06792_));
 sky130_fd_sc_hd__nand2_2 _28813_ (.A(_06624_),
    .B(_06792_),
    .Y(_06793_));
 sky130_fd_sc_hd__nand2_2 _28814_ (.A(_06272_),
    .B(_19627_),
    .Y(_06794_));
 sky130_fd_sc_hd__nor2_2 _28815_ (.A(_06793_),
    .B(_06794_),
    .Y(_06795_));
 sky130_fd_sc_hd__nand2_2 _28816_ (.A(_06446_),
    .B(_19625_),
    .Y(_06796_));
 sky130_fd_sc_hd__inv_2 _28817_ (.A(_06796_),
    .Y(_06797_));
 sky130_fd_sc_hd__o21ai_2 _28818_ (.A1(_06791_),
    .A2(_06795_),
    .B1(_06797_),
    .Y(_06798_));
 sky130_fd_sc_hd__nand3b_2 _28819_ (.A_N(_06793_),
    .B(_19366_),
    .C(_19628_),
    .Y(_06799_));
 sky130_fd_sc_hd__nand2_2 _28820_ (.A(_06793_),
    .B(_06794_),
    .Y(_06800_));
 sky130_fd_sc_hd__nand3_2 _28821_ (.A(_06799_),
    .B(_06796_),
    .C(_06800_),
    .Y(_06801_));
 sky130_fd_sc_hd__o21ai_2 _28822_ (.A1(_06625_),
    .A2(_06626_),
    .B1(_06630_),
    .Y(_06802_));
 sky130_fd_sc_hd__nand2_2 _28823_ (.A(_06802_),
    .B(_06633_),
    .Y(_06803_));
 sky130_fd_sc_hd__a21o_2 _28824_ (.A1(_06798_),
    .A2(_06801_),
    .B1(_06803_),
    .X(_06804_));
 sky130_fd_sc_hd__nand3_2 _28825_ (.A(_06798_),
    .B(_06801_),
    .C(_06803_),
    .Y(_06805_));
 sky130_fd_sc_hd__nand2_2 _28826_ (.A(_06804_),
    .B(_06805_),
    .Y(_06806_));
 sky130_fd_sc_hd__nand2_2 _28827_ (.A(_19370_),
    .B(_05958_),
    .Y(_06807_));
 sky130_fd_sc_hd__buf_1 _28828_ (.A(_05419_),
    .X(_06808_));
 sky130_fd_sc_hd__nand2_2 _28829_ (.A(_06808_),
    .B(_06609_),
    .Y(_06809_));
 sky130_fd_sc_hd__nor2_2 _28830_ (.A(_06807_),
    .B(_06809_),
    .Y(_06810_));
 sky130_fd_sc_hd__nand2_2 _28831_ (.A(_05672_),
    .B(_05408_),
    .Y(_06811_));
 sky130_fd_sc_hd__a22o_2 _28832_ (.A1(_06256_),
    .A2(_05422_),
    .B1(_06258_),
    .B2(_19619_),
    .X(_06812_));
 sky130_fd_sc_hd__nand3b_2 _28833_ (.A_N(_06810_),
    .B(_06811_),
    .C(_06812_),
    .Y(_06813_));
 sky130_fd_sc_hd__a22oi_2 _28834_ (.A1(_05801_),
    .A2(_05425_),
    .B1(_05803_),
    .B2(_06617_),
    .Y(_06814_));
 sky130_fd_sc_hd__inv_2 _28835_ (.A(_06811_),
    .Y(_06815_));
 sky130_fd_sc_hd__o21ai_2 _28836_ (.A1(_06814_),
    .A2(_06810_),
    .B1(_06815_),
    .Y(_06816_));
 sky130_fd_sc_hd__nand2_2 _28837_ (.A(_06813_),
    .B(_06816_),
    .Y(_06817_));
 sky130_fd_sc_hd__nand2_2 _28838_ (.A(_06806_),
    .B(_06817_),
    .Y(_06818_));
 sky130_fd_sc_hd__nand3b_2 _28839_ (.A_N(_06817_),
    .B(_06804_),
    .C(_06805_),
    .Y(_06819_));
 sky130_fd_sc_hd__nand2_2 _28840_ (.A(_06818_),
    .B(_06819_),
    .Y(_06820_));
 sky130_fd_sc_hd__buf_1 _28841_ (.A(\pcpi_mul.rs2[17] ),
    .X(_06821_));
 sky130_fd_sc_hd__buf_1 _28842_ (.A(_06821_),
    .X(_06822_));
 sky130_fd_sc_hd__buf_1 _28843_ (.A(\pcpi_mul.rs2[16] ),
    .X(_06823_));
 sky130_fd_sc_hd__buf_1 _28844_ (.A(_06823_),
    .X(_06824_));
 sky130_fd_sc_hd__and4_2 _28845_ (.A(_06822_),
    .B(_06824_),
    .C(_19636_),
    .D(_19640_),
    .X(_06825_));
 sky130_fd_sc_hd__inv_2 _28846_ (.A(_19354_),
    .Y(_06826_));
 sky130_fd_sc_hd__buf_1 _28847_ (.A(_19356_),
    .X(_06827_));
 sky130_fd_sc_hd__buf_1 _28848_ (.A(_06827_),
    .X(_06828_));
 sky130_fd_sc_hd__nand2_2 _28849_ (.A(_06828_),
    .B(_05804_),
    .Y(_06829_));
 sky130_fd_sc_hd__o21ai_2 _28850_ (.A1(_06826_),
    .A2(_04838_),
    .B1(_06829_),
    .Y(_06830_));
 sky130_fd_sc_hd__inv_2 _28851_ (.A(\pcpi_mul.rs2[15] ),
    .Y(_06831_));
 sky130_fd_sc_hd__nor2_2 _28852_ (.A(_06831_),
    .B(_05256_),
    .Y(_06832_));
 sky130_fd_sc_hd__nand2_2 _28853_ (.A(_06830_),
    .B(_06832_),
    .Y(_06833_));
 sky130_fd_sc_hd__o21a_2 _28854_ (.A1(_06826_),
    .A2(_04838_),
    .B1(_06829_),
    .X(_06834_));
 sky130_fd_sc_hd__o21bai_2 _28855_ (.A1(_06825_),
    .A2(_06834_),
    .B1_N(_06832_),
    .Y(_06835_));
 sky130_fd_sc_hd__o21ai_2 _28856_ (.A1(_06825_),
    .A2(_06833_),
    .B1(_06835_),
    .Y(_06836_));
 sky130_fd_sc_hd__nand2_2 _28857_ (.A(_06836_),
    .B(_06601_),
    .Y(_06837_));
 sky130_fd_sc_hd__or2_2 _28858_ (.A(_06601_),
    .B(_06836_),
    .X(_06838_));
 sky130_fd_sc_hd__nand3b_2 _28859_ (.A_N(_06820_),
    .B(_06837_),
    .C(_06838_),
    .Y(_06839_));
 sky130_fd_sc_hd__a22o_2 _28860_ (.A1(_06818_),
    .A2(_06819_),
    .B1(_06837_),
    .B2(_06838_),
    .X(_06840_));
 sky130_fd_sc_hd__nand2_2 _28861_ (.A(_06839_),
    .B(_06840_),
    .Y(_06841_));
 sky130_fd_sc_hd__or2b_2 _28862_ (.A(_06841_),
    .B_N(_06640_),
    .X(_06842_));
 sky130_fd_sc_hd__nand2_2 _28863_ (.A(_06644_),
    .B(_06841_),
    .Y(_06843_));
 sky130_fd_sc_hd__nand2_2 _28864_ (.A(_06842_),
    .B(_06843_),
    .Y(_06844_));
 sky130_fd_sc_hd__inv_2 _28865_ (.A(_06844_),
    .Y(_06845_));
 sky130_fd_sc_hd__a21oi_2 _28866_ (.A1(_06786_),
    .A2(_06789_),
    .B1(_06845_),
    .Y(_06846_));
 sky130_fd_sc_hd__a21oi_2 _28867_ (.A1(_06780_),
    .A2(_06783_),
    .B1(_06787_),
    .Y(_06847_));
 sky130_fd_sc_hd__nand2_2 _28868_ (.A(_06788_),
    .B(_06845_),
    .Y(_06848_));
 sky130_fd_sc_hd__o21bai_2 _28869_ (.A1(_06847_),
    .A2(_06848_),
    .B1_N(_06653_),
    .Y(_06849_));
 sky130_fd_sc_hd__nor2_2 _28870_ (.A(_06846_),
    .B(_06849_),
    .Y(_06850_));
 sky130_fd_sc_hd__nor2_2 _28871_ (.A(_06841_),
    .B(_06644_),
    .Y(_06851_));
 sky130_fd_sc_hd__inv_2 _28872_ (.A(_06843_),
    .Y(_06852_));
 sky130_fd_sc_hd__and3_2 _28873_ (.A(_06780_),
    .B(_06784_),
    .C(_06787_),
    .X(_06853_));
 sky130_fd_sc_hd__o22ai_2 _28874_ (.A1(_06851_),
    .A2(_06852_),
    .B1(_06847_),
    .B2(_06853_),
    .Y(_06854_));
 sky130_fd_sc_hd__nand3_2 _28875_ (.A(_06786_),
    .B(_06845_),
    .C(_06789_),
    .Y(_06855_));
 sky130_fd_sc_hd__a21oi_2 _28876_ (.A1(_06854_),
    .A2(_06855_),
    .B1(_06650_),
    .Y(_06856_));
 sky130_fd_sc_hd__o22ai_2 _28877_ (.A1(_06682_),
    .A2(_06683_),
    .B1(_06850_),
    .B2(_06856_),
    .Y(_06857_));
 sky130_fd_sc_hd__nor2_2 _28878_ (.A(_06847_),
    .B(_06848_),
    .Y(_06858_));
 sky130_fd_sc_hd__o21ai_2 _28879_ (.A1(_06858_),
    .A2(_06846_),
    .B1(_06653_),
    .Y(_06859_));
 sky130_fd_sc_hd__nor2_2 _28880_ (.A(_06682_),
    .B(_06683_),
    .Y(_06860_));
 sky130_fd_sc_hd__nand3_2 _28881_ (.A(_06854_),
    .B(_06650_),
    .C(_06855_),
    .Y(_06861_));
 sky130_fd_sc_hd__nand3_2 _28882_ (.A(_06859_),
    .B(_06860_),
    .C(_06861_),
    .Y(_06862_));
 sky130_fd_sc_hd__a21oi_2 _28883_ (.A1(_06652_),
    .A2(_06653_),
    .B1(_06471_),
    .Y(_06863_));
 sky130_fd_sc_hd__o21ai_2 _28884_ (.A1(_06660_),
    .A2(_06863_),
    .B1(_06654_),
    .Y(_06864_));
 sky130_fd_sc_hd__nand3_2 _28885_ (.A(_06857_),
    .B(_06862_),
    .C(_06864_),
    .Y(_06865_));
 sky130_fd_sc_hd__o21ai_2 _28886_ (.A1(_06850_),
    .A2(_06856_),
    .B1(_06860_),
    .Y(_06866_));
 sky130_fd_sc_hd__o21a_2 _28887_ (.A1(_06660_),
    .A2(_06863_),
    .B1(_06654_),
    .X(_06867_));
 sky130_fd_sc_hd__inv_2 _28888_ (.A(_06860_),
    .Y(_06868_));
 sky130_fd_sc_hd__nand3_2 _28889_ (.A(_06859_),
    .B(_06868_),
    .C(_06861_),
    .Y(_06869_));
 sky130_fd_sc_hd__nand3_2 _28890_ (.A(_06866_),
    .B(_06867_),
    .C(_06869_),
    .Y(_06870_));
 sky130_fd_sc_hd__o2bb2ai_2 _28891_ (.A1_N(_06865_),
    .A2_N(_06870_),
    .B1(_06427_),
    .B2(_06658_),
    .Y(_06871_));
 sky130_fd_sc_hd__nor2_2 _28892_ (.A(_06658_),
    .B(_06427_),
    .Y(_06872_));
 sky130_fd_sc_hd__nand2_2 _28893_ (.A(_06870_),
    .B(_06872_),
    .Y(_06873_));
 sky130_fd_sc_hd__nand2_2 _28894_ (.A(_06676_),
    .B(_06664_),
    .Y(_06874_));
 sky130_fd_sc_hd__a21oi_2 _28895_ (.A1(_06871_),
    .A2(_06873_),
    .B1(_06874_),
    .Y(_06875_));
 sky130_fd_sc_hd__nand3_2 _28896_ (.A(_06871_),
    .B(_06874_),
    .C(_06873_),
    .Y(_06876_));
 sky130_fd_sc_hd__and2b_2 _28897_ (.A_N(_06875_),
    .B(_06876_),
    .X(_06877_));
 sky130_fd_sc_hd__nand2_2 _28898_ (.A(_06679_),
    .B(_06677_),
    .Y(_06878_));
 sky130_fd_sc_hd__xor2_2 _28899_ (.A(_06877_),
    .B(_06878_),
    .X(_02636_));
 sky130_fd_sc_hd__inv_2 _28900_ (.A(_06761_),
    .Y(_06879_));
 sky130_fd_sc_hd__o21a_2 _28901_ (.A1(_06766_),
    .A2(_06879_),
    .B1(_06763_),
    .X(_06880_));
 sky130_fd_sc_hd__inv_2 _28902_ (.A(_06880_),
    .Y(_06881_));
 sky130_fd_sc_hd__and2_2 _28903_ (.A(_06789_),
    .B(_06784_),
    .X(_06882_));
 sky130_fd_sc_hd__nor2_2 _28904_ (.A(_06881_),
    .B(_06882_),
    .Y(_06883_));
 sky130_fd_sc_hd__and3_2 _28905_ (.A(_06789_),
    .B(_06784_),
    .C(_06881_),
    .X(_06884_));
 sky130_fd_sc_hd__and2_2 _28906_ (.A(_06520_),
    .B(_06511_),
    .X(_06885_));
 sky130_fd_sc_hd__nand2_2 _28907_ (.A(_06719_),
    .B(_06885_),
    .Y(_06886_));
 sky130_fd_sc_hd__inv_2 _28908_ (.A(_06706_),
    .Y(_06887_));
 sky130_fd_sc_hd__and2_2 _28909_ (.A(_06702_),
    .B(_06709_),
    .X(_06888_));
 sky130_fd_sc_hd__buf_1 _28910_ (.A(_05597_),
    .X(_06889_));
 sky130_fd_sc_hd__a22oi_2 _28911_ (.A1(_05851_),
    .A2(_06889_),
    .B1(_06508_),
    .B2(_05717_),
    .Y(_06890_));
 sky130_fd_sc_hd__nand3_2 _28912_ (.A(_19379_),
    .B(_06334_),
    .C(_19608_),
    .Y(_06891_));
 sky130_fd_sc_hd__nor2_2 _28913_ (.A(_06224_),
    .B(_06891_),
    .Y(_06892_));
 sky130_fd_sc_hd__nand2_2 _28914_ (.A(_05763_),
    .B(_05896_),
    .Y(_06893_));
 sky130_fd_sc_hd__o21ai_2 _28915_ (.A1(_06890_),
    .A2(_06892_),
    .B1(_06893_),
    .Y(_06894_));
 sky130_fd_sc_hd__inv_2 _28916_ (.A(_06893_),
    .Y(_06895_));
 sky130_fd_sc_hd__buf_1 _28917_ (.A(_19382_),
    .X(_06896_));
 sky130_fd_sc_hd__a22o_2 _28918_ (.A1(_05857_),
    .A2(_19609_),
    .B1(_06896_),
    .B2(_06540_),
    .X(_06897_));
 sky130_fd_sc_hd__o211ai_2 _28919_ (.A1(_06688_),
    .A2(_06891_),
    .B1(_06895_),
    .C1(_06897_),
    .Y(_06898_));
 sky130_fd_sc_hd__o22ai_2 _28920_ (.A1(_06807_),
    .A2(_06809_),
    .B1(_06811_),
    .B2(_06814_),
    .Y(_06899_));
 sky130_fd_sc_hd__nand3_2 _28921_ (.A(_06894_),
    .B(_06898_),
    .C(_06899_),
    .Y(_06900_));
 sky130_fd_sc_hd__o21ai_2 _28922_ (.A1(_06890_),
    .A2(_06892_),
    .B1(_06895_),
    .Y(_06901_));
 sky130_fd_sc_hd__a21oi_2 _28923_ (.A1(_06812_),
    .A2(_06815_),
    .B1(_06810_),
    .Y(_06902_));
 sky130_fd_sc_hd__o211ai_2 _28924_ (.A1(_06688_),
    .A2(_06891_),
    .B1(_06893_),
    .C1(_06897_),
    .Y(_06903_));
 sky130_fd_sc_hd__nand3_2 _28925_ (.A(_06901_),
    .B(_06902_),
    .C(_06903_),
    .Y(_06904_));
 sky130_fd_sc_hd__nor2_2 _28926_ (.A(_06698_),
    .B(_06692_),
    .Y(_06905_));
 sky130_fd_sc_hd__o2bb2ai_2 _28927_ (.A1_N(_06900_),
    .A2_N(_06904_),
    .B1(_06689_),
    .B2(_06905_),
    .Y(_06906_));
 sky130_fd_sc_hd__nor2_2 _28928_ (.A(_06689_),
    .B(_06905_),
    .Y(_06907_));
 sky130_fd_sc_hd__nand3_2 _28929_ (.A(_06904_),
    .B(_06900_),
    .C(_06907_),
    .Y(_06908_));
 sky130_fd_sc_hd__o21a_2 _28930_ (.A1(_06791_),
    .A2(_06795_),
    .B1(_06796_),
    .X(_06909_));
 sky130_fd_sc_hd__nand2_2 _28931_ (.A(_06799_),
    .B(_06797_),
    .Y(_06910_));
 sky130_fd_sc_hd__and2_2 _28932_ (.A(_06802_),
    .B(_06633_),
    .X(_06911_));
 sky130_fd_sc_hd__o21ai_2 _28933_ (.A1(_06791_),
    .A2(_06910_),
    .B1(_06911_),
    .Y(_06912_));
 sky130_fd_sc_hd__o2bb2ai_2 _28934_ (.A1_N(_06805_),
    .A2_N(_06817_),
    .B1(_06909_),
    .B2(_06912_),
    .Y(_06913_));
 sky130_fd_sc_hd__a21oi_2 _28935_ (.A1(_06906_),
    .A2(_06908_),
    .B1(_06913_),
    .Y(_06914_));
 sky130_fd_sc_hd__and3_2 _28936_ (.A(_06894_),
    .B(_06898_),
    .C(_06899_),
    .X(_06915_));
 sky130_fd_sc_hd__nand2_2 _28937_ (.A(_06904_),
    .B(_06907_),
    .Y(_06916_));
 sky130_fd_sc_hd__o211a_2 _28938_ (.A1(_06915_),
    .A2(_06916_),
    .B1(_06906_),
    .C1(_06913_),
    .X(_06917_));
 sky130_fd_sc_hd__o22ai_2 _28939_ (.A1(_06887_),
    .A2(_06888_),
    .B1(_06914_),
    .B2(_06917_),
    .Y(_06918_));
 sky130_fd_sc_hd__nand2_2 _28940_ (.A(_06906_),
    .B(_06908_),
    .Y(_06919_));
 sky130_fd_sc_hd__o2bb2a_2 _28941_ (.A1_N(_06805_),
    .A2_N(_06817_),
    .B1(_06909_),
    .B2(_06912_),
    .X(_06920_));
 sky130_fd_sc_hd__nand2_2 _28942_ (.A(_06919_),
    .B(_06920_),
    .Y(_06921_));
 sky130_fd_sc_hd__nand3_2 _28943_ (.A(_06913_),
    .B(_06906_),
    .C(_06908_),
    .Y(_06922_));
 sky130_fd_sc_hd__nand2_2 _28944_ (.A(_06710_),
    .B(_06702_),
    .Y(_06923_));
 sky130_fd_sc_hd__nand3_2 _28945_ (.A(_06921_),
    .B(_06922_),
    .C(_06923_),
    .Y(_06924_));
 sky130_fd_sc_hd__a22oi_2 _28946_ (.A1(_06718_),
    .A2(_06886_),
    .B1(_06918_),
    .B2(_06924_),
    .Y(_06925_));
 sky130_fd_sc_hd__nor2_2 _28947_ (.A(_06885_),
    .B(_06713_),
    .Y(_06926_));
 sky130_fd_sc_hd__o211a_2 _28948_ (.A1(_06716_),
    .A2(_06926_),
    .B1(_06924_),
    .C1(_06918_),
    .X(_06927_));
 sky130_fd_sc_hd__o21ai_2 _28949_ (.A1(_06729_),
    .A2(_06725_),
    .B1(_06734_),
    .Y(_06928_));
 sky130_fd_sc_hd__nand2_2 _28950_ (.A(_19387_),
    .B(\pcpi_mul.rs1[13] ),
    .Y(_06929_));
 sky130_fd_sc_hd__nand2_2 _28951_ (.A(_19390_),
    .B(_06205_),
    .Y(_06930_));
 sky130_fd_sc_hd__or2_2 _28952_ (.A(_06929_),
    .B(_06930_),
    .X(_06931_));
 sky130_fd_sc_hd__nand2_2 _28953_ (.A(_06929_),
    .B(_06930_),
    .Y(_06932_));
 sky130_fd_sc_hd__nand2_2 _28954_ (.A(_05157_),
    .B(\pcpi_mul.rs1[18] ),
    .Y(_06933_));
 sky130_fd_sc_hd__nand3_2 _28955_ (.A(_06931_),
    .B(_06932_),
    .C(_06933_),
    .Y(_06934_));
 sky130_fd_sc_hd__buf_1 _28956_ (.A(_06387_),
    .X(_06935_));
 sky130_fd_sc_hd__a22oi_2 _28957_ (.A1(_06735_),
    .A2(_06736_),
    .B1(_05403_),
    .B2(_06935_),
    .Y(_06936_));
 sky130_fd_sc_hd__nor2_2 _28958_ (.A(_06929_),
    .B(_06930_),
    .Y(_06937_));
 sky130_fd_sc_hd__inv_2 _28959_ (.A(_06933_),
    .Y(_06938_));
 sky130_fd_sc_hd__o21ai_2 _28960_ (.A1(_06936_),
    .A2(_06937_),
    .B1(_06938_),
    .Y(_06939_));
 sky130_fd_sc_hd__nand3b_2 _28961_ (.A_N(_06928_),
    .B(_06934_),
    .C(_06939_),
    .Y(_06940_));
 sky130_fd_sc_hd__nand2_2 _28962_ (.A(_06938_),
    .B(_06932_),
    .Y(_06941_));
 sky130_fd_sc_hd__o21ai_2 _28963_ (.A1(_06936_),
    .A2(_06937_),
    .B1(_06933_),
    .Y(_06942_));
 sky130_fd_sc_hd__o211ai_2 _28964_ (.A1(_06937_),
    .A2(_06941_),
    .B1(_06928_),
    .C1(_06942_),
    .Y(_06943_));
 sky130_fd_sc_hd__buf_1 _28965_ (.A(\pcpi_mul.rs1[17] ),
    .X(_06944_));
 sky130_fd_sc_hd__buf_1 _28966_ (.A(_06944_),
    .X(_06945_));
 sky130_fd_sc_hd__buf_1 _28967_ (.A(\pcpi_mul.rs1[16] ),
    .X(_06946_));
 sky130_fd_sc_hd__nand2_2 _28968_ (.A(_05268_),
    .B(_06946_),
    .Y(_06947_));
 sky130_fd_sc_hd__a21o_2 _28969_ (.A1(_05909_),
    .A2(_06945_),
    .B1(_06947_),
    .X(_06948_));
 sky130_fd_sc_hd__buf_1 _28970_ (.A(\pcpi_mul.rs1[16] ),
    .X(_06949_));
 sky130_fd_sc_hd__buf_1 _28971_ (.A(_06949_),
    .X(_06950_));
 sky130_fd_sc_hd__buf_1 _28972_ (.A(\pcpi_mul.rs1[17] ),
    .X(_06951_));
 sky130_fd_sc_hd__nand2_2 _28973_ (.A(_05221_),
    .B(_06951_),
    .Y(_06952_));
 sky130_fd_sc_hd__a21o_2 _28974_ (.A1(_19398_),
    .A2(_06950_),
    .B1(_06952_),
    .X(_06953_));
 sky130_fd_sc_hd__buf_1 _28975_ (.A(_06373_),
    .X(_06954_));
 sky130_fd_sc_hd__nand2_2 _28976_ (.A(_19394_),
    .B(_06954_),
    .Y(_06955_));
 sky130_fd_sc_hd__a21oi_2 _28977_ (.A1(_06948_),
    .A2(_06953_),
    .B1(_06955_),
    .Y(_06956_));
 sky130_fd_sc_hd__buf_1 _28978_ (.A(_06372_),
    .X(_06957_));
 sky130_fd_sc_hd__inv_2 _28979_ (.A(_06957_),
    .Y(_06958_));
 sky130_fd_sc_hd__buf_1 _28980_ (.A(_06958_),
    .X(_06959_));
 sky130_fd_sc_hd__o211a_2 _28981_ (.A1(_05150_),
    .A2(_06959_),
    .B1(_06953_),
    .C1(_06948_),
    .X(_06960_));
 sky130_fd_sc_hd__nor2_2 _28982_ (.A(_06956_),
    .B(_06960_),
    .Y(_06961_));
 sky130_fd_sc_hd__a21oi_2 _28983_ (.A1(_06940_),
    .A2(_06943_),
    .B1(_06961_),
    .Y(_06962_));
 sky130_fd_sc_hd__o21a_2 _28984_ (.A1(_06936_),
    .A2(_06937_),
    .B1(_06933_),
    .X(_06963_));
 sky130_fd_sc_hd__o21ai_2 _28985_ (.A1(_06937_),
    .A2(_06941_),
    .B1(_06928_),
    .Y(_06964_));
 sky130_fd_sc_hd__o211a_2 _28986_ (.A1(_06963_),
    .A2(_06964_),
    .B1(_06940_),
    .C1(_06961_),
    .X(_06965_));
 sky130_fd_sc_hd__nand2_2 _28987_ (.A(_06756_),
    .B(_06745_),
    .Y(_06966_));
 sky130_fd_sc_hd__nand2_2 _28988_ (.A(_06966_),
    .B(_06741_),
    .Y(_06967_));
 sky130_fd_sc_hd__o21bai_2 _28989_ (.A1(_06962_),
    .A2(_06965_),
    .B1_N(_06967_),
    .Y(_06968_));
 sky130_fd_sc_hd__nor2_2 _28990_ (.A(_06963_),
    .B(_06964_),
    .Y(_06969_));
 sky130_fd_sc_hd__nand2_2 _28991_ (.A(_06961_),
    .B(_06940_),
    .Y(_06970_));
 sky130_fd_sc_hd__a21o_2 _28992_ (.A1(_06940_),
    .A2(_06943_),
    .B1(_06961_),
    .X(_06971_));
 sky130_fd_sc_hd__o211ai_2 _28993_ (.A1(_06969_),
    .A2(_06970_),
    .B1(_06967_),
    .C1(_06971_),
    .Y(_06972_));
 sky130_fd_sc_hd__a41o_2 _28994_ (.A1(_19399_),
    .A2(_19402_),
    .A3(_19591_),
    .A4(_19595_),
    .B1(_06754_),
    .X(_06973_));
 sky130_fd_sc_hd__a21oi_2 _28995_ (.A1(_06968_),
    .A2(_06972_),
    .B1(_06973_),
    .Y(_06974_));
 sky130_fd_sc_hd__nand2_2 _28996_ (.A(_06971_),
    .B(_06967_),
    .Y(_06975_));
 sky130_fd_sc_hd__o211a_2 _28997_ (.A1(_06965_),
    .A2(_06975_),
    .B1(_06973_),
    .C1(_06968_),
    .X(_06976_));
 sky130_fd_sc_hd__nor2_2 _28998_ (.A(_06974_),
    .B(_06976_),
    .Y(_06977_));
 sky130_fd_sc_hd__o21ai_2 _28999_ (.A1(_06925_),
    .A2(_06927_),
    .B1(_06977_),
    .Y(_06978_));
 sky130_fd_sc_hd__a21o_2 _29000_ (.A1(_06968_),
    .A2(_06972_),
    .B1(_06973_),
    .X(_06979_));
 sky130_fd_sc_hd__nand3_2 _29001_ (.A(_06968_),
    .B(_06972_),
    .C(_06973_),
    .Y(_06980_));
 sky130_fd_sc_hd__nand2_2 _29002_ (.A(_06979_),
    .B(_06980_),
    .Y(_06981_));
 sky130_fd_sc_hd__inv_2 _29003_ (.A(_06886_),
    .Y(_06982_));
 sky130_fd_sc_hd__o2bb2ai_2 _29004_ (.A1_N(_06924_),
    .A2_N(_06918_),
    .B1(_06713_),
    .B2(_06982_),
    .Y(_06983_));
 sky130_fd_sc_hd__o211ai_2 _29005_ (.A1(_06716_),
    .A2(_06926_),
    .B1(_06924_),
    .C1(_06918_),
    .Y(_06984_));
 sky130_fd_sc_hd__nand3_2 _29006_ (.A(_06981_),
    .B(_06983_),
    .C(_06984_),
    .Y(_06985_));
 sky130_fd_sc_hd__nand3_2 _29007_ (.A(_06978_),
    .B(_06842_),
    .C(_06985_),
    .Y(_06986_));
 sky130_fd_sc_hd__o22ai_2 _29008_ (.A1(_06976_),
    .A2(_06974_),
    .B1(_06925_),
    .B2(_06927_),
    .Y(_06987_));
 sky130_fd_sc_hd__nand3_2 _29009_ (.A(_06977_),
    .B(_06983_),
    .C(_06984_),
    .Y(_06988_));
 sky130_fd_sc_hd__nand3_2 _29010_ (.A(_06987_),
    .B(_06851_),
    .C(_06988_),
    .Y(_06989_));
 sky130_fd_sc_hd__nor2_2 _29011_ (.A(_06770_),
    .B(_06723_),
    .Y(_06990_));
 sky130_fd_sc_hd__nor2_2 _29012_ (.A(_06722_),
    .B(_06990_),
    .Y(_06991_));
 sky130_fd_sc_hd__nand3_2 _29013_ (.A(_06986_),
    .B(_06989_),
    .C(_06991_),
    .Y(_06992_));
 sky130_fd_sc_hd__buf_1 _29014_ (.A(_06992_),
    .X(_06993_));
 sky130_fd_sc_hd__o2bb2ai_2 _29015_ (.A1_N(_06989_),
    .A2_N(_06986_),
    .B1(_06722_),
    .B2(_06990_),
    .Y(_06994_));
 sky130_fd_sc_hd__a21oi_2 _29016_ (.A1(_06830_),
    .A2(_06832_),
    .B1(_06825_),
    .Y(_06995_));
 sky130_fd_sc_hd__and4_2 _29017_ (.A(_06821_),
    .B(_06823_),
    .C(_05248_),
    .D(_19635_),
    .X(_06996_));
 sky130_fd_sc_hd__inv_2 _29018_ (.A(_06996_),
    .Y(_06997_));
 sky130_fd_sc_hd__inv_2 _29019_ (.A(_06823_),
    .Y(_06998_));
 sky130_fd_sc_hd__nand2_2 _29020_ (.A(_19354_),
    .B(_05190_),
    .Y(_06999_));
 sky130_fd_sc_hd__o21ai_2 _29021_ (.A1(_06998_),
    .A2(_05256_),
    .B1(_06999_),
    .Y(_07000_));
 sky130_fd_sc_hd__nor2_2 _29022_ (.A(_06831_),
    .B(_05319_),
    .Y(_07001_));
 sky130_fd_sc_hd__nand3_2 _29023_ (.A(_06997_),
    .B(_07000_),
    .C(_07001_),
    .Y(_07002_));
 sky130_fd_sc_hd__o21a_2 _29024_ (.A1(_06998_),
    .A2(_05256_),
    .B1(_06999_),
    .X(_07003_));
 sky130_fd_sc_hd__inv_2 _29025_ (.A(_07001_),
    .Y(_07004_));
 sky130_fd_sc_hd__o21ai_2 _29026_ (.A1(_06996_),
    .A2(_07003_),
    .B1(_07004_),
    .Y(_07005_));
 sky130_fd_sc_hd__nand3b_2 _29027_ (.A_N(_06995_),
    .B(_07002_),
    .C(_07005_),
    .Y(_07006_));
 sky130_fd_sc_hd__nor2_2 _29028_ (.A(_06832_),
    .B(_06825_),
    .Y(_07007_));
 sky130_fd_sc_hd__o2bb2ai_2 _29029_ (.A1_N(_07002_),
    .A2_N(_07005_),
    .B1(_06834_),
    .B2(_07007_),
    .Y(_07008_));
 sky130_fd_sc_hd__o2bb2ai_2 _29030_ (.A1_N(_07006_),
    .A2_N(_07008_),
    .B1(_06602_),
    .B2(_06836_),
    .Y(_07009_));
 sky130_fd_sc_hd__nor2_2 _29031_ (.A(_06602_),
    .B(_06836_),
    .Y(_07010_));
 sky130_fd_sc_hd__nand3_2 _29032_ (.A(_07010_),
    .B(_07006_),
    .C(_07008_),
    .Y(_07011_));
 sky130_fd_sc_hd__buf_1 _29033_ (.A(_06269_),
    .X(_07012_));
 sky130_fd_sc_hd__a22oi_2 _29034_ (.A1(_07012_),
    .A2(_05338_),
    .B1(_06276_),
    .B2(_05765_),
    .Y(_07013_));
 sky130_fd_sc_hd__nand2_2 _29035_ (.A(_06624_),
    .B(_05206_),
    .Y(_07014_));
 sky130_fd_sc_hd__buf_1 _29036_ (.A(\pcpi_mul.rs2[13] ),
    .X(_07015_));
 sky130_fd_sc_hd__nand2_2 _29037_ (.A(_07015_),
    .B(_05340_),
    .Y(_07016_));
 sky130_fd_sc_hd__nor2_2 _29038_ (.A(_07014_),
    .B(_07016_),
    .Y(_07017_));
 sky130_fd_sc_hd__and2_2 _29039_ (.A(_19367_),
    .B(_05347_),
    .X(_07018_));
 sky130_fd_sc_hd__o21ai_2 _29040_ (.A1(_07013_),
    .A2(_07017_),
    .B1(_07018_),
    .Y(_07019_));
 sky130_fd_sc_hd__buf_1 _29041_ (.A(_06275_),
    .X(_07020_));
 sky130_fd_sc_hd__nand3_2 _29042_ (.A(_19363_),
    .B(_07020_),
    .C(_05338_),
    .Y(_07021_));
 sky130_fd_sc_hd__nand2_2 _29043_ (.A(_07014_),
    .B(_07016_),
    .Y(_07022_));
 sky130_fd_sc_hd__o221ai_2 _29044_ (.A1(_06118_),
    .A2(_05261_),
    .B1(_05856_),
    .B2(_07021_),
    .C1(_07022_),
    .Y(_07023_));
 sky130_fd_sc_hd__o21ai_2 _29045_ (.A1(_06793_),
    .A2(_06794_),
    .B1(_06796_),
    .Y(_07024_));
 sky130_fd_sc_hd__nand2_2 _29046_ (.A(_07024_),
    .B(_06800_),
    .Y(_07025_));
 sky130_fd_sc_hd__a21o_2 _29047_ (.A1(_07019_),
    .A2(_07023_),
    .B1(_07025_),
    .X(_07026_));
 sky130_fd_sc_hd__nand3_2 _29048_ (.A(_07019_),
    .B(_07025_),
    .C(_07023_),
    .Y(_07027_));
 sky130_fd_sc_hd__a22oi_2 _29049_ (.A1(_05800_),
    .A2(_05502_),
    .B1(_05958_),
    .B2(_05506_),
    .Y(_07028_));
 sky130_fd_sc_hd__nand2_2 _29050_ (.A(\pcpi_mul.rs2[11] ),
    .B(\pcpi_mul.rs1[7] ),
    .Y(_07029_));
 sky130_fd_sc_hd__nand2_2 _29051_ (.A(_19372_),
    .B(_19615_),
    .Y(_07030_));
 sky130_fd_sc_hd__nor2_2 _29052_ (.A(_07029_),
    .B(_07030_),
    .Y(_07031_));
 sky130_fd_sc_hd__nand2_2 _29053_ (.A(_05672_),
    .B(_05614_),
    .Y(_07032_));
 sky130_fd_sc_hd__o21bai_2 _29054_ (.A1(_07028_),
    .A2(_07031_),
    .B1_N(_07032_),
    .Y(_07033_));
 sky130_fd_sc_hd__buf_1 _29055_ (.A(_19372_),
    .X(_07034_));
 sky130_fd_sc_hd__nand3b_2 _29056_ (.A_N(_07029_),
    .B(_07034_),
    .C(_06507_),
    .Y(_07035_));
 sky130_fd_sc_hd__nand2_2 _29057_ (.A(_07029_),
    .B(_07030_),
    .Y(_07036_));
 sky130_fd_sc_hd__nand3_2 _29058_ (.A(_07035_),
    .B(_07032_),
    .C(_07036_),
    .Y(_07037_));
 sky130_fd_sc_hd__nand2_2 _29059_ (.A(_07033_),
    .B(_07037_),
    .Y(_07038_));
 sky130_fd_sc_hd__a21o_2 _29060_ (.A1(_07026_),
    .A2(_07027_),
    .B1(_07038_),
    .X(_07039_));
 sky130_fd_sc_hd__a32oi_2 _29061_ (.A1(_07019_),
    .A2(_07025_),
    .A3(_07023_),
    .B1(_07033_),
    .B2(_07037_),
    .Y(_07040_));
 sky130_fd_sc_hd__nand2_2 _29062_ (.A(_07040_),
    .B(_07026_),
    .Y(_07041_));
 sky130_fd_sc_hd__nand2_2 _29063_ (.A(_07039_),
    .B(_07041_),
    .Y(_07042_));
 sky130_fd_sc_hd__a21o_2 _29064_ (.A1(_07009_),
    .A2(_07011_),
    .B1(_07042_),
    .X(_07043_));
 sky130_fd_sc_hd__nand3_2 _29065_ (.A(_07042_),
    .B(_07009_),
    .C(_07011_),
    .Y(_07044_));
 sky130_fd_sc_hd__nand3_2 _29066_ (.A(_07043_),
    .B(_07044_),
    .C(_06840_),
    .Y(_07045_));
 sky130_fd_sc_hd__a22o_2 _29067_ (.A1(_07041_),
    .A2(_07039_),
    .B1(_07009_),
    .B2(_07011_),
    .X(_07046_));
 sky130_fd_sc_hd__a22oi_2 _29068_ (.A1(_06818_),
    .A2(_06819_),
    .B1(_06837_),
    .B2(_06838_),
    .Y(_07047_));
 sky130_fd_sc_hd__a21oi_2 _29069_ (.A1(_07019_),
    .A2(_07023_),
    .B1(_07025_),
    .Y(_07048_));
 sky130_fd_sc_hd__nand2_2 _29070_ (.A(_07027_),
    .B(_07038_),
    .Y(_07049_));
 sky130_fd_sc_hd__o2111ai_2 _29071_ (.A1(_07048_),
    .A2(_07049_),
    .B1(_07039_),
    .C1(_07011_),
    .D1(_07009_),
    .Y(_07050_));
 sky130_fd_sc_hd__nand3_2 _29072_ (.A(_07046_),
    .B(_07047_),
    .C(_07050_),
    .Y(_07051_));
 sky130_fd_sc_hd__inv_2 _29073_ (.A(\pcpi_mul.rs2[18] ),
    .Y(_07052_));
 sky130_fd_sc_hd__buf_1 _29074_ (.A(_07052_),
    .X(_07053_));
 sky130_fd_sc_hd__nor2_2 _29075_ (.A(_07053_),
    .B(_04840_),
    .Y(_07054_));
 sky130_fd_sc_hd__nand3_2 _29076_ (.A(_07045_),
    .B(_07051_),
    .C(_07054_),
    .Y(_07055_));
 sky130_fd_sc_hd__inv_2 _29077_ (.A(_07055_),
    .Y(_07056_));
 sky130_fd_sc_hd__nand2_2 _29078_ (.A(_07045_),
    .B(_07051_),
    .Y(_07057_));
 sky130_fd_sc_hd__inv_2 _29079_ (.A(_07054_),
    .Y(_07058_));
 sky130_fd_sc_hd__nand2_2 _29080_ (.A(_07057_),
    .B(_07058_),
    .Y(_07059_));
 sky130_fd_sc_hd__inv_2 _29081_ (.A(_07059_),
    .Y(_07060_));
 sky130_fd_sc_hd__o2bb2ai_2 _29082_ (.A1_N(_06993_),
    .A2_N(_06994_),
    .B1(_07056_),
    .B2(_07060_),
    .Y(_07061_));
 sky130_fd_sc_hd__nand2_2 _29083_ (.A(_07059_),
    .B(_07055_),
    .Y(_07062_));
 sky130_fd_sc_hd__inv_2 _29084_ (.A(_07062_),
    .Y(_07063_));
 sky130_fd_sc_hd__nand3_2 _29085_ (.A(_06994_),
    .B(_07063_),
    .C(_06993_),
    .Y(_07064_));
 sky130_fd_sc_hd__a21oi_2 _29086_ (.A1(_07061_),
    .A2(_07064_),
    .B1(_06858_),
    .Y(_07065_));
 sky130_fd_sc_hd__a21oi_2 _29087_ (.A1(_06986_),
    .A2(_06989_),
    .B1(_06991_),
    .Y(_07066_));
 sky130_fd_sc_hd__nand2_2 _29088_ (.A(_06993_),
    .B(_07063_),
    .Y(_07067_));
 sky130_fd_sc_hd__o211a_2 _29089_ (.A1(_07066_),
    .A2(_07067_),
    .B1(_06858_),
    .C1(_07061_),
    .X(_07068_));
 sky130_fd_sc_hd__o22ai_2 _29090_ (.A1(_06883_),
    .A2(_06884_),
    .B1(_07065_),
    .B2(_07068_),
    .Y(_07069_));
 sky130_fd_sc_hd__a21oi_2 _29091_ (.A1(_06859_),
    .A2(_06860_),
    .B1(_06850_),
    .Y(_07070_));
 sky130_fd_sc_hd__nand2_2 _29092_ (.A(_06994_),
    .B(_06993_),
    .Y(_07071_));
 sky130_fd_sc_hd__a21oi_2 _29093_ (.A1(_07071_),
    .A2(_07062_),
    .B1(_06855_),
    .Y(_07072_));
 sky130_fd_sc_hd__nand2_2 _29094_ (.A(_07072_),
    .B(_07064_),
    .Y(_07073_));
 sky130_fd_sc_hd__a21o_2 _29095_ (.A1(_06789_),
    .A2(_06784_),
    .B1(_06880_),
    .X(_07074_));
 sky130_fd_sc_hd__nand3_2 _29096_ (.A(_06789_),
    .B(_06784_),
    .C(_06880_),
    .Y(_07075_));
 sky130_fd_sc_hd__nand2_2 _29097_ (.A(_07074_),
    .B(_07075_),
    .Y(_07076_));
 sky130_fd_sc_hd__a22oi_2 _29098_ (.A1(_07055_),
    .A2(_07059_),
    .B1(_06994_),
    .B2(_06993_),
    .Y(_07077_));
 sky130_fd_sc_hd__nor2_2 _29099_ (.A(_07066_),
    .B(_07067_),
    .Y(_07078_));
 sky130_fd_sc_hd__o22ai_2 _29100_ (.A1(_06847_),
    .A2(_06848_),
    .B1(_07077_),
    .B2(_07078_),
    .Y(_07079_));
 sky130_fd_sc_hd__nand3_2 _29101_ (.A(_07073_),
    .B(_07076_),
    .C(_07079_),
    .Y(_07080_));
 sky130_fd_sc_hd__nand3_2 _29102_ (.A(_07069_),
    .B(_07070_),
    .C(_07080_),
    .Y(_07081_));
 sky130_fd_sc_hd__nand2_2 _29103_ (.A(_07081_),
    .B(_06682_),
    .Y(_07082_));
 sky130_fd_sc_hd__o21ai_2 _29104_ (.A1(_07065_),
    .A2(_07068_),
    .B1(_07076_),
    .Y(_07083_));
 sky130_fd_sc_hd__o21ai_2 _29105_ (.A1(_06868_),
    .A2(_06856_),
    .B1(_06861_),
    .Y(_07084_));
 sky130_fd_sc_hd__and2_2 _29106_ (.A(_07074_),
    .B(_07075_),
    .X(_07085_));
 sky130_fd_sc_hd__nand3_2 _29107_ (.A(_07073_),
    .B(_07085_),
    .C(_07079_),
    .Y(_07086_));
 sky130_fd_sc_hd__nand3_2 _29108_ (.A(_07083_),
    .B(_07084_),
    .C(_07086_),
    .Y(_07087_));
 sky130_fd_sc_hd__nand2_2 _29109_ (.A(_07087_),
    .B(_07081_),
    .Y(_07088_));
 sky130_fd_sc_hd__inv_2 _29110_ (.A(_06682_),
    .Y(_07089_));
 sky130_fd_sc_hd__a22oi_2 _29111_ (.A1(_06873_),
    .A2(_06865_),
    .B1(_07088_),
    .B2(_07089_),
    .Y(_07090_));
 sky130_fd_sc_hd__o2bb2ai_2 _29112_ (.A1_N(_07081_),
    .A2_N(_07087_),
    .B1(_06597_),
    .B2(_06681_),
    .Y(_07091_));
 sky130_fd_sc_hd__nand2_2 _29113_ (.A(_06873_),
    .B(_06865_),
    .Y(_07092_));
 sky130_fd_sc_hd__a21oi_2 _29114_ (.A1(_07091_),
    .A2(_07082_),
    .B1(_07092_),
    .Y(_07093_));
 sky130_fd_sc_hd__a21oi_2 _29115_ (.A1(_07082_),
    .A2(_07090_),
    .B1(_07093_),
    .Y(_07094_));
 sky130_fd_sc_hd__a31oi_2 _29116_ (.A1(_06679_),
    .A2(_06677_),
    .A3(_06876_),
    .B1(_06875_),
    .Y(_07095_));
 sky130_fd_sc_hd__or2_2 _29117_ (.A(_07094_),
    .B(_07095_),
    .X(_07096_));
 sky130_fd_sc_hd__nand2_2 _29118_ (.A(_07095_),
    .B(_07094_),
    .Y(_07097_));
 sky130_fd_sc_hd__and2_2 _29119_ (.A(_07096_),
    .B(_07097_),
    .X(_02637_));
 sky130_fd_sc_hd__and2_2 _29120_ (.A(_06710_),
    .B(_06702_),
    .X(_07098_));
 sky130_fd_sc_hd__nand2_2 _29121_ (.A(_06922_),
    .B(_07098_),
    .Y(_07099_));
 sky130_fd_sc_hd__inv_2 _29122_ (.A(_06904_),
    .Y(_07100_));
 sky130_fd_sc_hd__nor2_2 _29123_ (.A(_06907_),
    .B(_06915_),
    .Y(_07101_));
 sky130_fd_sc_hd__a22oi_2 _29124_ (.A1(_06008_),
    .A2(_06539_),
    .B1(_06010_),
    .B2(_19602_),
    .Y(_07102_));
 sky130_fd_sc_hd__nand3_2 _29125_ (.A(_05447_),
    .B(_19382_),
    .C(\pcpi_mul.rs1[11] ),
    .Y(_07103_));
 sky130_fd_sc_hd__nor2_2 _29126_ (.A(_06390_),
    .B(_07103_),
    .Y(_07104_));
 sky130_fd_sc_hd__nand2_2 _29127_ (.A(_05763_),
    .B(\pcpi_mul.rs1[13] ),
    .Y(_07105_));
 sky130_fd_sc_hd__o21ai_2 _29128_ (.A1(_07102_),
    .A2(_07104_),
    .B1(_07105_),
    .Y(_07106_));
 sky130_fd_sc_hd__o21ai_2 _29129_ (.A1(_07032_),
    .A2(_07028_),
    .B1(_07035_),
    .Y(_07107_));
 sky130_fd_sc_hd__inv_2 _29130_ (.A(_07105_),
    .Y(_07108_));
 sky130_fd_sc_hd__buf_1 _29131_ (.A(\pcpi_mul.rs1[12] ),
    .X(_07109_));
 sky130_fd_sc_hd__a22o_2 _29132_ (.A1(_05639_),
    .A2(_06539_),
    .B1(_05641_),
    .B2(_07109_),
    .X(_07110_));
 sky130_fd_sc_hd__o211ai_2 _29133_ (.A1(_06390_),
    .A2(_07103_),
    .B1(_07108_),
    .C1(_07110_),
    .Y(_07111_));
 sky130_fd_sc_hd__nand3_2 _29134_ (.A(_07106_),
    .B(_07107_),
    .C(_07111_),
    .Y(_07112_));
 sky130_fd_sc_hd__o21ai_2 _29135_ (.A1(_07102_),
    .A2(_07104_),
    .B1(_07108_),
    .Y(_07113_));
 sky130_fd_sc_hd__o21ai_2 _29136_ (.A1(_07029_),
    .A2(_07030_),
    .B1(_07032_),
    .Y(_07114_));
 sky130_fd_sc_hd__nand2_2 _29137_ (.A(_07114_),
    .B(_07036_),
    .Y(_07115_));
 sky130_fd_sc_hd__o211ai_2 _29138_ (.A1(_06390_),
    .A2(_07103_),
    .B1(_07105_),
    .C1(_07110_),
    .Y(_07116_));
 sky130_fd_sc_hd__nand3_2 _29139_ (.A(_07113_),
    .B(_07115_),
    .C(_07116_),
    .Y(_07117_));
 sky130_fd_sc_hd__nor2_2 _29140_ (.A(_06895_),
    .B(_06892_),
    .Y(_07118_));
 sky130_fd_sc_hd__o2bb2ai_2 _29141_ (.A1_N(_07112_),
    .A2_N(_07117_),
    .B1(_06890_),
    .B2(_07118_),
    .Y(_07119_));
 sky130_fd_sc_hd__nor2_2 _29142_ (.A(_06890_),
    .B(_07118_),
    .Y(_07120_));
 sky130_fd_sc_hd__nand3_2 _29143_ (.A(_07112_),
    .B(_07117_),
    .C(_07120_),
    .Y(_07121_));
 sky130_fd_sc_hd__nand2_2 _29144_ (.A(_07049_),
    .B(_07026_),
    .Y(_07122_));
 sky130_fd_sc_hd__a21oi_2 _29145_ (.A1(_07119_),
    .A2(_07121_),
    .B1(_07122_),
    .Y(_07123_));
 sky130_fd_sc_hd__o211a_2 _29146_ (.A1(_07048_),
    .A2(_07040_),
    .B1(_07121_),
    .C1(_07119_),
    .X(_07124_));
 sky130_fd_sc_hd__o22ai_2 _29147_ (.A1(_07100_),
    .A2(_07101_),
    .B1(_07123_),
    .B2(_07124_),
    .Y(_07125_));
 sky130_fd_sc_hd__a21o_2 _29148_ (.A1(_07119_),
    .A2(_07121_),
    .B1(_07122_),
    .X(_07126_));
 sky130_fd_sc_hd__nand3_2 _29149_ (.A(_07122_),
    .B(_07119_),
    .C(_07121_),
    .Y(_07127_));
 sky130_fd_sc_hd__nand2_2 _29150_ (.A(_06916_),
    .B(_06900_),
    .Y(_07128_));
 sky130_fd_sc_hd__nand3_2 _29151_ (.A(_07126_),
    .B(_07127_),
    .C(_07128_),
    .Y(_07129_));
 sky130_fd_sc_hd__a22oi_2 _29152_ (.A1(_06921_),
    .A2(_07099_),
    .B1(_07125_),
    .B2(_07129_),
    .Y(_07130_));
 sky130_fd_sc_hd__a21oi_2 _29153_ (.A1(_06919_),
    .A2(_06920_),
    .B1(_07098_),
    .Y(_07131_));
 sky130_fd_sc_hd__o211a_2 _29154_ (.A1(_06917_),
    .A2(_07131_),
    .B1(_07129_),
    .C1(_07125_),
    .X(_07132_));
 sky130_fd_sc_hd__a21oi_2 _29155_ (.A1(_06961_),
    .A2(_06940_),
    .B1(_06969_),
    .Y(_07133_));
 sky130_fd_sc_hd__nand2_2 _29156_ (.A(_05321_),
    .B(_19596_),
    .Y(_07134_));
 sky130_fd_sc_hd__nand2_2 _29157_ (.A(_05322_),
    .B(_19593_),
    .Y(_07135_));
 sky130_fd_sc_hd__or2_2 _29158_ (.A(_07134_),
    .B(_07135_),
    .X(_07136_));
 sky130_fd_sc_hd__nand2_2 _29159_ (.A(_07134_),
    .B(_07135_),
    .Y(_07137_));
 sky130_fd_sc_hd__buf_1 _29160_ (.A(\pcpi_mul.rs1[19] ),
    .X(_07138_));
 sky130_fd_sc_hd__nand2_2 _29161_ (.A(_04834_),
    .B(_07138_),
    .Y(_07139_));
 sky130_fd_sc_hd__inv_2 _29162_ (.A(_07139_),
    .Y(_07140_));
 sky130_fd_sc_hd__nand3_2 _29163_ (.A(_07136_),
    .B(_07137_),
    .C(_07140_),
    .Y(_07141_));
 sky130_fd_sc_hd__nand2_2 _29164_ (.A(_06931_),
    .B(_06941_),
    .Y(_07142_));
 sky130_fd_sc_hd__buf_1 _29165_ (.A(_06205_),
    .X(_07143_));
 sky130_fd_sc_hd__a22oi_2 _29166_ (.A1(_06199_),
    .A2(_07143_),
    .B1(_06201_),
    .B2(_06748_),
    .Y(_07144_));
 sky130_fd_sc_hd__nor2_2 _29167_ (.A(_07134_),
    .B(_07135_),
    .Y(_07145_));
 sky130_fd_sc_hd__o21ai_2 _29168_ (.A1(_07144_),
    .A2(_07145_),
    .B1(_07139_),
    .Y(_07146_));
 sky130_fd_sc_hd__nand3_2 _29169_ (.A(_07141_),
    .B(_07142_),
    .C(_07146_),
    .Y(_07147_));
 sky130_fd_sc_hd__nand3_2 _29170_ (.A(_07136_),
    .B(_07137_),
    .C(_07139_),
    .Y(_07148_));
 sky130_fd_sc_hd__a21oi_2 _29171_ (.A1(_06938_),
    .A2(_06932_),
    .B1(_06937_),
    .Y(_07149_));
 sky130_fd_sc_hd__o21ai_2 _29172_ (.A1(_07144_),
    .A2(_07145_),
    .B1(_07140_),
    .Y(_07150_));
 sky130_fd_sc_hd__nand3_2 _29173_ (.A(_07148_),
    .B(_07149_),
    .C(_07150_),
    .Y(_07151_));
 sky130_fd_sc_hd__nand2_2 _29174_ (.A(_07147_),
    .B(_07151_),
    .Y(_07152_));
 sky130_fd_sc_hd__buf_1 _29175_ (.A(_19584_),
    .X(_07153_));
 sky130_fd_sc_hd__nand2_2 _29176_ (.A(_05268_),
    .B(_19588_),
    .Y(_07154_));
 sky130_fd_sc_hd__a21o_2 _29177_ (.A1(_05909_),
    .A2(_07153_),
    .B1(_07154_),
    .X(_07155_));
 sky130_fd_sc_hd__buf_1 _29178_ (.A(_19584_),
    .X(_07156_));
 sky130_fd_sc_hd__nand2_2 _29179_ (.A(_05221_),
    .B(_07156_),
    .Y(_07157_));
 sky130_fd_sc_hd__a21o_2 _29180_ (.A1(_05736_),
    .A2(_06945_),
    .B1(_07157_),
    .X(_07158_));
 sky130_fd_sc_hd__nand2_2 _29181_ (.A(_19393_),
    .B(_06950_),
    .Y(_07159_));
 sky130_fd_sc_hd__a21oi_2 _29182_ (.A1(_07155_),
    .A2(_07158_),
    .B1(_07159_),
    .Y(_07160_));
 sky130_fd_sc_hd__and3_2 _29183_ (.A(_07155_),
    .B(_07158_),
    .C(_07159_),
    .X(_07161_));
 sky130_fd_sc_hd__nor2_2 _29184_ (.A(_07160_),
    .B(_07161_),
    .Y(_07162_));
 sky130_fd_sc_hd__nand2_2 _29185_ (.A(_07152_),
    .B(_07162_),
    .Y(_07163_));
 sky130_fd_sc_hd__a21o_2 _29186_ (.A1(_07155_),
    .A2(_07158_),
    .B1(_07159_),
    .X(_07164_));
 sky130_fd_sc_hd__nand3_2 _29187_ (.A(_07155_),
    .B(_07158_),
    .C(_07159_),
    .Y(_07165_));
 sky130_fd_sc_hd__nand2_2 _29188_ (.A(_07164_),
    .B(_07165_),
    .Y(_07166_));
 sky130_fd_sc_hd__nand3_2 _29189_ (.A(_07166_),
    .B(_07147_),
    .C(_07151_),
    .Y(_07167_));
 sky130_fd_sc_hd__nand3_2 _29190_ (.A(_07133_),
    .B(_07163_),
    .C(_07167_),
    .Y(_07168_));
 sky130_fd_sc_hd__nor2_2 _29191_ (.A(_06947_),
    .B(_06952_),
    .Y(_07169_));
 sky130_fd_sc_hd__nor2_2 _29192_ (.A(_07169_),
    .B(_06956_),
    .Y(_07170_));
 sky130_fd_sc_hd__inv_2 _29193_ (.A(_07170_),
    .Y(_07171_));
 sky130_fd_sc_hd__and2_2 _29194_ (.A(_07168_),
    .B(_07171_),
    .X(_07172_));
 sky130_fd_sc_hd__a21oi_2 _29195_ (.A1(_07141_),
    .A2(_07146_),
    .B1(_07142_),
    .Y(_07173_));
 sky130_fd_sc_hd__nand2_2 _29196_ (.A(_07162_),
    .B(_07147_),
    .Y(_07174_));
 sky130_fd_sc_hd__nand2_2 _29197_ (.A(_07152_),
    .B(_07166_),
    .Y(_07175_));
 sky130_fd_sc_hd__nand2_2 _29198_ (.A(_06970_),
    .B(_06943_),
    .Y(_07176_));
 sky130_fd_sc_hd__o211ai_2 _29199_ (.A1(_07173_),
    .A2(_07174_),
    .B1(_07175_),
    .C1(_07176_),
    .Y(_07177_));
 sky130_fd_sc_hd__a21oi_2 _29200_ (.A1(_07177_),
    .A2(_07168_),
    .B1(_07171_),
    .Y(_07178_));
 sky130_fd_sc_hd__a21oi_2 _29201_ (.A1(_07172_),
    .A2(_07177_),
    .B1(_07178_),
    .Y(_07179_));
 sky130_fd_sc_hd__o21ai_2 _29202_ (.A1(_07130_),
    .A2(_07132_),
    .B1(_07179_),
    .Y(_07180_));
 sky130_fd_sc_hd__nand2_2 _29203_ (.A(_07125_),
    .B(_07129_),
    .Y(_07181_));
 sky130_fd_sc_hd__nand2_2 _29204_ (.A(_07099_),
    .B(_06921_),
    .Y(_07182_));
 sky130_fd_sc_hd__nand2_2 _29205_ (.A(_07181_),
    .B(_07182_),
    .Y(_07183_));
 sky130_fd_sc_hd__nand2_2 _29206_ (.A(_07168_),
    .B(_07171_),
    .Y(_07184_));
 sky130_fd_sc_hd__inv_2 _29207_ (.A(_07177_),
    .Y(_07185_));
 sky130_fd_sc_hd__nand2_2 _29208_ (.A(_07177_),
    .B(_07168_),
    .Y(_07186_));
 sky130_fd_sc_hd__nand2_2 _29209_ (.A(_07186_),
    .B(_07170_),
    .Y(_07187_));
 sky130_fd_sc_hd__o21ai_2 _29210_ (.A1(_07184_),
    .A2(_07185_),
    .B1(_07187_),
    .Y(_07188_));
 sky130_fd_sc_hd__nand3b_2 _29211_ (.A_N(_07182_),
    .B(_07129_),
    .C(_07125_),
    .Y(_07189_));
 sky130_fd_sc_hd__nand3_2 _29212_ (.A(_07183_),
    .B(_07188_),
    .C(_07189_),
    .Y(_07190_));
 sky130_fd_sc_hd__nand3_2 _29213_ (.A(_07180_),
    .B(_07051_),
    .C(_07190_),
    .Y(_07191_));
 sky130_fd_sc_hd__nor2_2 _29214_ (.A(_07170_),
    .B(_07186_),
    .Y(_07192_));
 sky130_fd_sc_hd__o22ai_2 _29215_ (.A1(_07192_),
    .A2(_07178_),
    .B1(_07130_),
    .B2(_07132_),
    .Y(_07193_));
 sky130_fd_sc_hd__inv_2 _29216_ (.A(_07051_),
    .Y(_07194_));
 sky130_fd_sc_hd__nand3_2 _29217_ (.A(_07183_),
    .B(_07179_),
    .C(_07189_),
    .Y(_07195_));
 sky130_fd_sc_hd__nand3_2 _29218_ (.A(_07193_),
    .B(_07194_),
    .C(_07195_),
    .Y(_07196_));
 sky130_fd_sc_hd__buf_1 _29219_ (.A(_07196_),
    .X(_07197_));
 sky130_fd_sc_hd__o21ai_2 _29220_ (.A1(_06925_),
    .A2(_06981_),
    .B1(_06984_),
    .Y(_07198_));
 sky130_fd_sc_hd__a21oi_2 _29221_ (.A1(_07191_),
    .A2(_07197_),
    .B1(_07198_),
    .Y(_07199_));
 sky130_fd_sc_hd__and3_2 _29222_ (.A(_07191_),
    .B(_07197_),
    .C(_07198_),
    .X(_07200_));
 sky130_fd_sc_hd__and3_2 _29223_ (.A(_07010_),
    .B(_07006_),
    .C(_07008_),
    .X(_07201_));
 sky130_fd_sc_hd__a31oi_2 _29224_ (.A1(_07041_),
    .A2(_07009_),
    .A3(_07039_),
    .B1(_07201_),
    .Y(_07202_));
 sky130_fd_sc_hd__buf_1 _29225_ (.A(_05955_),
    .X(_07203_));
 sky130_fd_sc_hd__a22oi_2 _29226_ (.A1(_07203_),
    .A2(_06162_),
    .B1(_06258_),
    .B2(_06492_),
    .Y(_07204_));
 sky130_fd_sc_hd__nand2_2 _29227_ (.A(_05955_),
    .B(_05730_),
    .Y(_07205_));
 sky130_fd_sc_hd__nand2_2 _29228_ (.A(_07034_),
    .B(_06327_),
    .Y(_07206_));
 sky130_fd_sc_hd__nor2_2 _29229_ (.A(_07205_),
    .B(_07206_),
    .Y(_07207_));
 sky130_fd_sc_hd__nand2_2 _29230_ (.A(_05673_),
    .B(_05733_),
    .Y(_07208_));
 sky130_fd_sc_hd__o21bai_2 _29231_ (.A1(_07204_),
    .A2(_07207_),
    .B1_N(_07208_),
    .Y(_07209_));
 sky130_fd_sc_hd__buf_1 _29232_ (.A(_05516_),
    .X(_07210_));
 sky130_fd_sc_hd__nand3b_2 _29233_ (.A_N(_07205_),
    .B(_06605_),
    .C(_07210_),
    .Y(_07211_));
 sky130_fd_sc_hd__nand2_2 _29234_ (.A(_07205_),
    .B(_07206_),
    .Y(_07212_));
 sky130_fd_sc_hd__nand3_2 _29235_ (.A(_07211_),
    .B(_07208_),
    .C(_07212_),
    .Y(_07213_));
 sky130_fd_sc_hd__and2_2 _29236_ (.A(_07209_),
    .B(_07213_),
    .X(_07214_));
 sky130_fd_sc_hd__a21o_2 _29237_ (.A1(_07018_),
    .A2(_07022_),
    .B1(_07017_),
    .X(_07215_));
 sky130_fd_sc_hd__a22oi_2 _29238_ (.A1(_06270_),
    .A2(_05345_),
    .B1(_06272_),
    .B2(_05347_),
    .Y(_07216_));
 sky130_fd_sc_hd__and4_2 _29239_ (.A(_06624_),
    .B(_07015_),
    .C(_06609_),
    .D(_05345_),
    .X(_07217_));
 sky130_fd_sc_hd__nand2_2 _29240_ (.A(_06117_),
    .B(_19618_),
    .Y(_07218_));
 sky130_fd_sc_hd__o21ai_2 _29241_ (.A1(_07216_),
    .A2(_07217_),
    .B1(_07218_),
    .Y(_07219_));
 sky130_fd_sc_hd__nand2_2 _29242_ (.A(_19362_),
    .B(_05193_),
    .Y(_07220_));
 sky130_fd_sc_hd__nand3b_2 _29243_ (.A_N(_07220_),
    .B(_06443_),
    .C(_05422_),
    .Y(_07221_));
 sky130_fd_sc_hd__a22o_2 _29244_ (.A1(_06270_),
    .A2(_05345_),
    .B1(_06272_),
    .B2(_05347_),
    .X(_07222_));
 sky130_fd_sc_hd__inv_2 _29245_ (.A(_07218_),
    .Y(_07223_));
 sky130_fd_sc_hd__nand3_2 _29246_ (.A(_07221_),
    .B(_07222_),
    .C(_07223_),
    .Y(_07224_));
 sky130_fd_sc_hd__nand3_2 _29247_ (.A(_07215_),
    .B(_07219_),
    .C(_07224_),
    .Y(_07225_));
 sky130_fd_sc_hd__o21ai_2 _29248_ (.A1(_07216_),
    .A2(_07217_),
    .B1(_07223_),
    .Y(_07226_));
 sky130_fd_sc_hd__nand3_2 _29249_ (.A(_07221_),
    .B(_07222_),
    .C(_07218_),
    .Y(_07227_));
 sky130_fd_sc_hd__a21oi_2 _29250_ (.A1(_07022_),
    .A2(_07018_),
    .B1(_07017_),
    .Y(_07228_));
 sky130_fd_sc_hd__nand3_2 _29251_ (.A(_07226_),
    .B(_07227_),
    .C(_07228_),
    .Y(_07229_));
 sky130_fd_sc_hd__nand2_2 _29252_ (.A(_07225_),
    .B(_07229_),
    .Y(_07230_));
 sky130_fd_sc_hd__or2_2 _29253_ (.A(_07214_),
    .B(_07230_),
    .X(_07231_));
 sky130_fd_sc_hd__nand2_2 _29254_ (.A(_07230_),
    .B(_07214_),
    .Y(_07232_));
 sky130_fd_sc_hd__nand2_2 _29255_ (.A(_07231_),
    .B(_07232_),
    .Y(_07233_));
 sky130_fd_sc_hd__nand2_2 _29256_ (.A(\pcpi_mul.rs2[17] ),
    .B(_19356_),
    .Y(_07234_));
 sky130_fd_sc_hd__nor2_2 _29257_ (.A(_05147_),
    .B(_07234_),
    .Y(_07235_));
 sky130_fd_sc_hd__buf_1 _29258_ (.A(\pcpi_mul.rs2[17] ),
    .X(_07236_));
 sky130_fd_sc_hd__a22o_2 _29259_ (.A1(_07236_),
    .A2(_19632_),
    .B1(_06823_),
    .B2(_19629_),
    .X(_07237_));
 sky130_fd_sc_hd__inv_2 _29260_ (.A(_07237_),
    .Y(_07238_));
 sky130_fd_sc_hd__nor2_2 _29261_ (.A(_06831_),
    .B(_05849_),
    .Y(_07239_));
 sky130_fd_sc_hd__inv_2 _29262_ (.A(_07239_),
    .Y(_07240_));
 sky130_fd_sc_hd__o21ai_2 _29263_ (.A1(_07235_),
    .A2(_07238_),
    .B1(_07240_),
    .Y(_07241_));
 sky130_fd_sc_hd__a21o_2 _29264_ (.A1(_07000_),
    .A2(_07001_),
    .B1(_06996_),
    .X(_07242_));
 sky130_fd_sc_hd__inv_2 _29265_ (.A(_07235_),
    .Y(_07243_));
 sky130_fd_sc_hd__nand3_2 _29266_ (.A(_07243_),
    .B(_07239_),
    .C(_07237_),
    .Y(_07244_));
 sky130_fd_sc_hd__nand3_2 _29267_ (.A(_07241_),
    .B(_07242_),
    .C(_07244_),
    .Y(_07245_));
 sky130_fd_sc_hd__o21ai_2 _29268_ (.A1(_07235_),
    .A2(_07238_),
    .B1(_07239_),
    .Y(_07246_));
 sky130_fd_sc_hd__a21oi_2 _29269_ (.A1(_07000_),
    .A2(_07001_),
    .B1(_06996_),
    .Y(_07247_));
 sky130_fd_sc_hd__nand3_2 _29270_ (.A(_07240_),
    .B(_07243_),
    .C(_07237_),
    .Y(_07248_));
 sky130_fd_sc_hd__nand3_2 _29271_ (.A(_07246_),
    .B(_07247_),
    .C(_07248_),
    .Y(_07249_));
 sky130_fd_sc_hd__nand2_2 _29272_ (.A(_07245_),
    .B(_07249_),
    .Y(_07250_));
 sky130_fd_sc_hd__nand2_2 _29273_ (.A(_07250_),
    .B(_07006_),
    .Y(_07251_));
 sky130_fd_sc_hd__nand3b_2 _29274_ (.A_N(_07006_),
    .B(_07245_),
    .C(_07249_),
    .Y(_07252_));
 sky130_fd_sc_hd__nand3_2 _29275_ (.A(_07233_),
    .B(_07251_),
    .C(_07252_),
    .Y(_07253_));
 sky130_fd_sc_hd__xor2_2 _29276_ (.A(_07214_),
    .B(_07230_),
    .X(_07254_));
 sky130_fd_sc_hd__nand2_2 _29277_ (.A(_07251_),
    .B(_07252_),
    .Y(_07255_));
 sky130_fd_sc_hd__nand2_2 _29278_ (.A(_07254_),
    .B(_07255_),
    .Y(_07256_));
 sky130_fd_sc_hd__nand3_2 _29279_ (.A(_07202_),
    .B(_07253_),
    .C(_07256_),
    .Y(_07257_));
 sky130_fd_sc_hd__nand2_2 _29280_ (.A(_07233_),
    .B(_07255_),
    .Y(_07258_));
 sky130_fd_sc_hd__nand3_2 _29281_ (.A(_07009_),
    .B(_07041_),
    .C(_07039_),
    .Y(_07259_));
 sky130_fd_sc_hd__nand2_2 _29282_ (.A(_07259_),
    .B(_07011_),
    .Y(_07260_));
 sky130_fd_sc_hd__nand3_2 _29283_ (.A(_07254_),
    .B(_07251_),
    .C(_07252_),
    .Y(_07261_));
 sky130_fd_sc_hd__nand3_2 _29284_ (.A(_07258_),
    .B(_07260_),
    .C(_07261_),
    .Y(_07262_));
 sky130_fd_sc_hd__nand2_2 _29285_ (.A(_07257_),
    .B(_07262_),
    .Y(_07263_));
 sky130_fd_sc_hd__nand2_2 _29286_ (.A(\pcpi_mul.rs2[19] ),
    .B(_19639_),
    .Y(_07264_));
 sky130_fd_sc_hd__nand2_2 _29287_ (.A(\pcpi_mul.rs2[18] ),
    .B(_05104_),
    .Y(_07265_));
 sky130_fd_sc_hd__nor2_2 _29288_ (.A(_07264_),
    .B(_07265_),
    .Y(_07266_));
 sky130_fd_sc_hd__inv_2 _29289_ (.A(_07266_),
    .Y(_07267_));
 sky130_fd_sc_hd__nand2_2 _29290_ (.A(_07264_),
    .B(_07265_),
    .Y(_07268_));
 sky130_fd_sc_hd__nand2_2 _29291_ (.A(_07267_),
    .B(_07268_),
    .Y(_07269_));
 sky130_fd_sc_hd__nand2_2 _29292_ (.A(_07263_),
    .B(_07269_),
    .Y(_07270_));
 sky130_fd_sc_hd__nand3b_2 _29293_ (.A_N(_07269_),
    .B(_07257_),
    .C(_07262_),
    .Y(_07271_));
 sky130_fd_sc_hd__nand2_2 _29294_ (.A(_07270_),
    .B(_07271_),
    .Y(_07272_));
 sky130_fd_sc_hd__nand2_2 _29295_ (.A(_07272_),
    .B(_07055_),
    .Y(_07273_));
 sky130_fd_sc_hd__nand3_2 _29296_ (.A(_07056_),
    .B(_07270_),
    .C(_07271_),
    .Y(_07274_));
 sky130_fd_sc_hd__nand2_2 _29297_ (.A(_07273_),
    .B(_07274_),
    .Y(_07275_));
 sky130_fd_sc_hd__o21ai_2 _29298_ (.A1(_07199_),
    .A2(_07200_),
    .B1(_07275_),
    .Y(_07276_));
 sky130_fd_sc_hd__nand3_2 _29299_ (.A(_07191_),
    .B(_07196_),
    .C(_07198_),
    .Y(_07277_));
 sky130_fd_sc_hd__a21o_2 _29300_ (.A1(_07191_),
    .A2(_07197_),
    .B1(_07198_),
    .X(_07278_));
 sky130_fd_sc_hd__nand3b_2 _29301_ (.A_N(_07275_),
    .B(_07277_),
    .C(_07278_),
    .Y(_07279_));
 sky130_fd_sc_hd__nand3_2 _29302_ (.A(_07276_),
    .B(_07279_),
    .C(_07078_),
    .Y(_07280_));
 sky130_fd_sc_hd__o21bai_2 _29303_ (.A1(_07199_),
    .A2(_07200_),
    .B1_N(_07275_),
    .Y(_07281_));
 sky130_fd_sc_hd__nand3_2 _29304_ (.A(_07278_),
    .B(_07275_),
    .C(_07277_),
    .Y(_07282_));
 sky130_fd_sc_hd__nand3_2 _29305_ (.A(_07281_),
    .B(_07064_),
    .C(_07282_),
    .Y(_07283_));
 sky130_fd_sc_hd__nand2_2 _29306_ (.A(_07280_),
    .B(_07283_),
    .Y(_07284_));
 sky130_fd_sc_hd__a21boi_2 _29307_ (.A1(_06968_),
    .A2(_06973_),
    .B1_N(_06972_),
    .Y(_07285_));
 sky130_fd_sc_hd__a21oi_2 _29308_ (.A1(_06993_),
    .A2(_06989_),
    .B1(_07285_),
    .Y(_07286_));
 sky130_fd_sc_hd__and3_2 _29309_ (.A(_06992_),
    .B(_06989_),
    .C(_07285_),
    .X(_07287_));
 sky130_fd_sc_hd__nor2_2 _29310_ (.A(_07286_),
    .B(_07287_),
    .Y(_07288_));
 sky130_fd_sc_hd__nand2_2 _29311_ (.A(_07284_),
    .B(_07288_),
    .Y(_07289_));
 sky130_fd_sc_hd__a22oi_2 _29312_ (.A1(_07064_),
    .A2(_07072_),
    .B1(_07079_),
    .B2(_07085_),
    .Y(_07290_));
 sky130_fd_sc_hd__nand3b_2 _29313_ (.A_N(_07288_),
    .B(_07283_),
    .C(_07280_),
    .Y(_07291_));
 sky130_fd_sc_hd__nand3_2 _29314_ (.A(_07289_),
    .B(_07290_),
    .C(_07291_),
    .Y(_07292_));
 sky130_fd_sc_hd__o21ai_2 _29315_ (.A1(_07076_),
    .A2(_07065_),
    .B1(_07073_),
    .Y(_07293_));
 sky130_fd_sc_hd__o2bb2ai_2 _29316_ (.A1_N(_07283_),
    .A2_N(_07280_),
    .B1(_07286_),
    .B2(_07287_),
    .Y(_07294_));
 sky130_fd_sc_hd__nand3_2 _29317_ (.A(_07280_),
    .B(_07283_),
    .C(_07288_),
    .Y(_07295_));
 sky130_fd_sc_hd__nand3_2 _29318_ (.A(_07293_),
    .B(_07294_),
    .C(_07295_),
    .Y(_07296_));
 sky130_fd_sc_hd__nand2_2 _29319_ (.A(_07292_),
    .B(_07296_),
    .Y(_07297_));
 sky130_fd_sc_hd__a22oi_2 _29320_ (.A1(_07297_),
    .A2(_07074_),
    .B1(_07087_),
    .B2(_07082_),
    .Y(_07298_));
 sky130_fd_sc_hd__inv_2 _29321_ (.A(_07074_),
    .Y(_07299_));
 sky130_fd_sc_hd__nand3_2 _29322_ (.A(_07292_),
    .B(_07296_),
    .C(_07299_),
    .Y(_07300_));
 sky130_fd_sc_hd__o2bb2ai_2 _29323_ (.A1_N(_07296_),
    .A2_N(_07292_),
    .B1(_06880_),
    .B2(_06882_),
    .Y(_07301_));
 sky130_fd_sc_hd__nand2_2 _29324_ (.A(_07082_),
    .B(_07087_),
    .Y(_07302_));
 sky130_fd_sc_hd__a21oi_2 _29325_ (.A1(_07301_),
    .A2(_07300_),
    .B1(_07302_),
    .Y(_07303_));
 sky130_fd_sc_hd__a21oi_2 _29326_ (.A1(_07298_),
    .A2(_07300_),
    .B1(_07303_),
    .Y(_07304_));
 sky130_fd_sc_hd__nand3_2 _29327_ (.A(_07091_),
    .B(_07092_),
    .C(_07082_),
    .Y(_07305_));
 sky130_fd_sc_hd__nand2_2 _29328_ (.A(_07097_),
    .B(_07305_),
    .Y(_07306_));
 sky130_fd_sc_hd__xor2_2 _29329_ (.A(_07304_),
    .B(_07306_),
    .X(_02638_));
 sky130_fd_sc_hd__nand2_2 _29330_ (.A(_07277_),
    .B(_07273_),
    .Y(_07307_));
 sky130_fd_sc_hd__o22ai_2 _29331_ (.A1(_07055_),
    .A2(_07272_),
    .B1(_07199_),
    .B2(_07307_),
    .Y(_07308_));
 sky130_fd_sc_hd__inv_2 _29332_ (.A(_07117_),
    .Y(_07309_));
 sky130_fd_sc_hd__o21a_2 _29333_ (.A1(_06890_),
    .A2(_07118_),
    .B1(_07112_),
    .X(_07310_));
 sky130_fd_sc_hd__buf_1 _29334_ (.A(\pcpi_mul.rs1[13] ),
    .X(_07311_));
 sky130_fd_sc_hd__a22oi_2 _29335_ (.A1(_05542_),
    .A2(_06732_),
    .B1(_06508_),
    .B2(_07311_),
    .Y(_07312_));
 sky130_fd_sc_hd__inv_2 _29336_ (.A(_19599_),
    .Y(_07313_));
 sky130_fd_sc_hd__nand3_2 _29337_ (.A(_06008_),
    .B(_06010_),
    .C(_19602_),
    .Y(_07314_));
 sky130_fd_sc_hd__nor2_2 _29338_ (.A(_07313_),
    .B(_07314_),
    .Y(_07315_));
 sky130_fd_sc_hd__o22ai_2 _29339_ (.A1(_05244_),
    .A2(_06396_),
    .B1(_07312_),
    .B2(_07315_),
    .Y(_07316_));
 sky130_fd_sc_hd__o21ai_2 _29340_ (.A1(_07208_),
    .A2(_07204_),
    .B1(_07211_),
    .Y(_07317_));
 sky130_fd_sc_hd__and2_2 _29341_ (.A(_06496_),
    .B(_19596_),
    .X(_07318_));
 sky130_fd_sc_hd__a22o_2 _29342_ (.A1(_05448_),
    .A2(_07109_),
    .B1(_05445_),
    .B2(_06058_),
    .X(_07319_));
 sky130_fd_sc_hd__o211ai_2 _29343_ (.A1(_07313_),
    .A2(_07314_),
    .B1(_07318_),
    .C1(_07319_),
    .Y(_07320_));
 sky130_fd_sc_hd__nand3_2 _29344_ (.A(_07316_),
    .B(_07317_),
    .C(_07320_),
    .Y(_07321_));
 sky130_fd_sc_hd__o21ai_2 _29345_ (.A1(_07312_),
    .A2(_07315_),
    .B1(_07318_),
    .Y(_07322_));
 sky130_fd_sc_hd__o21ai_2 _29346_ (.A1(_07205_),
    .A2(_07206_),
    .B1(_07208_),
    .Y(_07323_));
 sky130_fd_sc_hd__nand2_2 _29347_ (.A(_07323_),
    .B(_07212_),
    .Y(_07324_));
 sky130_fd_sc_hd__o221ai_2 _29348_ (.A1(_05244_),
    .A2(_06396_),
    .B1(_07313_),
    .B2(_07314_),
    .C1(_07319_),
    .Y(_07325_));
 sky130_fd_sc_hd__nand3_2 _29349_ (.A(_07322_),
    .B(_07324_),
    .C(_07325_),
    .Y(_07326_));
 sky130_fd_sc_hd__nor2_2 _29350_ (.A(_07108_),
    .B(_07104_),
    .Y(_07327_));
 sky130_fd_sc_hd__o2bb2ai_2 _29351_ (.A1_N(_07321_),
    .A2_N(_07326_),
    .B1(_07102_),
    .B2(_07327_),
    .Y(_07328_));
 sky130_fd_sc_hd__nor2_2 _29352_ (.A(_07102_),
    .B(_07327_),
    .Y(_07329_));
 sky130_fd_sc_hd__nand3_2 _29353_ (.A(_07326_),
    .B(_07321_),
    .C(_07329_),
    .Y(_07330_));
 sky130_fd_sc_hd__nand2_2 _29354_ (.A(_07209_),
    .B(_07213_),
    .Y(_07331_));
 sky130_fd_sc_hd__a21oi_2 _29355_ (.A1(_07221_),
    .A2(_07222_),
    .B1(_07223_),
    .Y(_07332_));
 sky130_fd_sc_hd__nand2_2 _29356_ (.A(_07215_),
    .B(_07224_),
    .Y(_07333_));
 sky130_fd_sc_hd__o2bb2ai_2 _29357_ (.A1_N(_07229_),
    .A2_N(_07331_),
    .B1(_07332_),
    .B2(_07333_),
    .Y(_07334_));
 sky130_fd_sc_hd__a21oi_2 _29358_ (.A1(_07328_),
    .A2(_07330_),
    .B1(_07334_),
    .Y(_07335_));
 sky130_fd_sc_hd__nand2_2 _29359_ (.A(_07326_),
    .B(_07329_),
    .Y(_07336_));
 sky130_fd_sc_hd__inv_2 _29360_ (.A(_07321_),
    .Y(_07337_));
 sky130_fd_sc_hd__o211a_2 _29361_ (.A1(_07336_),
    .A2(_07337_),
    .B1(_07328_),
    .C1(_07334_),
    .X(_07338_));
 sky130_fd_sc_hd__o22ai_2 _29362_ (.A1(_07309_),
    .A2(_07310_),
    .B1(_07335_),
    .B2(_07338_),
    .Y(_07339_));
 sky130_fd_sc_hd__inv_2 _29363_ (.A(_07121_),
    .Y(_07340_));
 sky130_fd_sc_hd__nand2_2 _29364_ (.A(_07122_),
    .B(_07119_),
    .Y(_07341_));
 sky130_fd_sc_hd__and2_2 _29365_ (.A(_06916_),
    .B(_06900_),
    .X(_07342_));
 sky130_fd_sc_hd__o22ai_2 _29366_ (.A1(_07340_),
    .A2(_07341_),
    .B1(_07342_),
    .B2(_07123_),
    .Y(_07343_));
 sky130_fd_sc_hd__a21o_2 _29367_ (.A1(_07328_),
    .A2(_07330_),
    .B1(_07334_),
    .X(_07344_));
 sky130_fd_sc_hd__nand3_2 _29368_ (.A(_07334_),
    .B(_07328_),
    .C(_07330_),
    .Y(_07345_));
 sky130_fd_sc_hd__nand2_2 _29369_ (.A(_07121_),
    .B(_07112_),
    .Y(_07346_));
 sky130_fd_sc_hd__nand3_2 _29370_ (.A(_07344_),
    .B(_07345_),
    .C(_07346_),
    .Y(_07347_));
 sky130_fd_sc_hd__nand3_2 _29371_ (.A(_07339_),
    .B(_07343_),
    .C(_07347_),
    .Y(_07348_));
 sky130_fd_sc_hd__buf_1 _29372_ (.A(_07348_),
    .X(_07349_));
 sky130_fd_sc_hd__o21ai_2 _29373_ (.A1(_07335_),
    .A2(_07338_),
    .B1(_07346_),
    .Y(_07350_));
 sky130_fd_sc_hd__nand2_2 _29374_ (.A(_07127_),
    .B(_07342_),
    .Y(_07351_));
 sky130_fd_sc_hd__nand2_2 _29375_ (.A(_07351_),
    .B(_07126_),
    .Y(_07352_));
 sky130_fd_sc_hd__inv_2 _29376_ (.A(_07346_),
    .Y(_07353_));
 sky130_fd_sc_hd__nand3_2 _29377_ (.A(_07344_),
    .B(_07345_),
    .C(_07353_),
    .Y(_07354_));
 sky130_fd_sc_hd__nand3_2 _29378_ (.A(_07350_),
    .B(_07352_),
    .C(_07354_),
    .Y(_07355_));
 sky130_fd_sc_hd__a21boi_2 _29379_ (.A1(_07162_),
    .A2(_07151_),
    .B1_N(_07147_),
    .Y(_07356_));
 sky130_fd_sc_hd__a21oi_2 _29380_ (.A1(_07140_),
    .A2(_07137_),
    .B1(_07145_),
    .Y(_07357_));
 sky130_fd_sc_hd__buf_1 _29381_ (.A(\pcpi_mul.rs1[20] ),
    .X(_07358_));
 sky130_fd_sc_hd__nand2_2 _29382_ (.A(_05192_),
    .B(_07358_),
    .Y(_07359_));
 sky130_fd_sc_hd__buf_1 _29383_ (.A(\pcpi_mul.rs1[16] ),
    .X(_07360_));
 sky130_fd_sc_hd__a22oi_2 _29384_ (.A1(_05321_),
    .A2(_19593_),
    .B1(_05322_),
    .B2(_07360_),
    .Y(_07361_));
 sky130_fd_sc_hd__nor2_2 _29385_ (.A(_07359_),
    .B(_07361_),
    .Y(_07362_));
 sky130_fd_sc_hd__nand2_2 _29386_ (.A(_06731_),
    .B(_06373_),
    .Y(_07363_));
 sky130_fd_sc_hd__nand2_2 _29387_ (.A(_05891_),
    .B(_06542_),
    .Y(_07364_));
 sky130_fd_sc_hd__or2_2 _29388_ (.A(_07363_),
    .B(_07364_),
    .X(_07365_));
 sky130_fd_sc_hd__nand2_2 _29389_ (.A(_07362_),
    .B(_07365_),
    .Y(_07366_));
 sky130_fd_sc_hd__nor2_2 _29390_ (.A(_07363_),
    .B(_07364_),
    .Y(_07367_));
 sky130_fd_sc_hd__o21ai_2 _29391_ (.A1(_07361_),
    .A2(_07367_),
    .B1(_07359_),
    .Y(_07368_));
 sky130_fd_sc_hd__nand3b_2 _29392_ (.A_N(_07357_),
    .B(_07366_),
    .C(_07368_),
    .Y(_07369_));
 sky130_fd_sc_hd__inv_2 _29393_ (.A(_07361_),
    .Y(_07370_));
 sky130_fd_sc_hd__nand3_2 _29394_ (.A(_07365_),
    .B(_07370_),
    .C(_07359_),
    .Y(_07371_));
 sky130_fd_sc_hd__o21bai_2 _29395_ (.A1(_07361_),
    .A2(_07367_),
    .B1_N(_07359_),
    .Y(_07372_));
 sky130_fd_sc_hd__nand3_2 _29396_ (.A(_07371_),
    .B(_07357_),
    .C(_07372_),
    .Y(_07373_));
 sky130_fd_sc_hd__nand2_2 _29397_ (.A(_07369_),
    .B(_07373_),
    .Y(_07374_));
 sky130_fd_sc_hd__nand2_2 _29398_ (.A(_05209_),
    .B(_07156_),
    .Y(_07375_));
 sky130_fd_sc_hd__a21o_2 _29399_ (.A1(_05143_),
    .A2(_19582_),
    .B1(_07375_),
    .X(_07376_));
 sky130_fd_sc_hd__buf_1 _29400_ (.A(\pcpi_mul.rs1[19] ),
    .X(_07377_));
 sky130_fd_sc_hd__nand2_2 _29401_ (.A(_05210_),
    .B(_07377_),
    .Y(_07378_));
 sky130_fd_sc_hd__a21o_2 _29402_ (.A1(_05203_),
    .A2(_19585_),
    .B1(_07378_),
    .X(_07379_));
 sky130_fd_sc_hd__buf_1 _29403_ (.A(_06951_),
    .X(_07380_));
 sky130_fd_sc_hd__nand2_2 _29404_ (.A(_19393_),
    .B(_07380_),
    .Y(_07381_));
 sky130_fd_sc_hd__a21oi_2 _29405_ (.A1(_07376_),
    .A2(_07379_),
    .B1(_07381_),
    .Y(_07382_));
 sky130_fd_sc_hd__and3_2 _29406_ (.A(_07376_),
    .B(_07379_),
    .C(_07381_),
    .X(_07383_));
 sky130_fd_sc_hd__nor2_2 _29407_ (.A(_07382_),
    .B(_07383_),
    .Y(_07384_));
 sky130_fd_sc_hd__nand2_2 _29408_ (.A(_07374_),
    .B(_07384_),
    .Y(_07385_));
 sky130_fd_sc_hd__o211ai_2 _29409_ (.A1(_07382_),
    .A2(_07383_),
    .B1(_07373_),
    .C1(_07369_),
    .Y(_07386_));
 sky130_fd_sc_hd__nand3_2 _29410_ (.A(_07356_),
    .B(_07385_),
    .C(_07386_),
    .Y(_07387_));
 sky130_fd_sc_hd__o21ai_2 _29411_ (.A1(_07166_),
    .A2(_07173_),
    .B1(_07147_),
    .Y(_07388_));
 sky130_fd_sc_hd__o2bb2ai_2 _29412_ (.A1_N(_07373_),
    .A2_N(_07369_),
    .B1(_07383_),
    .B2(_07382_),
    .Y(_07389_));
 sky130_fd_sc_hd__nand3_2 _29413_ (.A(_07384_),
    .B(_07373_),
    .C(_07369_),
    .Y(_07390_));
 sky130_fd_sc_hd__nand3_2 _29414_ (.A(_07388_),
    .B(_07389_),
    .C(_07390_),
    .Y(_07391_));
 sky130_fd_sc_hd__nor2_2 _29415_ (.A(_07154_),
    .B(_07157_),
    .Y(_07392_));
 sky130_fd_sc_hd__nor2_2 _29416_ (.A(_07392_),
    .B(_07160_),
    .Y(_07393_));
 sky130_fd_sc_hd__inv_2 _29417_ (.A(_07393_),
    .Y(_07394_));
 sky130_fd_sc_hd__and3_2 _29418_ (.A(_07387_),
    .B(_07391_),
    .C(_07394_),
    .X(_07395_));
 sky130_fd_sc_hd__a21oi_2 _29419_ (.A1(_07387_),
    .A2(_07391_),
    .B1(_07394_),
    .Y(_07396_));
 sky130_fd_sc_hd__o2bb2ai_2 _29420_ (.A1_N(_07349_),
    .A2_N(_07355_),
    .B1(_07395_),
    .B2(_07396_),
    .Y(_07397_));
 sky130_fd_sc_hd__inv_2 _29421_ (.A(_07262_),
    .Y(_07398_));
 sky130_fd_sc_hd__a31oi_2 _29422_ (.A1(_07356_),
    .A2(_07385_),
    .A3(_07386_),
    .B1(_07393_),
    .Y(_07399_));
 sky130_fd_sc_hd__a21oi_2 _29423_ (.A1(_07391_),
    .A2(_07399_),
    .B1(_07396_),
    .Y(_07400_));
 sky130_fd_sc_hd__nand3_2 _29424_ (.A(_07400_),
    .B(_07355_),
    .C(_07349_),
    .Y(_07401_));
 sky130_fd_sc_hd__nand3_2 _29425_ (.A(_07397_),
    .B(_07398_),
    .C(_07401_),
    .Y(_07402_));
 sky130_fd_sc_hd__buf_1 _29426_ (.A(_07402_),
    .X(_07403_));
 sky130_fd_sc_hd__nand2_2 _29427_ (.A(_07355_),
    .B(_07348_),
    .Y(_07404_));
 sky130_fd_sc_hd__nand2_2 _29428_ (.A(_07404_),
    .B(_07400_),
    .Y(_07405_));
 sky130_fd_sc_hd__o211ai_2 _29429_ (.A1(_07396_),
    .A2(_07395_),
    .B1(_07349_),
    .C1(_07355_),
    .Y(_07406_));
 sky130_fd_sc_hd__nand3_2 _29430_ (.A(_07405_),
    .B(_07262_),
    .C(_07406_),
    .Y(_07407_));
 sky130_fd_sc_hd__nor2_2 _29431_ (.A(_07179_),
    .B(_07132_),
    .Y(_07408_));
 sky130_fd_sc_hd__o2bb2ai_2 _29432_ (.A1_N(_07403_),
    .A2_N(_07407_),
    .B1(_07130_),
    .B2(_07408_),
    .Y(_07409_));
 sky130_fd_sc_hd__o21ai_2 _29433_ (.A1(_07130_),
    .A2(_07188_),
    .B1(_07189_),
    .Y(_07410_));
 sky130_fd_sc_hd__nand3_2 _29434_ (.A(_07407_),
    .B(_07402_),
    .C(_07410_),
    .Y(_07411_));
 sky130_fd_sc_hd__nand2_2 _29435_ (.A(_07409_),
    .B(_07411_),
    .Y(_07412_));
 sky130_fd_sc_hd__nand2_2 _29436_ (.A(_07241_),
    .B(_07244_),
    .Y(_07413_));
 sky130_fd_sc_hd__nand3_2 _29437_ (.A(\pcpi_mul.rs2[17] ),
    .B(_19356_),
    .C(_19629_),
    .Y(_07414_));
 sky130_fd_sc_hd__nor2_2 _29438_ (.A(_05849_),
    .B(_07414_),
    .Y(_07415_));
 sky130_fd_sc_hd__buf_1 _29439_ (.A(\pcpi_mul.rs2[17] ),
    .X(_07416_));
 sky130_fd_sc_hd__buf_1 _29440_ (.A(_19356_),
    .X(_07417_));
 sky130_fd_sc_hd__a22o_2 _29441_ (.A1(_07416_),
    .A2(_05271_),
    .B1(_07417_),
    .B2(_05158_),
    .X(_07418_));
 sky130_fd_sc_hd__nand2_2 _29442_ (.A(\pcpi_mul.rs2[15] ),
    .B(_19624_),
    .Y(_07419_));
 sky130_fd_sc_hd__inv_2 _29443_ (.A(_07419_),
    .Y(_07420_));
 sky130_fd_sc_hd__nand2_2 _29444_ (.A(_07418_),
    .B(_07420_),
    .Y(_07421_));
 sky130_fd_sc_hd__a22oi_2 _29445_ (.A1(_07416_),
    .A2(_05271_),
    .B1(_07417_),
    .B2(_05206_),
    .Y(_07422_));
 sky130_fd_sc_hd__o21ai_2 _29446_ (.A1(_07422_),
    .A2(_07415_),
    .B1(_07419_),
    .Y(_07423_));
 sky130_fd_sc_hd__o211ai_2 _29447_ (.A1(_07415_),
    .A2(_07421_),
    .B1(_07266_),
    .C1(_07423_),
    .Y(_07424_));
 sky130_fd_sc_hd__o21ai_2 _29448_ (.A1(_07422_),
    .A2(_07415_),
    .B1(_07420_),
    .Y(_07425_));
 sky130_fd_sc_hd__o211ai_2 _29449_ (.A1(_06105_),
    .A2(_07414_),
    .B1(_07419_),
    .C1(_07418_),
    .Y(_07426_));
 sky130_fd_sc_hd__nand3_2 _29450_ (.A(_07425_),
    .B(_07267_),
    .C(_07426_),
    .Y(_07427_));
 sky130_fd_sc_hd__a21o_2 _29451_ (.A1(_07239_),
    .A2(_07237_),
    .B1(_07235_),
    .X(_07428_));
 sky130_fd_sc_hd__a21oi_2 _29452_ (.A1(_07424_),
    .A2(_07427_),
    .B1(_07428_),
    .Y(_07429_));
 sky130_fd_sc_hd__and3_2 _29453_ (.A(_07424_),
    .B(_07427_),
    .C(_07428_),
    .X(_07430_));
 sky130_fd_sc_hd__o22ai_2 _29454_ (.A1(_07247_),
    .A2(_07413_),
    .B1(_07429_),
    .B2(_07430_),
    .Y(_07431_));
 sky130_fd_sc_hd__a21o_2 _29455_ (.A1(_07424_),
    .A2(_07427_),
    .B1(_07428_),
    .X(_07432_));
 sky130_fd_sc_hd__and3_2 _29456_ (.A(_07241_),
    .B(_07242_),
    .C(_07244_),
    .X(_07433_));
 sky130_fd_sc_hd__nand3_2 _29457_ (.A(_07424_),
    .B(_07427_),
    .C(_07428_),
    .Y(_07434_));
 sky130_fd_sc_hd__nand3_2 _29458_ (.A(_07432_),
    .B(_07433_),
    .C(_07434_),
    .Y(_07435_));
 sky130_fd_sc_hd__and4_2 _29459_ (.A(_05800_),
    .B(_06432_),
    .C(_05598_),
    .D(_05614_),
    .X(_07436_));
 sky130_fd_sc_hd__a22o_2 _29460_ (.A1(_05956_),
    .A2(_06327_),
    .B1(_07034_),
    .B2(_06889_),
    .X(_07437_));
 sky130_fd_sc_hd__nand2_2 _29461_ (.A(_05672_),
    .B(_19605_),
    .Y(_07438_));
 sky130_fd_sc_hd__inv_2 _29462_ (.A(_07438_),
    .Y(_07439_));
 sky130_fd_sc_hd__nand2_2 _29463_ (.A(_07437_),
    .B(_07439_),
    .Y(_07440_));
 sky130_fd_sc_hd__a22oi_2 _29464_ (.A1(_07203_),
    .A2(_06492_),
    .B1(_19373_),
    .B2(_06889_),
    .Y(_07441_));
 sky130_fd_sc_hd__o21ai_2 _29465_ (.A1(_07441_),
    .A2(_07436_),
    .B1(_07438_),
    .Y(_07442_));
 sky130_fd_sc_hd__o21ai_2 _29466_ (.A1(_07436_),
    .A2(_07440_),
    .B1(_07442_),
    .Y(_07443_));
 sky130_fd_sc_hd__a22oi_2 _29467_ (.A1(_06441_),
    .A2(_19622_),
    .B1(_06443_),
    .B2(_05426_),
    .Y(_07444_));
 sky130_fd_sc_hd__nand2_2 _29468_ (.A(_06269_),
    .B(_19621_),
    .Y(_07445_));
 sky130_fd_sc_hd__nand2_2 _29469_ (.A(\pcpi_mul.rs2[13] ),
    .B(_05419_),
    .Y(_07446_));
 sky130_fd_sc_hd__nor2_2 _29470_ (.A(_07445_),
    .B(_07446_),
    .Y(_07447_));
 sky130_fd_sc_hd__nand2_2 _29471_ (.A(_06117_),
    .B(_05730_),
    .Y(_07448_));
 sky130_fd_sc_hd__o21ai_2 _29472_ (.A1(_07444_),
    .A2(_07447_),
    .B1(_07448_),
    .Y(_07449_));
 sky130_fd_sc_hd__buf_1 _29473_ (.A(_06275_),
    .X(_07450_));
 sky130_fd_sc_hd__nand3b_2 _29474_ (.A_N(_07445_),
    .B(_07450_),
    .C(_19619_),
    .Y(_07451_));
 sky130_fd_sc_hd__inv_2 _29475_ (.A(_07448_),
    .Y(_07452_));
 sky130_fd_sc_hd__nand2_2 _29476_ (.A(_07445_),
    .B(_07446_),
    .Y(_07453_));
 sky130_fd_sc_hd__nand3_2 _29477_ (.A(_07451_),
    .B(_07452_),
    .C(_07453_),
    .Y(_07454_));
 sky130_fd_sc_hd__o21ai_2 _29478_ (.A1(_07218_),
    .A2(_07216_),
    .B1(_07221_),
    .Y(_07455_));
 sky130_fd_sc_hd__a21oi_2 _29479_ (.A1(_07449_),
    .A2(_07454_),
    .B1(_07455_),
    .Y(_07456_));
 sky130_fd_sc_hd__nor2_2 _29480_ (.A(_07443_),
    .B(_07456_),
    .Y(_07457_));
 sky130_fd_sc_hd__nand3_2 _29481_ (.A(_07449_),
    .B(_07454_),
    .C(_07455_),
    .Y(_07458_));
 sky130_fd_sc_hd__o21ai_2 _29482_ (.A1(_07444_),
    .A2(_07447_),
    .B1(_07452_),
    .Y(_07459_));
 sky130_fd_sc_hd__nand3_2 _29483_ (.A(_07451_),
    .B(_07448_),
    .C(_07453_),
    .Y(_07460_));
 sky130_fd_sc_hd__nand3b_2 _29484_ (.A_N(_07455_),
    .B(_07459_),
    .C(_07460_),
    .Y(_07461_));
 sky130_fd_sc_hd__a21boi_2 _29485_ (.A1(_07461_),
    .A2(_07458_),
    .B1_N(_07443_),
    .Y(_07462_));
 sky130_fd_sc_hd__a21oi_2 _29486_ (.A1(_07457_),
    .A2(_07458_),
    .B1(_07462_),
    .Y(_07463_));
 sky130_fd_sc_hd__a21oi_2 _29487_ (.A1(_07431_),
    .A2(_07435_),
    .B1(_07463_),
    .Y(_07464_));
 sky130_fd_sc_hd__nand2_2 _29488_ (.A(_07433_),
    .B(_07434_),
    .Y(_07465_));
 sky130_fd_sc_hd__o211a_2 _29489_ (.A1(_07429_),
    .A2(_07465_),
    .B1(_07463_),
    .C1(_07431_),
    .X(_07466_));
 sky130_fd_sc_hd__nor2_2 _29490_ (.A(_07006_),
    .B(_07250_),
    .Y(_07467_));
 sky130_fd_sc_hd__a21oi_2 _29491_ (.A1(_07254_),
    .A2(_07251_),
    .B1(_07467_),
    .Y(_07468_));
 sky130_fd_sc_hd__o21ai_2 _29492_ (.A1(_07464_),
    .A2(_07466_),
    .B1(_07468_),
    .Y(_07469_));
 sky130_fd_sc_hd__nor2_2 _29493_ (.A(_07429_),
    .B(_07465_),
    .Y(_07470_));
 sky130_fd_sc_hd__nand2_2 _29494_ (.A(_07431_),
    .B(_07463_),
    .Y(_07471_));
 sky130_fd_sc_hd__a31o_2 _29495_ (.A1(_07231_),
    .A2(_07251_),
    .A3(_07232_),
    .B1(_07467_),
    .X(_07472_));
 sky130_fd_sc_hd__a21o_2 _29496_ (.A1(_07431_),
    .A2(_07435_),
    .B1(_07463_),
    .X(_07473_));
 sky130_fd_sc_hd__o211ai_2 _29497_ (.A1(_07470_),
    .A2(_07471_),
    .B1(_07472_),
    .C1(_07473_),
    .Y(_07474_));
 sky130_fd_sc_hd__buf_1 _29498_ (.A(\pcpi_mul.rs2[18] ),
    .X(_07475_));
 sky130_fd_sc_hd__nand2_2 _29499_ (.A(_07475_),
    .B(_05119_),
    .Y(_07476_));
 sky130_fd_sc_hd__inv_2 _29500_ (.A(_07476_),
    .Y(_07477_));
 sky130_fd_sc_hd__buf_1 _29501_ (.A(\pcpi_mul.rs2[19] ),
    .X(_07478_));
 sky130_fd_sc_hd__nand2_2 _29502_ (.A(_07478_),
    .B(_05190_),
    .Y(_07479_));
 sky130_fd_sc_hd__buf_1 _29503_ (.A(\pcpi_mul.rs2[20] ),
    .X(_07480_));
 sky130_fd_sc_hd__buf_1 _29504_ (.A(_07480_),
    .X(_07481_));
 sky130_fd_sc_hd__nand3b_2 _29505_ (.A_N(_07479_),
    .B(_07481_),
    .C(_06598_),
    .Y(_07482_));
 sky130_fd_sc_hd__buf_1 _29506_ (.A(_19346_),
    .X(_07483_));
 sky130_fd_sc_hd__nand2_2 _29507_ (.A(_07483_),
    .B(_05188_),
    .Y(_07484_));
 sky130_fd_sc_hd__nand2_2 _29508_ (.A(_07479_),
    .B(_07484_),
    .Y(_07485_));
 sky130_fd_sc_hd__nand2_2 _29509_ (.A(_07482_),
    .B(_07485_),
    .Y(_07486_));
 sky130_fd_sc_hd__nor2_2 _29510_ (.A(_07477_),
    .B(_07486_),
    .Y(_07487_));
 sky130_fd_sc_hd__and2_2 _29511_ (.A(_07486_),
    .B(_07477_),
    .X(_07488_));
 sky130_fd_sc_hd__nor2_2 _29512_ (.A(_07487_),
    .B(_07488_),
    .Y(_07489_));
 sky130_fd_sc_hd__inv_2 _29513_ (.A(_07489_),
    .Y(_07490_));
 sky130_fd_sc_hd__a21oi_2 _29514_ (.A1(_07469_),
    .A2(_07474_),
    .B1(_07490_),
    .Y(_07491_));
 sky130_fd_sc_hd__and3_2 _29515_ (.A(_07469_),
    .B(_07474_),
    .C(_07490_),
    .X(_07492_));
 sky130_fd_sc_hd__buf_1 _29516_ (.A(_07492_),
    .X(_07493_));
 sky130_fd_sc_hd__o22ai_2 _29517_ (.A1(_07263_),
    .A2(_07269_),
    .B1(_07491_),
    .B2(_07493_),
    .Y(_07494_));
 sky130_fd_sc_hd__inv_2 _29518_ (.A(_07271_),
    .Y(_07495_));
 sky130_fd_sc_hd__nand2_2 _29519_ (.A(_07469_),
    .B(_07474_),
    .Y(_07496_));
 sky130_fd_sc_hd__nand2_2 _29520_ (.A(_07496_),
    .B(_07489_),
    .Y(_07497_));
 sky130_fd_sc_hd__nand3_2 _29521_ (.A(_07469_),
    .B(_07474_),
    .C(_07490_),
    .Y(_07498_));
 sky130_fd_sc_hd__nand3_2 _29522_ (.A(_07495_),
    .B(_07497_),
    .C(_07498_),
    .Y(_07499_));
 sky130_fd_sc_hd__nand2_2 _29523_ (.A(_07494_),
    .B(_07499_),
    .Y(_07500_));
 sky130_fd_sc_hd__nand2_2 _29524_ (.A(_07412_),
    .B(_07500_),
    .Y(_07501_));
 sky130_fd_sc_hd__nand2_2 _29525_ (.A(_07495_),
    .B(_07497_),
    .Y(_07502_));
 sky130_fd_sc_hd__buf_1 _29526_ (.A(_07411_),
    .X(_07503_));
 sky130_fd_sc_hd__o2111ai_2 _29527_ (.A1(_07493_),
    .A2(_07502_),
    .B1(_07494_),
    .C1(_07503_),
    .D1(_07409_),
    .Y(_07504_));
 sky130_fd_sc_hd__nand3_2 _29528_ (.A(_07308_),
    .B(_07501_),
    .C(_07504_),
    .Y(_07505_));
 sky130_fd_sc_hd__a22oi_2 _29529_ (.A1(_07494_),
    .A2(_07499_),
    .B1(_07409_),
    .B2(_07503_),
    .Y(_07506_));
 sky130_fd_sc_hd__a21oi_2 _29530_ (.A1(_07407_),
    .A2(_07403_),
    .B1(_07410_),
    .Y(_07507_));
 sky130_fd_sc_hd__nand3_2 _29531_ (.A(_07494_),
    .B(_07411_),
    .C(_07499_),
    .Y(_07508_));
 sky130_fd_sc_hd__nor2_2 _29532_ (.A(_07507_),
    .B(_07508_),
    .Y(_07509_));
 sky130_fd_sc_hd__a21oi_2 _29533_ (.A1(_07270_),
    .A2(_07271_),
    .B1(_07056_),
    .Y(_07510_));
 sky130_fd_sc_hd__a31oi_2 _29534_ (.A1(_07191_),
    .A2(_07197_),
    .A3(_07198_),
    .B1(_07510_),
    .Y(_07511_));
 sky130_fd_sc_hd__a21boi_2 _29535_ (.A1(_07511_),
    .A2(_07278_),
    .B1_N(_07274_),
    .Y(_07512_));
 sky130_fd_sc_hd__o21ai_2 _29536_ (.A1(_07506_),
    .A2(_07509_),
    .B1(_07512_),
    .Y(_07513_));
 sky130_fd_sc_hd__nor2_2 _29537_ (.A(_07185_),
    .B(_07172_),
    .Y(_07514_));
 sky130_fd_sc_hd__a21oi_2 _29538_ (.A1(_07277_),
    .A2(_07197_),
    .B1(_07514_),
    .Y(_07515_));
 sky130_fd_sc_hd__buf_1 _29539_ (.A(_07515_),
    .X(_07516_));
 sky130_fd_sc_hd__and3_2 _29540_ (.A(_07277_),
    .B(_07197_),
    .C(_07514_),
    .X(_07517_));
 sky130_fd_sc_hd__o2bb2ai_2 _29541_ (.A1_N(_07505_),
    .A2_N(_07513_),
    .B1(_07516_),
    .B2(_07517_),
    .Y(_07518_));
 sky130_fd_sc_hd__nor2_2 _29542_ (.A(_07515_),
    .B(_07517_),
    .Y(_07519_));
 sky130_fd_sc_hd__nand3_2 _29543_ (.A(_07513_),
    .B(_07505_),
    .C(_07519_),
    .Y(_07520_));
 sky130_fd_sc_hd__nand2_2 _29544_ (.A(_07283_),
    .B(_07288_),
    .Y(_07521_));
 sky130_fd_sc_hd__nand2_2 _29545_ (.A(_07521_),
    .B(_07280_),
    .Y(_07522_));
 sky130_fd_sc_hd__a21oi_2 _29546_ (.A1(_07518_),
    .A2(_07520_),
    .B1(_07522_),
    .Y(_07523_));
 sky130_fd_sc_hd__nand2_2 _29547_ (.A(_07513_),
    .B(_07519_),
    .Y(_07524_));
 sky130_fd_sc_hd__inv_2 _29548_ (.A(_07505_),
    .Y(_07525_));
 sky130_fd_sc_hd__o211a_2 _29549_ (.A1(_07524_),
    .A2(_07525_),
    .B1(_07518_),
    .C1(_07522_),
    .X(_07526_));
 sky130_fd_sc_hd__o21ai_2 _29550_ (.A1(_07523_),
    .A2(_07526_),
    .B1(_07286_),
    .Y(_07527_));
 sky130_fd_sc_hd__a21boi_2 _29551_ (.A1(_07292_),
    .A2(_07299_),
    .B1_N(_07296_),
    .Y(_07528_));
 sky130_fd_sc_hd__nand2_2 _29552_ (.A(_07518_),
    .B(_07520_),
    .Y(_07529_));
 sky130_fd_sc_hd__a21boi_2 _29553_ (.A1(_07288_),
    .A2(_07283_),
    .B1_N(_07280_),
    .Y(_07530_));
 sky130_fd_sc_hd__nand2_2 _29554_ (.A(_07529_),
    .B(_07530_),
    .Y(_07531_));
 sky130_fd_sc_hd__inv_2 _29555_ (.A(_07286_),
    .Y(_07532_));
 sky130_fd_sc_hd__nand3_2 _29556_ (.A(_07522_),
    .B(_07518_),
    .C(_07520_),
    .Y(_07533_));
 sky130_fd_sc_hd__nand3_2 _29557_ (.A(_07531_),
    .B(_07532_),
    .C(_07533_),
    .Y(_07534_));
 sky130_fd_sc_hd__nand3_2 _29558_ (.A(_07527_),
    .B(_07528_),
    .C(_07534_),
    .Y(_07535_));
 sky130_fd_sc_hd__o21ai_2 _29559_ (.A1(_07523_),
    .A2(_07526_),
    .B1(_07532_),
    .Y(_07536_));
 sky130_fd_sc_hd__nand2_2 _29560_ (.A(_07292_),
    .B(_07299_),
    .Y(_07537_));
 sky130_fd_sc_hd__nand2_2 _29561_ (.A(_07537_),
    .B(_07296_),
    .Y(_07538_));
 sky130_fd_sc_hd__nand3_2 _29562_ (.A(_07531_),
    .B(_07286_),
    .C(_07533_),
    .Y(_07539_));
 sky130_fd_sc_hd__nand3_2 _29563_ (.A(_07536_),
    .B(_07538_),
    .C(_07539_),
    .Y(_07540_));
 sky130_fd_sc_hd__and2_2 _29564_ (.A(_07535_),
    .B(_07540_),
    .X(_07541_));
 sky130_fd_sc_hd__nand3_2 _29565_ (.A(_06876_),
    .B(_06675_),
    .C(_06677_),
    .Y(_07542_));
 sky130_fd_sc_hd__nor2_2 _29566_ (.A(_06875_),
    .B(_07542_),
    .Y(_07543_));
 sky130_fd_sc_hd__nand3_2 _29567_ (.A(_07543_),
    .B(_07094_),
    .C(_07304_),
    .Y(_07544_));
 sky130_fd_sc_hd__a21oi_2 _29568_ (.A1(_06677_),
    .A2(_06876_),
    .B1(_06875_),
    .Y(_07545_));
 sky130_fd_sc_hd__o2bb2ai_2 _29569_ (.A1_N(_07300_),
    .A2_N(_07298_),
    .B1(_07305_),
    .B2(_07303_),
    .Y(_07546_));
 sky130_fd_sc_hd__a31oi_2 _29570_ (.A1(_07094_),
    .A2(_07304_),
    .A3(_07545_),
    .B1(_07546_),
    .Y(_07547_));
 sky130_fd_sc_hd__o21a_2 _29571_ (.A1(_07544_),
    .A2(_06491_),
    .B1(_07547_),
    .X(_07548_));
 sky130_fd_sc_hd__xnor2_2 _29572_ (.A(_07541_),
    .B(_07548_),
    .Y(_02639_));
 sky130_fd_sc_hd__nand2_2 _29573_ (.A(_07524_),
    .B(_07505_),
    .Y(_07549_));
 sky130_fd_sc_hd__o21ai_2 _29574_ (.A1(_07507_),
    .A2(_07508_),
    .B1(_07499_),
    .Y(_07550_));
 sky130_fd_sc_hd__o21ai_2 _29575_ (.A1(_07443_),
    .A2(_07456_),
    .B1(_07458_),
    .Y(_07551_));
 sky130_fd_sc_hd__a22oi_2 _29576_ (.A1(_05758_),
    .A2(_06058_),
    .B1(_05760_),
    .B2(_06387_),
    .Y(_07552_));
 sky130_fd_sc_hd__nand3_2 _29577_ (.A(_19379_),
    .B(_06334_),
    .C(_19599_),
    .Y(_07553_));
 sky130_fd_sc_hd__nor2_2 _29578_ (.A(_06395_),
    .B(_07553_),
    .Y(_07554_));
 sky130_fd_sc_hd__nand2_2 _29579_ (.A(_05763_),
    .B(_06372_),
    .Y(_07555_));
 sky130_fd_sc_hd__inv_2 _29580_ (.A(_07555_),
    .Y(_07556_));
 sky130_fd_sc_hd__o21ai_2 _29581_ (.A1(_07552_),
    .A2(_07554_),
    .B1(_07556_),
    .Y(_07557_));
 sky130_fd_sc_hd__a21oi_2 _29582_ (.A1(_07437_),
    .A2(_07439_),
    .B1(_07436_),
    .Y(_07558_));
 sky130_fd_sc_hd__a22o_2 _29583_ (.A1(_05448_),
    .A2(_06058_),
    .B1(_05445_),
    .B2(_06387_),
    .X(_07559_));
 sky130_fd_sc_hd__o211ai_2 _29584_ (.A1(_06396_),
    .A2(_07553_),
    .B1(_07555_),
    .C1(_07559_),
    .Y(_07560_));
 sky130_fd_sc_hd__nand3_2 _29585_ (.A(_07557_),
    .B(_07558_),
    .C(_07560_),
    .Y(_07561_));
 sky130_fd_sc_hd__o21ai_2 _29586_ (.A1(_07552_),
    .A2(_07554_),
    .B1(_07555_),
    .Y(_07562_));
 sky130_fd_sc_hd__nand2_2 _29587_ (.A(_05800_),
    .B(_05614_),
    .Y(_07563_));
 sky130_fd_sc_hd__nand3b_2 _29588_ (.A_N(_07563_),
    .B(_05803_),
    .C(_05738_),
    .Y(_07564_));
 sky130_fd_sc_hd__o21ai_2 _29589_ (.A1(_07438_),
    .A2(_07441_),
    .B1(_07564_),
    .Y(_07565_));
 sky130_fd_sc_hd__o211ai_2 _29590_ (.A1(_06396_),
    .A2(_07553_),
    .B1(_07556_),
    .C1(_07559_),
    .Y(_07566_));
 sky130_fd_sc_hd__nand3_2 _29591_ (.A(_07562_),
    .B(_07565_),
    .C(_07566_),
    .Y(_07567_));
 sky130_fd_sc_hd__a21o_2 _29592_ (.A1(_07319_),
    .A2(_07318_),
    .B1(_07315_),
    .X(_07568_));
 sky130_fd_sc_hd__a21o_2 _29593_ (.A1(_07561_),
    .A2(_07567_),
    .B1(_07568_),
    .X(_07569_));
 sky130_fd_sc_hd__nand3_2 _29594_ (.A(_07561_),
    .B(_07567_),
    .C(_07568_),
    .Y(_07570_));
 sky130_fd_sc_hd__nand3_2 _29595_ (.A(_07551_),
    .B(_07569_),
    .C(_07570_),
    .Y(_07571_));
 sky130_fd_sc_hd__and2_2 _29596_ (.A(_07458_),
    .B(_07443_),
    .X(_07572_));
 sky130_fd_sc_hd__a21oi_2 _29597_ (.A1(_07561_),
    .A2(_07567_),
    .B1(_07568_),
    .Y(_07573_));
 sky130_fd_sc_hd__and3_2 _29598_ (.A(_07561_),
    .B(_07567_),
    .C(_07568_),
    .X(_07574_));
 sky130_fd_sc_hd__o22ai_2 _29599_ (.A1(_07456_),
    .A2(_07572_),
    .B1(_07573_),
    .B2(_07574_),
    .Y(_07575_));
 sky130_fd_sc_hd__and2_2 _29600_ (.A(_07326_),
    .B(_07329_),
    .X(_07576_));
 sky130_fd_sc_hd__o2bb2ai_2 _29601_ (.A1_N(_07571_),
    .A2_N(_07575_),
    .B1(_07337_),
    .B2(_07576_),
    .Y(_07577_));
 sky130_fd_sc_hd__a21oi_2 _29602_ (.A1(_07344_),
    .A2(_07346_),
    .B1(_07338_),
    .Y(_07578_));
 sky130_fd_sc_hd__and2_2 _29603_ (.A(_07336_),
    .B(_07321_),
    .X(_07579_));
 sky130_fd_sc_hd__nand3_2 _29604_ (.A(_07575_),
    .B(_07571_),
    .C(_07579_),
    .Y(_07580_));
 sky130_fd_sc_hd__nand3_2 _29605_ (.A(_07577_),
    .B(_07578_),
    .C(_07580_),
    .Y(_07581_));
 sky130_fd_sc_hd__inv_2 _29606_ (.A(_07326_),
    .Y(_07582_));
 sky130_fd_sc_hd__nor2_2 _29607_ (.A(_07329_),
    .B(_07337_),
    .Y(_07583_));
 sky130_fd_sc_hd__o2bb2ai_2 _29608_ (.A1_N(_07571_),
    .A2_N(_07575_),
    .B1(_07582_),
    .B2(_07583_),
    .Y(_07584_));
 sky130_fd_sc_hd__o21ai_2 _29609_ (.A1(_07335_),
    .A2(_07353_),
    .B1(_07345_),
    .Y(_07585_));
 sky130_fd_sc_hd__nand3b_2 _29610_ (.A_N(_07579_),
    .B(_07575_),
    .C(_07571_),
    .Y(_07586_));
 sky130_fd_sc_hd__nand3_2 _29611_ (.A(_07584_),
    .B(_07585_),
    .C(_07586_),
    .Y(_07587_));
 sky130_fd_sc_hd__nand2_2 _29612_ (.A(_07581_),
    .B(_07587_),
    .Y(_07588_));
 sky130_fd_sc_hd__a21boi_2 _29613_ (.A1(_07384_),
    .A2(_07373_),
    .B1_N(_07369_),
    .Y(_07589_));
 sky130_fd_sc_hd__buf_1 _29614_ (.A(\pcpi_mul.rs1[20] ),
    .X(_07590_));
 sky130_fd_sc_hd__nand2_2 _29615_ (.A(_05209_),
    .B(_07138_),
    .Y(_07591_));
 sky130_fd_sc_hd__a21o_2 _29616_ (.A1(_05143_),
    .A2(_07590_),
    .B1(_07591_),
    .X(_07592_));
 sky130_fd_sc_hd__buf_1 _29617_ (.A(\pcpi_mul.rs1[19] ),
    .X(_07593_));
 sky130_fd_sc_hd__buf_1 _29618_ (.A(\pcpi_mul.rs1[20] ),
    .X(_07594_));
 sky130_fd_sc_hd__nand2_2 _29619_ (.A(_19400_),
    .B(_07594_),
    .Y(_07595_));
 sky130_fd_sc_hd__a21o_2 _29620_ (.A1(_05203_),
    .A2(_07593_),
    .B1(_07595_),
    .X(_07596_));
 sky130_fd_sc_hd__nand2_2 _29621_ (.A(_19393_),
    .B(_07153_),
    .Y(_07597_));
 sky130_fd_sc_hd__a21oi_2 _29622_ (.A1(_07592_),
    .A2(_07596_),
    .B1(_07597_),
    .Y(_07598_));
 sky130_fd_sc_hd__and3_2 _29623_ (.A(_07592_),
    .B(_07596_),
    .C(_07597_),
    .X(_07599_));
 sky130_fd_sc_hd__nor2_2 _29624_ (.A(_07598_),
    .B(_07599_),
    .Y(_07600_));
 sky130_fd_sc_hd__nand2_2 _29625_ (.A(_05321_),
    .B(_07360_),
    .Y(_07601_));
 sky130_fd_sc_hd__nand2_2 _29626_ (.A(_05322_),
    .B(_19587_),
    .Y(_07602_));
 sky130_fd_sc_hd__nor2_2 _29627_ (.A(_07601_),
    .B(_07602_),
    .Y(_07603_));
 sky130_fd_sc_hd__and2_2 _29628_ (.A(_07601_),
    .B(_07602_),
    .X(_07604_));
 sky130_fd_sc_hd__buf_1 _29629_ (.A(\pcpi_mul.rs1[21] ),
    .X(_07605_));
 sky130_fd_sc_hd__nand2_2 _29630_ (.A(_19403_),
    .B(_07605_),
    .Y(_07606_));
 sky130_fd_sc_hd__o21ai_2 _29631_ (.A1(_07603_),
    .A2(_07604_),
    .B1(_07606_),
    .Y(_07607_));
 sky130_fd_sc_hd__or2_2 _29632_ (.A(_07601_),
    .B(_07602_),
    .X(_07608_));
 sky130_fd_sc_hd__inv_2 _29633_ (.A(_07606_),
    .Y(_07609_));
 sky130_fd_sc_hd__nand2_2 _29634_ (.A(_07601_),
    .B(_07602_),
    .Y(_07610_));
 sky130_fd_sc_hd__nand3_2 _29635_ (.A(_07608_),
    .B(_07609_),
    .C(_07610_),
    .Y(_07611_));
 sky130_fd_sc_hd__o21ai_2 _29636_ (.A1(_07361_),
    .A2(_07359_),
    .B1(_07365_),
    .Y(_07612_));
 sky130_fd_sc_hd__nand3_2 _29637_ (.A(_07607_),
    .B(_07611_),
    .C(_07612_),
    .Y(_07613_));
 sky130_fd_sc_hd__nor2_2 _29638_ (.A(_07367_),
    .B(_07362_),
    .Y(_07614_));
 sky130_fd_sc_hd__o21ai_2 _29639_ (.A1(_07603_),
    .A2(_07604_),
    .B1(_07609_),
    .Y(_07615_));
 sky130_fd_sc_hd__nand3_2 _29640_ (.A(_07608_),
    .B(_07606_),
    .C(_07610_),
    .Y(_07616_));
 sky130_fd_sc_hd__nand3_2 _29641_ (.A(_07614_),
    .B(_07615_),
    .C(_07616_),
    .Y(_07617_));
 sky130_fd_sc_hd__nand3b_2 _29642_ (.A_N(_07600_),
    .B(_07613_),
    .C(_07617_),
    .Y(_07618_));
 sky130_fd_sc_hd__nand2_2 _29643_ (.A(_07617_),
    .B(_07613_),
    .Y(_07619_));
 sky130_fd_sc_hd__nand2_2 _29644_ (.A(_07619_),
    .B(_07600_),
    .Y(_07620_));
 sky130_fd_sc_hd__and3_2 _29645_ (.A(_07589_),
    .B(_07618_),
    .C(_07620_),
    .X(_07621_));
 sky130_fd_sc_hd__a21bo_2 _29646_ (.A1(_07384_),
    .A2(_07373_),
    .B1_N(_07369_),
    .X(_07622_));
 sky130_fd_sc_hd__o21ai_2 _29647_ (.A1(_07599_),
    .A2(_07598_),
    .B1(_07619_),
    .Y(_07623_));
 sky130_fd_sc_hd__nand3_2 _29648_ (.A(_07600_),
    .B(_07613_),
    .C(_07617_),
    .Y(_07624_));
 sky130_fd_sc_hd__nand3_2 _29649_ (.A(_07622_),
    .B(_07623_),
    .C(_07624_),
    .Y(_07625_));
 sky130_fd_sc_hd__nor2_2 _29650_ (.A(_07375_),
    .B(_07378_),
    .Y(_07626_));
 sky130_fd_sc_hd__nor2_2 _29651_ (.A(_07626_),
    .B(_07382_),
    .Y(_07627_));
 sky130_fd_sc_hd__inv_2 _29652_ (.A(_07627_),
    .Y(_07628_));
 sky130_fd_sc_hd__nand2_2 _29653_ (.A(_07625_),
    .B(_07628_),
    .Y(_07629_));
 sky130_fd_sc_hd__nand3_2 _29654_ (.A(_07618_),
    .B(_07589_),
    .C(_07620_),
    .Y(_07630_));
 sky130_fd_sc_hd__nand2_2 _29655_ (.A(_07625_),
    .B(_07630_),
    .Y(_07631_));
 sky130_fd_sc_hd__nand2_2 _29656_ (.A(_07631_),
    .B(_07627_),
    .Y(_07632_));
 sky130_fd_sc_hd__o21ai_2 _29657_ (.A1(_07621_),
    .A2(_07629_),
    .B1(_07632_),
    .Y(_07633_));
 sky130_fd_sc_hd__nand2_2 _29658_ (.A(_07588_),
    .B(_07633_),
    .Y(_07634_));
 sky130_fd_sc_hd__inv_2 _29659_ (.A(_07474_),
    .Y(_07635_));
 sky130_fd_sc_hd__nand2_2 _29660_ (.A(_07631_),
    .B(_07628_),
    .Y(_07636_));
 sky130_fd_sc_hd__nand3_2 _29661_ (.A(_07625_),
    .B(_07630_),
    .C(_07627_),
    .Y(_07637_));
 sky130_fd_sc_hd__nand2_2 _29662_ (.A(_07636_),
    .B(_07637_),
    .Y(_07638_));
 sky130_fd_sc_hd__nand3_2 _29663_ (.A(_07638_),
    .B(_07581_),
    .C(_07587_),
    .Y(_07639_));
 sky130_fd_sc_hd__nand3_2 _29664_ (.A(_07634_),
    .B(_07635_),
    .C(_07639_),
    .Y(_07640_));
 sky130_fd_sc_hd__inv_2 _29665_ (.A(_07637_),
    .Y(_07641_));
 sky130_fd_sc_hd__and2_2 _29666_ (.A(_07631_),
    .B(_07628_),
    .X(_07642_));
 sky130_fd_sc_hd__o2bb2ai_2 _29667_ (.A1_N(_07587_),
    .A2_N(_07581_),
    .B1(_07641_),
    .B2(_07642_),
    .Y(_07643_));
 sky130_fd_sc_hd__nand3_2 _29668_ (.A(_07633_),
    .B(_07581_),
    .C(_07587_),
    .Y(_07644_));
 sky130_fd_sc_hd__nand3_2 _29669_ (.A(_07643_),
    .B(_07474_),
    .C(_07644_),
    .Y(_07645_));
 sky130_fd_sc_hd__nand2_2 _29670_ (.A(_07401_),
    .B(_07349_),
    .Y(_07646_));
 sky130_fd_sc_hd__a21oi_2 _29671_ (.A1(_07640_),
    .A2(_07645_),
    .B1(_07646_),
    .Y(_07647_));
 sky130_fd_sc_hd__inv_2 _29672_ (.A(_07349_),
    .Y(_07648_));
 sky130_fd_sc_hd__and3_2 _29673_ (.A(_07400_),
    .B(_07355_),
    .C(_07349_),
    .X(_07649_));
 sky130_fd_sc_hd__o211a_2 _29674_ (.A1(_07648_),
    .A2(_07649_),
    .B1(_07645_),
    .C1(_07640_),
    .X(_07650_));
 sky130_fd_sc_hd__buf_1 _29675_ (.A(_05266_),
    .X(_07651_));
 sky130_fd_sc_hd__buf_1 _29676_ (.A(_19356_),
    .X(_07652_));
 sky130_fd_sc_hd__a22o_2 _29677_ (.A1(_19354_),
    .A2(_19627_),
    .B1(_07652_),
    .B2(_19625_),
    .X(_07653_));
 sky130_fd_sc_hd__o21ai_2 _29678_ (.A1(_07651_),
    .A2(_07234_),
    .B1(_07653_),
    .Y(_07654_));
 sky130_fd_sc_hd__nand2_2 _29679_ (.A(\pcpi_mul.rs2[15] ),
    .B(_05251_),
    .Y(_07655_));
 sky130_fd_sc_hd__inv_2 _29680_ (.A(_07655_),
    .Y(_07656_));
 sky130_fd_sc_hd__nand2_2 _29681_ (.A(_07654_),
    .B(_07656_),
    .Y(_07657_));
 sky130_fd_sc_hd__o21ai_2 _29682_ (.A1(_07479_),
    .A2(_07484_),
    .B1(_07476_),
    .Y(_07658_));
 sky130_fd_sc_hd__nand2_2 _29683_ (.A(_07658_),
    .B(_07485_),
    .Y(_07659_));
 sky130_fd_sc_hd__o211ai_2 _29684_ (.A1(_07651_),
    .A2(_07234_),
    .B1(_07655_),
    .C1(_07653_),
    .Y(_07660_));
 sky130_fd_sc_hd__nand3_2 _29685_ (.A(_07657_),
    .B(_07659_),
    .C(_07660_),
    .Y(_07661_));
 sky130_fd_sc_hd__nand2_2 _29686_ (.A(_07654_),
    .B(_07655_),
    .Y(_07662_));
 sky130_fd_sc_hd__nor2_2 _29687_ (.A(_07651_),
    .B(_07234_),
    .Y(_07663_));
 sky130_fd_sc_hd__nand3b_2 _29688_ (.A_N(_07663_),
    .B(_07656_),
    .C(_07653_),
    .Y(_07664_));
 sky130_fd_sc_hd__nand2_2 _29689_ (.A(_07477_),
    .B(_07485_),
    .Y(_07665_));
 sky130_fd_sc_hd__nand2_2 _29690_ (.A(_07665_),
    .B(_07482_),
    .Y(_07666_));
 sky130_fd_sc_hd__nand3_2 _29691_ (.A(_07662_),
    .B(_07664_),
    .C(_07666_),
    .Y(_07667_));
 sky130_fd_sc_hd__nor2_2 _29692_ (.A(_07420_),
    .B(_07415_),
    .Y(_07668_));
 sky130_fd_sc_hd__o2bb2ai_2 _29693_ (.A1_N(_07661_),
    .A2_N(_07667_),
    .B1(_07422_),
    .B2(_07668_),
    .Y(_07669_));
 sky130_fd_sc_hd__a21oi_2 _29694_ (.A1(_07418_),
    .A2(_07420_),
    .B1(_07415_),
    .Y(_07670_));
 sky130_fd_sc_hd__inv_2 _29695_ (.A(_07670_),
    .Y(_07671_));
 sky130_fd_sc_hd__nand3_2 _29696_ (.A(_07667_),
    .B(_07661_),
    .C(_07671_),
    .Y(_07672_));
 sky130_fd_sc_hd__nand2_2 _29697_ (.A(_07427_),
    .B(_07428_),
    .Y(_07673_));
 sky130_fd_sc_hd__nand2_2 _29698_ (.A(_07673_),
    .B(_07424_),
    .Y(_07674_));
 sky130_fd_sc_hd__a21oi_2 _29699_ (.A1(_07669_),
    .A2(_07672_),
    .B1(_07674_),
    .Y(_07675_));
 sky130_fd_sc_hd__and3_2 _29700_ (.A(_07669_),
    .B(_07674_),
    .C(_07672_),
    .X(_07676_));
 sky130_fd_sc_hd__o21ai_2 _29701_ (.A1(_07445_),
    .A2(_07446_),
    .B1(_07448_),
    .Y(_07677_));
 sky130_fd_sc_hd__and2_2 _29702_ (.A(_07677_),
    .B(_07453_),
    .X(_07678_));
 sky130_fd_sc_hd__nand2_2 _29703_ (.A(_06269_),
    .B(_05419_),
    .Y(_07679_));
 sky130_fd_sc_hd__nand3b_2 _29704_ (.A_N(_07679_),
    .B(_07020_),
    .C(_06507_),
    .Y(_07680_));
 sky130_fd_sc_hd__nand2_2 _29705_ (.A(_06275_),
    .B(_05730_),
    .Y(_07681_));
 sky130_fd_sc_hd__nand2_2 _29706_ (.A(_07679_),
    .B(_07681_),
    .Y(_07682_));
 sky130_fd_sc_hd__nand2_2 _29707_ (.A(_06117_),
    .B(_19612_),
    .Y(_07683_));
 sky130_fd_sc_hd__inv_2 _29708_ (.A(_07683_),
    .Y(_07684_));
 sky130_fd_sc_hd__nand3_2 _29709_ (.A(_07680_),
    .B(_07682_),
    .C(_07684_),
    .Y(_07685_));
 sky130_fd_sc_hd__a22oi_2 _29710_ (.A1(_06270_),
    .A2(_05420_),
    .B1(_19365_),
    .B2(_06162_),
    .Y(_07686_));
 sky130_fd_sc_hd__nor2_2 _29711_ (.A(_07679_),
    .B(_07681_),
    .Y(_07687_));
 sky130_fd_sc_hd__o21ai_2 _29712_ (.A1(_07686_),
    .A2(_07687_),
    .B1(_07683_),
    .Y(_07688_));
 sky130_fd_sc_hd__nand3_2 _29713_ (.A(_07678_),
    .B(_07685_),
    .C(_07688_),
    .Y(_07689_));
 sky130_fd_sc_hd__o21ai_2 _29714_ (.A1(_07686_),
    .A2(_07687_),
    .B1(_07684_),
    .Y(_07690_));
 sky130_fd_sc_hd__nand3_2 _29715_ (.A(_07680_),
    .B(_07682_),
    .C(_07683_),
    .Y(_07691_));
 sky130_fd_sc_hd__nand2_2 _29716_ (.A(_07677_),
    .B(_07453_),
    .Y(_07692_));
 sky130_fd_sc_hd__nand3_2 _29717_ (.A(_07690_),
    .B(_07691_),
    .C(_07692_),
    .Y(_07693_));
 sky130_fd_sc_hd__nand2_2 _29718_ (.A(_06430_),
    .B(_19608_),
    .Y(_07694_));
 sky130_fd_sc_hd__nand2_2 _29719_ (.A(_06432_),
    .B(_19605_),
    .Y(_07695_));
 sky130_fd_sc_hd__nor2_2 _29720_ (.A(_07694_),
    .B(_07695_),
    .Y(_07696_));
 sky130_fd_sc_hd__nand2_2 _29721_ (.A(_19375_),
    .B(_07109_),
    .Y(_07697_));
 sky130_fd_sc_hd__a21o_2 _29722_ (.A1(_07694_),
    .A2(_07695_),
    .B1(_07697_),
    .X(_07698_));
 sky130_fd_sc_hd__a22oi_2 _29723_ (.A1(_07203_),
    .A2(_06889_),
    .B1(_06258_),
    .B2(_05717_),
    .Y(_07699_));
 sky130_fd_sc_hd__o21ai_2 _29724_ (.A1(_07699_),
    .A2(_07696_),
    .B1(_07697_),
    .Y(_07700_));
 sky130_fd_sc_hd__o21a_2 _29725_ (.A1(_07696_),
    .A2(_07698_),
    .B1(_07700_),
    .X(_07701_));
 sky130_fd_sc_hd__a21o_2 _29726_ (.A1(_07689_),
    .A2(_07693_),
    .B1(_07701_),
    .X(_07702_));
 sky130_fd_sc_hd__nand3_2 _29727_ (.A(_07689_),
    .B(_07701_),
    .C(_07693_),
    .Y(_07703_));
 sky130_fd_sc_hd__nand2_2 _29728_ (.A(_07702_),
    .B(_07703_),
    .Y(_07704_));
 sky130_fd_sc_hd__o21ai_2 _29729_ (.A1(_07675_),
    .A2(_07676_),
    .B1(_07704_),
    .Y(_07705_));
 sky130_fd_sc_hd__inv_2 _29730_ (.A(_07704_),
    .Y(_07706_));
 sky130_fd_sc_hd__a21o_2 _29731_ (.A1(_07669_),
    .A2(_07672_),
    .B1(_07674_),
    .X(_07707_));
 sky130_fd_sc_hd__nand3_2 _29732_ (.A(_07669_),
    .B(_07674_),
    .C(_07672_),
    .Y(_07708_));
 sky130_fd_sc_hd__nand3_2 _29733_ (.A(_07706_),
    .B(_07707_),
    .C(_07708_),
    .Y(_07709_));
 sky130_fd_sc_hd__nand2_2 _29734_ (.A(_07471_),
    .B(_07435_),
    .Y(_07710_));
 sky130_fd_sc_hd__nand3_2 _29735_ (.A(_07705_),
    .B(_07709_),
    .C(_07710_),
    .Y(_07711_));
 sky130_fd_sc_hd__buf_1 _29736_ (.A(_07711_),
    .X(_07712_));
 sky130_fd_sc_hd__o21ai_2 _29737_ (.A1(_07675_),
    .A2(_07676_),
    .B1(_07706_),
    .Y(_07713_));
 sky130_fd_sc_hd__a21oi_2 _29738_ (.A1(_07431_),
    .A2(_07463_),
    .B1(_07470_),
    .Y(_07714_));
 sky130_fd_sc_hd__nand3_2 _29739_ (.A(_07707_),
    .B(_07708_),
    .C(_07704_),
    .Y(_07715_));
 sky130_fd_sc_hd__nand3_2 _29740_ (.A(_07713_),
    .B(_07714_),
    .C(_07715_),
    .Y(_07716_));
 sky130_fd_sc_hd__inv_2 _29741_ (.A(\pcpi_mul.rs2[21] ),
    .Y(_07717_));
 sky130_fd_sc_hd__buf_1 _29742_ (.A(_07717_),
    .X(_07718_));
 sky130_fd_sc_hd__nor2_2 _29743_ (.A(_07718_),
    .B(_04838_),
    .Y(_07719_));
 sky130_fd_sc_hd__nand2_2 _29744_ (.A(\pcpi_mul.rs2[18] ),
    .B(_05218_),
    .Y(_07720_));
 sky130_fd_sc_hd__inv_2 _29745_ (.A(_07720_),
    .Y(_07721_));
 sky130_fd_sc_hd__buf_1 _29746_ (.A(\pcpi_mul.rs2[20] ),
    .X(_07722_));
 sky130_fd_sc_hd__buf_1 _29747_ (.A(\pcpi_mul.rs2[19] ),
    .X(_07723_));
 sky130_fd_sc_hd__a22oi_2 _29748_ (.A1(_07722_),
    .A2(_05190_),
    .B1(_07723_),
    .B2(_05545_),
    .Y(_07724_));
 sky130_fd_sc_hd__and4_2 _29749_ (.A(_07480_),
    .B(_19349_),
    .C(_05248_),
    .D(_19635_),
    .X(_07725_));
 sky130_fd_sc_hd__nor2_2 _29750_ (.A(_07724_),
    .B(_07725_),
    .Y(_07726_));
 sky130_fd_sc_hd__or2_2 _29751_ (.A(_07721_),
    .B(_07726_),
    .X(_07727_));
 sky130_fd_sc_hd__nand2_2 _29752_ (.A(_07726_),
    .B(_07721_),
    .Y(_07728_));
 sky130_fd_sc_hd__nand2_2 _29753_ (.A(_07727_),
    .B(_07728_),
    .Y(_07729_));
 sky130_fd_sc_hd__nor2_2 _29754_ (.A(_07719_),
    .B(_07729_),
    .Y(_07730_));
 sky130_fd_sc_hd__and2_2 _29755_ (.A(_07729_),
    .B(_07719_),
    .X(_07731_));
 sky130_fd_sc_hd__nor2_2 _29756_ (.A(_07730_),
    .B(_07731_),
    .Y(_07732_));
 sky130_fd_sc_hd__inv_2 _29757_ (.A(_07732_),
    .Y(_07733_));
 sky130_fd_sc_hd__a21oi_2 _29758_ (.A1(_07712_),
    .A2(_07716_),
    .B1(_07733_),
    .Y(_07734_));
 sky130_fd_sc_hd__and3_2 _29759_ (.A(_07712_),
    .B(_07716_),
    .C(_07733_),
    .X(_07735_));
 sky130_fd_sc_hd__o21ai_2 _29760_ (.A1(_07734_),
    .A2(_07735_),
    .B1(_07498_),
    .Y(_07736_));
 sky130_fd_sc_hd__a21o_2 _29761_ (.A1(_07712_),
    .A2(_07716_),
    .B1(_07733_),
    .X(_07737_));
 sky130_fd_sc_hd__nand3_2 _29762_ (.A(_07712_),
    .B(_07716_),
    .C(_07733_),
    .Y(_07738_));
 sky130_fd_sc_hd__nand3_2 _29763_ (.A(_07493_),
    .B(_07737_),
    .C(_07738_),
    .Y(_07739_));
 sky130_fd_sc_hd__nand2_2 _29764_ (.A(_07736_),
    .B(_07739_),
    .Y(_07740_));
 sky130_fd_sc_hd__o21ai_2 _29765_ (.A1(_07647_),
    .A2(_07650_),
    .B1(_07740_),
    .Y(_07741_));
 sky130_fd_sc_hd__nor2_2 _29766_ (.A(_07498_),
    .B(_07734_),
    .Y(_07742_));
 sky130_fd_sc_hd__a21oi_2 _29767_ (.A1(_07737_),
    .A2(_07738_),
    .B1(_07493_),
    .Y(_07743_));
 sky130_fd_sc_hd__a21oi_2 _29768_ (.A1(_07742_),
    .A2(_07738_),
    .B1(_07743_),
    .Y(_07744_));
 sky130_fd_sc_hd__a21o_2 _29769_ (.A1(_07640_),
    .A2(_07645_),
    .B1(_07646_),
    .X(_07745_));
 sky130_fd_sc_hd__nand3_2 _29770_ (.A(_07640_),
    .B(_07645_),
    .C(_07646_),
    .Y(_07746_));
 sky130_fd_sc_hd__nand3_2 _29771_ (.A(_07744_),
    .B(_07745_),
    .C(_07746_),
    .Y(_07747_));
 sky130_fd_sc_hd__nand3_2 _29772_ (.A(_07550_),
    .B(_07741_),
    .C(_07747_),
    .Y(_07748_));
 sky130_fd_sc_hd__o21ai_2 _29773_ (.A1(_07647_),
    .A2(_07650_),
    .B1(_07744_),
    .Y(_07749_));
 sky130_fd_sc_hd__nor2_2 _29774_ (.A(_07493_),
    .B(_07502_),
    .Y(_07750_));
 sky130_fd_sc_hd__a31oi_2 _29775_ (.A1(_07409_),
    .A2(_07494_),
    .A3(_07503_),
    .B1(_07750_),
    .Y(_07751_));
 sky130_fd_sc_hd__nand3_2 _29776_ (.A(_07745_),
    .B(_07740_),
    .C(_07746_),
    .Y(_07752_));
 sky130_fd_sc_hd__nand3_2 _29777_ (.A(_07749_),
    .B(_07751_),
    .C(_07752_),
    .Y(_07753_));
 sky130_fd_sc_hd__nand2_2 _29778_ (.A(_07748_),
    .B(_07753_),
    .Y(_07754_));
 sky130_fd_sc_hd__inv_2 _29779_ (.A(_07399_),
    .Y(_07755_));
 sky130_fd_sc_hd__nand2_2 _29780_ (.A(_07755_),
    .B(_07391_),
    .Y(_07756_));
 sky130_fd_sc_hd__inv_2 _29781_ (.A(_07756_),
    .Y(_07757_));
 sky130_fd_sc_hd__a21o_2 _29782_ (.A1(_07411_),
    .A2(_07403_),
    .B1(_07757_),
    .X(_07758_));
 sky130_fd_sc_hd__nand3_2 _29783_ (.A(_07503_),
    .B(_07403_),
    .C(_07757_),
    .Y(_07759_));
 sky130_fd_sc_hd__nand2_2 _29784_ (.A(_07758_),
    .B(_07759_),
    .Y(_07760_));
 sky130_fd_sc_hd__nand2_2 _29785_ (.A(_07754_),
    .B(_07760_),
    .Y(_07761_));
 sky130_fd_sc_hd__and2_2 _29786_ (.A(_07758_),
    .B(_07759_),
    .X(_07762_));
 sky130_fd_sc_hd__nand3_2 _29787_ (.A(_07748_),
    .B(_07753_),
    .C(_07762_),
    .Y(_07763_));
 sky130_fd_sc_hd__nand3_2 _29788_ (.A(_07549_),
    .B(_07761_),
    .C(_07763_),
    .Y(_07764_));
 sky130_fd_sc_hd__a21boi_2 _29789_ (.A1(_07513_),
    .A2(_07519_),
    .B1_N(_07505_),
    .Y(_07765_));
 sky130_fd_sc_hd__and2_2 _29790_ (.A(_07503_),
    .B(_07403_),
    .X(_07766_));
 sky130_fd_sc_hd__nor2_2 _29791_ (.A(_07756_),
    .B(_07766_),
    .Y(_07767_));
 sky130_fd_sc_hd__and3_2 _29792_ (.A(_07503_),
    .B(_07403_),
    .C(_07756_),
    .X(_07768_));
 sky130_fd_sc_hd__o2bb2ai_2 _29793_ (.A1_N(_07753_),
    .A2_N(_07748_),
    .B1(_07767_),
    .B2(_07768_),
    .Y(_07769_));
 sky130_fd_sc_hd__nand3_2 _29794_ (.A(_07748_),
    .B(_07753_),
    .C(_07760_),
    .Y(_07770_));
 sky130_fd_sc_hd__nand3_2 _29795_ (.A(_07765_),
    .B(_07769_),
    .C(_07770_),
    .Y(_07771_));
 sky130_fd_sc_hd__a21oi_2 _29796_ (.A1(_07764_),
    .A2(_07771_),
    .B1(_07516_),
    .Y(_07772_));
 sky130_fd_sc_hd__and3_2 _29797_ (.A(_07764_),
    .B(_07771_),
    .C(_07516_),
    .X(_07773_));
 sky130_fd_sc_hd__a21oi_2 _29798_ (.A1(_07529_),
    .A2(_07530_),
    .B1(_07532_),
    .Y(_07774_));
 sky130_fd_sc_hd__nor2_2 _29799_ (.A(_07526_),
    .B(_07774_),
    .Y(_07775_));
 sky130_fd_sc_hd__o21ai_2 _29800_ (.A1(_07772_),
    .A2(_07773_),
    .B1(_07775_),
    .Y(_07776_));
 sky130_fd_sc_hd__o21ai_2 _29801_ (.A1(_07532_),
    .A2(_07523_),
    .B1(_07533_),
    .Y(_07777_));
 sky130_fd_sc_hd__nand2_2 _29802_ (.A(_07764_),
    .B(_07771_),
    .Y(_07778_));
 sky130_fd_sc_hd__inv_2 _29803_ (.A(_07516_),
    .Y(_07779_));
 sky130_fd_sc_hd__nand2_2 _29804_ (.A(_07778_),
    .B(_07779_),
    .Y(_07780_));
 sky130_fd_sc_hd__nand3_2 _29805_ (.A(_07764_),
    .B(_07771_),
    .C(_07516_),
    .Y(_07781_));
 sky130_fd_sc_hd__nand3_2 _29806_ (.A(_07777_),
    .B(_07780_),
    .C(_07781_),
    .Y(_07782_));
 sky130_fd_sc_hd__nand2_2 _29807_ (.A(_07776_),
    .B(_07782_),
    .Y(_07783_));
 sky130_fd_sc_hd__nand2_2 _29808_ (.A(_07548_),
    .B(_07540_),
    .Y(_07784_));
 sky130_fd_sc_hd__nand2_2 _29809_ (.A(_07784_),
    .B(_07535_),
    .Y(_07785_));
 sky130_fd_sc_hd__xor2_2 _29810_ (.A(_07783_),
    .B(_07785_),
    .X(_02640_));
 sky130_fd_sc_hd__inv_2 _29811_ (.A(_07688_),
    .Y(_07786_));
 sky130_fd_sc_hd__nand2_2 _29812_ (.A(_07678_),
    .B(_07685_),
    .Y(_07787_));
 sky130_fd_sc_hd__o2bb2ai_2 _29813_ (.A1_N(_07693_),
    .A2_N(_07701_),
    .B1(_07786_),
    .B2(_07787_),
    .Y(_07788_));
 sky130_fd_sc_hd__a22oi_2 _29814_ (.A1(_19380_),
    .A2(_07143_),
    .B1(_06896_),
    .B2(_06748_),
    .Y(_07789_));
 sky130_fd_sc_hd__nand3_2 _29815_ (.A(_05639_),
    .B(_06010_),
    .C(_19596_),
    .Y(_07790_));
 sky130_fd_sc_hd__nor2_2 _29816_ (.A(_06958_),
    .B(_07790_),
    .Y(_07791_));
 sky130_fd_sc_hd__nand2_2 _29817_ (.A(_06496_),
    .B(_07360_),
    .Y(_07792_));
 sky130_fd_sc_hd__o21ai_2 _29818_ (.A1(_07789_),
    .A2(_07791_),
    .B1(_07792_),
    .Y(_07793_));
 sky130_fd_sc_hd__nand3b_2 _29819_ (.A_N(_07694_),
    .B(_19374_),
    .C(_19607_),
    .Y(_07794_));
 sky130_fd_sc_hd__nand2_2 _29820_ (.A(_07698_),
    .B(_07794_),
    .Y(_07795_));
 sky130_fd_sc_hd__inv_2 _29821_ (.A(_07792_),
    .Y(_07796_));
 sky130_fd_sc_hd__buf_1 _29822_ (.A(_05639_),
    .X(_07797_));
 sky130_fd_sc_hd__buf_1 _29823_ (.A(_06372_),
    .X(_07798_));
 sky130_fd_sc_hd__a22o_2 _29824_ (.A1(_07797_),
    .A2(_19597_),
    .B1(_06896_),
    .B2(_07798_),
    .X(_07799_));
 sky130_fd_sc_hd__o211ai_2 _29825_ (.A1(_06959_),
    .A2(_07790_),
    .B1(_07796_),
    .C1(_07799_),
    .Y(_07800_));
 sky130_fd_sc_hd__nand3_2 _29826_ (.A(_07793_),
    .B(_07795_),
    .C(_07800_),
    .Y(_07801_));
 sky130_fd_sc_hd__o21ai_2 _29827_ (.A1(_07789_),
    .A2(_07791_),
    .B1(_07796_),
    .Y(_07802_));
 sky130_fd_sc_hd__nand2_2 _29828_ (.A(_07694_),
    .B(_07695_),
    .Y(_07803_));
 sky130_fd_sc_hd__a31oi_2 _29829_ (.A1(_07803_),
    .A2(_06020_),
    .A3(_06073_),
    .B1(_07696_),
    .Y(_07804_));
 sky130_fd_sc_hd__o211ai_2 _29830_ (.A1(_06958_),
    .A2(_07790_),
    .B1(_07792_),
    .C1(_07799_),
    .Y(_07805_));
 sky130_fd_sc_hd__nand3_2 _29831_ (.A(_07802_),
    .B(_07804_),
    .C(_07805_),
    .Y(_07806_));
 sky130_fd_sc_hd__nor2_2 _29832_ (.A(_07556_),
    .B(_07554_),
    .Y(_07807_));
 sky130_fd_sc_hd__o2bb2ai_2 _29833_ (.A1_N(_07801_),
    .A2_N(_07806_),
    .B1(_07552_),
    .B2(_07807_),
    .Y(_07808_));
 sky130_fd_sc_hd__nor2_2 _29834_ (.A(_07552_),
    .B(_07807_),
    .Y(_07809_));
 sky130_fd_sc_hd__nand3_2 _29835_ (.A(_07806_),
    .B(_07801_),
    .C(_07809_),
    .Y(_07810_));
 sky130_fd_sc_hd__nand3_2 _29836_ (.A(_07788_),
    .B(_07808_),
    .C(_07810_),
    .Y(_07811_));
 sky130_fd_sc_hd__inv_2 _29837_ (.A(_07693_),
    .Y(_07812_));
 sky130_fd_sc_hd__a31oi_2 _29838_ (.A1(_07678_),
    .A2(_07685_),
    .A3(_07688_),
    .B1(_07701_),
    .Y(_07813_));
 sky130_fd_sc_hd__o2bb2ai_2 _29839_ (.A1_N(_07810_),
    .A2_N(_07808_),
    .B1(_07812_),
    .B2(_07813_),
    .Y(_07814_));
 sky130_fd_sc_hd__inv_2 _29840_ (.A(_07567_),
    .Y(_07815_));
 sky130_fd_sc_hd__and2_2 _29841_ (.A(_07561_),
    .B(_07568_),
    .X(_07816_));
 sky130_fd_sc_hd__o2bb2ai_2 _29842_ (.A1_N(_07811_),
    .A2_N(_07814_),
    .B1(_07815_),
    .B2(_07816_),
    .Y(_07817_));
 sky130_fd_sc_hd__nand2_2 _29843_ (.A(_07571_),
    .B(_07579_),
    .Y(_07818_));
 sky130_fd_sc_hd__nand2_2 _29844_ (.A(_07818_),
    .B(_07575_),
    .Y(_07819_));
 sky130_fd_sc_hd__nor2_2 _29845_ (.A(_07815_),
    .B(_07816_),
    .Y(_07820_));
 sky130_fd_sc_hd__nand3_2 _29846_ (.A(_07814_),
    .B(_07811_),
    .C(_07820_),
    .Y(_07821_));
 sky130_fd_sc_hd__nand3_2 _29847_ (.A(_07817_),
    .B(_07819_),
    .C(_07821_),
    .Y(_07822_));
 sky130_fd_sc_hd__inv_2 _29848_ (.A(_07561_),
    .Y(_07823_));
 sky130_fd_sc_hd__nor2_2 _29849_ (.A(_07568_),
    .B(_07815_),
    .Y(_07824_));
 sky130_fd_sc_hd__o2bb2ai_2 _29850_ (.A1_N(_07811_),
    .A2_N(_07814_),
    .B1(_07823_),
    .B2(_07824_),
    .Y(_07825_));
 sky130_fd_sc_hd__nand2_2 _29851_ (.A(_07551_),
    .B(_07569_),
    .Y(_07826_));
 sky130_fd_sc_hd__a21oi_2 _29852_ (.A1(_07569_),
    .A2(_07570_),
    .B1(_07551_),
    .Y(_07827_));
 sky130_fd_sc_hd__o22ai_2 _29853_ (.A1(_07574_),
    .A2(_07826_),
    .B1(_07579_),
    .B2(_07827_),
    .Y(_07828_));
 sky130_fd_sc_hd__nand3b_2 _29854_ (.A_N(_07820_),
    .B(_07814_),
    .C(_07811_),
    .Y(_07829_));
 sky130_fd_sc_hd__nand3_2 _29855_ (.A(_07825_),
    .B(_07828_),
    .C(_07829_),
    .Y(_07830_));
 sky130_fd_sc_hd__nand2_2 _29856_ (.A(_07822_),
    .B(_07830_),
    .Y(_07831_));
 sky130_fd_sc_hd__inv_2 _29857_ (.A(\pcpi_mul.rs1[17] ),
    .Y(_07832_));
 sky130_fd_sc_hd__buf_1 _29858_ (.A(_07832_),
    .X(_07833_));
 sky130_fd_sc_hd__nand3_2 _29859_ (.A(_06199_),
    .B(_06201_),
    .C(_07153_),
    .Y(_07834_));
 sky130_fd_sc_hd__a22o_2 _29860_ (.A1(_06731_),
    .A2(_19588_),
    .B1(_05891_),
    .B2(_07156_),
    .X(_07835_));
 sky130_fd_sc_hd__o21ai_2 _29861_ (.A1(_07833_),
    .A2(_07834_),
    .B1(_07835_),
    .Y(_07836_));
 sky130_fd_sc_hd__buf_1 _29862_ (.A(\pcpi_mul.rs1[22] ),
    .X(_07837_));
 sky130_fd_sc_hd__nand2_2 _29863_ (.A(_19403_),
    .B(_07837_),
    .Y(_07838_));
 sky130_fd_sc_hd__nand2_2 _29864_ (.A(_07836_),
    .B(_07838_),
    .Y(_07839_));
 sky130_fd_sc_hd__inv_2 _29865_ (.A(_07838_),
    .Y(_07840_));
 sky130_fd_sc_hd__o211ai_2 _29866_ (.A1(_07833_),
    .A2(_07834_),
    .B1(_07840_),
    .C1(_07835_),
    .Y(_07841_));
 sky130_fd_sc_hd__a21o_2 _29867_ (.A1(_07609_),
    .A2(_07610_),
    .B1(_07603_),
    .X(_07842_));
 sky130_fd_sc_hd__a21oi_2 _29868_ (.A1(_07839_),
    .A2(_07841_),
    .B1(_07842_),
    .Y(_07843_));
 sky130_fd_sc_hd__and3_2 _29869_ (.A(_07839_),
    .B(_07842_),
    .C(_07841_),
    .X(_07844_));
 sky130_fd_sc_hd__buf_1 _29870_ (.A(_19577_),
    .X(_07845_));
 sky130_fd_sc_hd__nand2_2 _29871_ (.A(_05736_),
    .B(_19580_),
    .Y(_07846_));
 sky130_fd_sc_hd__a21o_2 _29872_ (.A1(_06220_),
    .A2(_07845_),
    .B1(_07846_),
    .X(_07847_));
 sky130_fd_sc_hd__buf_1 _29873_ (.A(_07358_),
    .X(_07848_));
 sky130_fd_sc_hd__buf_1 _29874_ (.A(_07605_),
    .X(_07849_));
 sky130_fd_sc_hd__nand2_2 _29875_ (.A(_05205_),
    .B(_07849_),
    .Y(_07850_));
 sky130_fd_sc_hd__a21o_2 _29876_ (.A1(_06072_),
    .A2(_07848_),
    .B1(_07850_),
    .X(_07851_));
 sky130_fd_sc_hd__buf_1 _29877_ (.A(_07377_),
    .X(_07852_));
 sky130_fd_sc_hd__nand2_2 _29878_ (.A(_19394_),
    .B(_07852_),
    .Y(_07853_));
 sky130_fd_sc_hd__a21o_2 _29879_ (.A1(_07847_),
    .A2(_07851_),
    .B1(_07853_),
    .X(_07854_));
 sky130_fd_sc_hd__nand3_2 _29880_ (.A(_07847_),
    .B(_07851_),
    .C(_07853_),
    .Y(_07855_));
 sky130_fd_sc_hd__nand2_2 _29881_ (.A(_07854_),
    .B(_07855_),
    .Y(_07856_));
 sky130_fd_sc_hd__o21ai_2 _29882_ (.A1(_07843_),
    .A2(_07844_),
    .B1(_07856_),
    .Y(_07857_));
 sky130_fd_sc_hd__inv_2 _29883_ (.A(_07607_),
    .Y(_07858_));
 sky130_fd_sc_hd__nand2_2 _29884_ (.A(_07611_),
    .B(_07612_),
    .Y(_07859_));
 sky130_fd_sc_hd__o2bb2ai_2 _29885_ (.A1_N(_07617_),
    .A2_N(_07600_),
    .B1(_07858_),
    .B2(_07859_),
    .Y(_07860_));
 sky130_fd_sc_hd__and2_2 _29886_ (.A(_07854_),
    .B(_07855_),
    .X(_07861_));
 sky130_fd_sc_hd__a21o_2 _29887_ (.A1(_07839_),
    .A2(_07841_),
    .B1(_07842_),
    .X(_07862_));
 sky130_fd_sc_hd__nand3_2 _29888_ (.A(_07839_),
    .B(_07842_),
    .C(_07841_),
    .Y(_07863_));
 sky130_fd_sc_hd__nand3_2 _29889_ (.A(_07861_),
    .B(_07862_),
    .C(_07863_),
    .Y(_07864_));
 sky130_fd_sc_hd__nand3_2 _29890_ (.A(_07857_),
    .B(_07860_),
    .C(_07864_),
    .Y(_07865_));
 sky130_fd_sc_hd__o21ai_2 _29891_ (.A1(_07843_),
    .A2(_07844_),
    .B1(_07861_),
    .Y(_07866_));
 sky130_fd_sc_hd__a21boi_2 _29892_ (.A1(_07600_),
    .A2(_07617_),
    .B1_N(_07613_),
    .Y(_07867_));
 sky130_fd_sc_hd__nand3_2 _29893_ (.A(_07862_),
    .B(_07856_),
    .C(_07863_),
    .Y(_07868_));
 sky130_fd_sc_hd__o21ba_2 _29894_ (.A1(_07591_),
    .A2(_07595_),
    .B1_N(_07598_),
    .X(_07869_));
 sky130_fd_sc_hd__a31oi_2 _29895_ (.A1(_07866_),
    .A2(_07867_),
    .A3(_07868_),
    .B1(_07869_),
    .Y(_07870_));
 sky130_fd_sc_hd__nand3_2 _29896_ (.A(_07866_),
    .B(_07867_),
    .C(_07868_),
    .Y(_07871_));
 sky130_fd_sc_hd__a21boi_2 _29897_ (.A1(_07865_),
    .A2(_07871_),
    .B1_N(_07869_),
    .Y(_07872_));
 sky130_fd_sc_hd__a21oi_2 _29898_ (.A1(_07865_),
    .A2(_07870_),
    .B1(_07872_),
    .Y(_07873_));
 sky130_fd_sc_hd__nand2_2 _29899_ (.A(_07831_),
    .B(_07873_),
    .Y(_07874_));
 sky130_fd_sc_hd__nand2_2 _29900_ (.A(_07865_),
    .B(_07871_),
    .Y(_07875_));
 sky130_fd_sc_hd__nor2_2 _29901_ (.A(_07869_),
    .B(_07875_),
    .Y(_07876_));
 sky130_fd_sc_hd__o211ai_2 _29902_ (.A1(_07872_),
    .A2(_07876_),
    .B1(_07822_),
    .C1(_07830_),
    .Y(_07877_));
 sky130_fd_sc_hd__nand3_2 _29903_ (.A(_07874_),
    .B(_07712_),
    .C(_07877_),
    .Y(_07878_));
 sky130_fd_sc_hd__o2bb2ai_2 _29904_ (.A1_N(_07830_),
    .A2_N(_07822_),
    .B1(_07876_),
    .B2(_07872_),
    .Y(_07879_));
 sky130_fd_sc_hd__nand3_2 _29905_ (.A(_07873_),
    .B(_07822_),
    .C(_07830_),
    .Y(_07880_));
 sky130_fd_sc_hd__inv_2 _29906_ (.A(_07711_),
    .Y(_07881_));
 sky130_fd_sc_hd__nand3_2 _29907_ (.A(_07879_),
    .B(_07880_),
    .C(_07881_),
    .Y(_07882_));
 sky130_fd_sc_hd__a21bo_2 _29908_ (.A1(_07638_),
    .A2(_07581_),
    .B1_N(_07587_),
    .X(_07883_));
 sky130_fd_sc_hd__a21oi_2 _29909_ (.A1(_07878_),
    .A2(_07882_),
    .B1(_07883_),
    .Y(_07884_));
 sky130_fd_sc_hd__and3_2 _29910_ (.A(_07878_),
    .B(_07882_),
    .C(_07883_),
    .X(_07885_));
 sky130_fd_sc_hd__buf_1 _29911_ (.A(_07236_),
    .X(_07886_));
 sky130_fd_sc_hd__a22oi_2 _29912_ (.A1(_07886_),
    .A2(_05765_),
    .B1(_06824_),
    .B2(_06606_),
    .Y(_07887_));
 sky130_fd_sc_hd__nand3_2 _29913_ (.A(_07416_),
    .B(_07417_),
    .C(_05184_),
    .Y(_07888_));
 sky130_fd_sc_hd__nor2_2 _29914_ (.A(_05261_),
    .B(_07888_),
    .Y(_07889_));
 sky130_fd_sc_hd__buf_1 _29915_ (.A(\pcpi_mul.rs2[15] ),
    .X(_07890_));
 sky130_fd_sc_hd__nand2_2 _29916_ (.A(_07890_),
    .B(_05420_),
    .Y(_07891_));
 sky130_fd_sc_hd__inv_2 _29917_ (.A(_07891_),
    .Y(_07892_));
 sky130_fd_sc_hd__o21ai_2 _29918_ (.A1(_07887_),
    .A2(_07889_),
    .B1(_07892_),
    .Y(_07893_));
 sky130_fd_sc_hd__buf_1 _29919_ (.A(_19346_),
    .X(_07894_));
 sky130_fd_sc_hd__buf_1 _29920_ (.A(_19349_),
    .X(_07895_));
 sky130_fd_sc_hd__a22o_2 _29921_ (.A1(_07894_),
    .A2(_19636_),
    .B1(_07895_),
    .B2(_19633_),
    .X(_07896_));
 sky130_fd_sc_hd__a21oi_2 _29922_ (.A1(_07896_),
    .A2(_07721_),
    .B1(_07725_),
    .Y(_07897_));
 sky130_fd_sc_hd__buf_1 _29923_ (.A(_07236_),
    .X(_07898_));
 sky130_fd_sc_hd__a22o_2 _29924_ (.A1(_07898_),
    .A2(_05269_),
    .B1(_06824_),
    .B2(_06606_),
    .X(_07899_));
 sky130_fd_sc_hd__o211ai_2 _29925_ (.A1(_05501_),
    .A2(_07888_),
    .B1(_07891_),
    .C1(_07899_),
    .Y(_07900_));
 sky130_fd_sc_hd__nand3_2 _29926_ (.A(_07893_),
    .B(_07897_),
    .C(_07900_),
    .Y(_07901_));
 sky130_fd_sc_hd__o21ai_2 _29927_ (.A1(_07887_),
    .A2(_07889_),
    .B1(_07891_),
    .Y(_07902_));
 sky130_fd_sc_hd__buf_1 _29928_ (.A(_19346_),
    .X(_07903_));
 sky130_fd_sc_hd__buf_1 _29929_ (.A(_05104_),
    .X(_07904_));
 sky130_fd_sc_hd__nand2_2 _29930_ (.A(_07903_),
    .B(_07904_),
    .Y(_07905_));
 sky130_fd_sc_hd__buf_1 _29931_ (.A(\pcpi_mul.rs2[19] ),
    .X(_07906_));
 sky130_fd_sc_hd__buf_1 _29932_ (.A(_07906_),
    .X(_07907_));
 sky130_fd_sc_hd__nand3b_2 _29933_ (.A_N(_07905_),
    .B(_07907_),
    .C(_05120_),
    .Y(_07908_));
 sky130_fd_sc_hd__o21ai_2 _29934_ (.A1(_07720_),
    .A2(_07724_),
    .B1(_07908_),
    .Y(_07909_));
 sky130_fd_sc_hd__o211ai_2 _29935_ (.A1(_05501_),
    .A2(_07888_),
    .B1(_07892_),
    .C1(_07899_),
    .Y(_07910_));
 sky130_fd_sc_hd__nand3_2 _29936_ (.A(_07902_),
    .B(_07909_),
    .C(_07910_),
    .Y(_07911_));
 sky130_fd_sc_hd__a21oi_2 _29937_ (.A1(_07653_),
    .A2(_07656_),
    .B1(_07663_),
    .Y(_07912_));
 sky130_fd_sc_hd__inv_2 _29938_ (.A(_07912_),
    .Y(_07913_));
 sky130_fd_sc_hd__a21o_2 _29939_ (.A1(_07901_),
    .A2(_07911_),
    .B1(_07913_),
    .X(_07914_));
 sky130_fd_sc_hd__nand3_2 _29940_ (.A(_07901_),
    .B(_07911_),
    .C(_07913_),
    .Y(_07915_));
 sky130_fd_sc_hd__nand2_2 _29941_ (.A(_07661_),
    .B(_07671_),
    .Y(_07916_));
 sky130_fd_sc_hd__nand2_2 _29942_ (.A(_07916_),
    .B(_07667_),
    .Y(_07917_));
 sky130_fd_sc_hd__a21oi_2 _29943_ (.A1(_07914_),
    .A2(_07915_),
    .B1(_07917_),
    .Y(_07918_));
 sky130_fd_sc_hd__and3_2 _29944_ (.A(_07902_),
    .B(_07909_),
    .C(_07910_),
    .X(_07919_));
 sky130_fd_sc_hd__nand2_2 _29945_ (.A(_07901_),
    .B(_07913_),
    .Y(_07920_));
 sky130_fd_sc_hd__o211a_2 _29946_ (.A1(_07919_),
    .A2(_07920_),
    .B1(_07914_),
    .C1(_07917_),
    .X(_07921_));
 sky130_fd_sc_hd__nand2_2 _29947_ (.A(_19362_),
    .B(_05730_),
    .Y(_07922_));
 sky130_fd_sc_hd__nand2_2 _29948_ (.A(_06275_),
    .B(_05516_),
    .Y(_07923_));
 sky130_fd_sc_hd__nor2_2 _29949_ (.A(_07922_),
    .B(_07923_),
    .Y(_07924_));
 sky130_fd_sc_hd__nand2_2 _29950_ (.A(_19367_),
    .B(_19608_),
    .Y(_07925_));
 sky130_fd_sc_hd__inv_2 _29951_ (.A(_07925_),
    .Y(_07926_));
 sky130_fd_sc_hd__nand2_2 _29952_ (.A(_07922_),
    .B(_07923_),
    .Y(_07927_));
 sky130_fd_sc_hd__nand2_2 _29953_ (.A(_07926_),
    .B(_07927_),
    .Y(_07928_));
 sky130_fd_sc_hd__o21ai_2 _29954_ (.A1(_07679_),
    .A2(_07681_),
    .B1(_07683_),
    .Y(_07929_));
 sky130_fd_sc_hd__a22oi_2 _29955_ (.A1(_06441_),
    .A2(_06507_),
    .B1(_07020_),
    .B2(_06492_),
    .Y(_07930_));
 sky130_fd_sc_hd__o21ai_2 _29956_ (.A1(_07930_),
    .A2(_07924_),
    .B1(_07925_),
    .Y(_07931_));
 sky130_fd_sc_hd__o2111ai_2 _29957_ (.A1(_07924_),
    .A2(_07928_),
    .B1(_07682_),
    .C1(_07929_),
    .D1(_07931_),
    .Y(_07932_));
 sky130_fd_sc_hd__o21ai_2 _29958_ (.A1(_07930_),
    .A2(_07924_),
    .B1(_07926_),
    .Y(_07933_));
 sky130_fd_sc_hd__buf_1 _29959_ (.A(_07015_),
    .X(_07934_));
 sky130_fd_sc_hd__nand3b_2 _29960_ (.A_N(_07922_),
    .B(_07934_),
    .C(_05615_),
    .Y(_07935_));
 sky130_fd_sc_hd__nand3_2 _29961_ (.A(_07935_),
    .B(_07927_),
    .C(_07925_),
    .Y(_07936_));
 sky130_fd_sc_hd__nand2_2 _29962_ (.A(_07929_),
    .B(_07682_),
    .Y(_07937_));
 sky130_fd_sc_hd__nand3_2 _29963_ (.A(_07933_),
    .B(_07936_),
    .C(_07937_),
    .Y(_07938_));
 sky130_fd_sc_hd__buf_1 _29964_ (.A(_05896_),
    .X(_07939_));
 sky130_fd_sc_hd__a22oi_2 _29965_ (.A1(_07203_),
    .A2(_06369_),
    .B1(_06258_),
    .B2(_07939_),
    .Y(_07940_));
 sky130_fd_sc_hd__nand2_2 _29966_ (.A(_05955_),
    .B(_19605_),
    .Y(_07941_));
 sky130_fd_sc_hd__nand2_2 _29967_ (.A(_06432_),
    .B(_19602_),
    .Y(_07942_));
 sky130_fd_sc_hd__nor2_2 _29968_ (.A(_07941_),
    .B(_07942_),
    .Y(_07943_));
 sky130_fd_sc_hd__nand2_2 _29969_ (.A(_19375_),
    .B(_06058_),
    .Y(_07944_));
 sky130_fd_sc_hd__o21bai_2 _29970_ (.A1(_07940_),
    .A2(_07943_),
    .B1_N(_07944_),
    .Y(_07945_));
 sky130_fd_sc_hd__nand3b_2 _29971_ (.A_N(_07941_),
    .B(_06605_),
    .C(_06538_),
    .Y(_07946_));
 sky130_fd_sc_hd__nand2_2 _29972_ (.A(_07941_),
    .B(_07942_),
    .Y(_07947_));
 sky130_fd_sc_hd__nand3_2 _29973_ (.A(_07946_),
    .B(_07947_),
    .C(_07944_),
    .Y(_07948_));
 sky130_fd_sc_hd__nand2_2 _29974_ (.A(_07945_),
    .B(_07948_),
    .Y(_07949_));
 sky130_fd_sc_hd__a21oi_2 _29975_ (.A1(_07932_),
    .A2(_07938_),
    .B1(_07949_),
    .Y(_07950_));
 sky130_fd_sc_hd__and3_2 _29976_ (.A(_07932_),
    .B(_07938_),
    .C(_07949_),
    .X(_07951_));
 sky130_fd_sc_hd__nor2_2 _29977_ (.A(_07950_),
    .B(_07951_),
    .Y(_07952_));
 sky130_fd_sc_hd__o21ai_2 _29978_ (.A1(_07918_),
    .A2(_07921_),
    .B1(_07952_),
    .Y(_07953_));
 sky130_fd_sc_hd__nand2_2 _29979_ (.A(_07704_),
    .B(_07708_),
    .Y(_07954_));
 sky130_fd_sc_hd__nand2_2 _29980_ (.A(_07954_),
    .B(_07707_),
    .Y(_07955_));
 sky130_fd_sc_hd__a21o_2 _29981_ (.A1(_07914_),
    .A2(_07915_),
    .B1(_07917_),
    .X(_07956_));
 sky130_fd_sc_hd__and2_2 _29982_ (.A(_07932_),
    .B(_07949_),
    .X(_07957_));
 sky130_fd_sc_hd__a21o_2 _29983_ (.A1(_07957_),
    .A2(_07938_),
    .B1(_07950_),
    .X(_07958_));
 sky130_fd_sc_hd__nand3_2 _29984_ (.A(_07917_),
    .B(_07914_),
    .C(_07915_),
    .Y(_07959_));
 sky130_fd_sc_hd__nand3_2 _29985_ (.A(_07956_),
    .B(_07958_),
    .C(_07959_),
    .Y(_07960_));
 sky130_fd_sc_hd__nand3_2 _29986_ (.A(_07953_),
    .B(_07955_),
    .C(_07960_),
    .Y(_07961_));
 sky130_fd_sc_hd__o22ai_2 _29987_ (.A1(_07951_),
    .A2(_07950_),
    .B1(_07918_),
    .B2(_07921_),
    .Y(_07962_));
 sky130_fd_sc_hd__o21ai_2 _29988_ (.A1(_07704_),
    .A2(_07675_),
    .B1(_07708_),
    .Y(_07963_));
 sky130_fd_sc_hd__nand3_2 _29989_ (.A(_07956_),
    .B(_07959_),
    .C(_07952_),
    .Y(_07964_));
 sky130_fd_sc_hd__nand3_2 _29990_ (.A(_07962_),
    .B(_07963_),
    .C(_07964_),
    .Y(_07965_));
 sky130_fd_sc_hd__nand2_2 _29991_ (.A(_07475_),
    .B(_05212_),
    .Y(_07966_));
 sky130_fd_sc_hd__a22oi_2 _29992_ (.A1(_07903_),
    .A2(_05215_),
    .B1(_07895_),
    .B2(_19630_),
    .Y(_07967_));
 sky130_fd_sc_hd__nand2_2 _29993_ (.A(_19346_),
    .B(_05248_),
    .Y(_07968_));
 sky130_fd_sc_hd__nand2_2 _29994_ (.A(_07478_),
    .B(_06447_),
    .Y(_07969_));
 sky130_fd_sc_hd__nor2_2 _29995_ (.A(_07968_),
    .B(_07969_),
    .Y(_07970_));
 sky130_fd_sc_hd__or3_2 _29996_ (.A(_07966_),
    .B(_07967_),
    .C(_07970_),
    .X(_07971_));
 sky130_fd_sc_hd__o21ai_2 _29997_ (.A1(_07967_),
    .A2(_07970_),
    .B1(_07966_),
    .Y(_07972_));
 sky130_fd_sc_hd__nand2_2 _29998_ (.A(_07971_),
    .B(_07972_),
    .Y(_07973_));
 sky130_fd_sc_hd__buf_1 _29999_ (.A(\pcpi_mul.rs2[22] ),
    .X(_07974_));
 sky130_fd_sc_hd__nand2_2 _30000_ (.A(_07974_),
    .B(_19640_),
    .Y(_07975_));
 sky130_fd_sc_hd__buf_1 _30001_ (.A(\pcpi_mul.rs2[21] ),
    .X(_07976_));
 sky130_fd_sc_hd__nand2_2 _30002_ (.A(_07976_),
    .B(_19636_),
    .Y(_07977_));
 sky130_fd_sc_hd__or2_2 _30003_ (.A(_07975_),
    .B(_07977_),
    .X(_07978_));
 sky130_fd_sc_hd__nand2_2 _30004_ (.A(_07975_),
    .B(_07977_),
    .Y(_07979_));
 sky130_fd_sc_hd__nand2_2 _30005_ (.A(_07978_),
    .B(_07979_),
    .Y(_07980_));
 sky130_fd_sc_hd__nand2_2 _30006_ (.A(_07973_),
    .B(_07980_),
    .Y(_07981_));
 sky130_fd_sc_hd__nand3b_2 _30007_ (.A_N(_07980_),
    .B(_07971_),
    .C(_07972_),
    .Y(_07982_));
 sky130_fd_sc_hd__and3_2 _30008_ (.A(_07727_),
    .B(_07719_),
    .C(_07728_),
    .X(_07983_));
 sky130_fd_sc_hd__a21oi_2 _30009_ (.A1(_07981_),
    .A2(_07982_),
    .B1(_07983_),
    .Y(_07984_));
 sky130_fd_sc_hd__nand3_2 _30010_ (.A(_07983_),
    .B(_07981_),
    .C(_07982_),
    .Y(_07985_));
 sky130_fd_sc_hd__inv_2 _30011_ (.A(_07985_),
    .Y(_07986_));
 sky130_fd_sc_hd__nor2_2 _30012_ (.A(_07984_),
    .B(_07986_),
    .Y(_07987_));
 sky130_fd_sc_hd__nand3_2 _30013_ (.A(_07961_),
    .B(_07965_),
    .C(_07987_),
    .Y(_07988_));
 sky130_fd_sc_hd__nand2_2 _30014_ (.A(_07961_),
    .B(_07965_),
    .Y(_07989_));
 sky130_fd_sc_hd__inv_2 _30015_ (.A(_07987_),
    .Y(_07990_));
 sky130_fd_sc_hd__a21oi_2 _30016_ (.A1(_07989_),
    .A2(_07990_),
    .B1(_07738_),
    .Y(_07991_));
 sky130_fd_sc_hd__a31oi_2 _30017_ (.A1(_07713_),
    .A2(_07714_),
    .A3(_07715_),
    .B1(_07732_),
    .Y(_07992_));
 sky130_fd_sc_hd__o2bb2ai_2 _30018_ (.A1_N(_07965_),
    .A2_N(_07961_),
    .B1(_07986_),
    .B2(_07984_),
    .Y(_07993_));
 sky130_fd_sc_hd__a22oi_2 _30019_ (.A1(_07712_),
    .A2(_07992_),
    .B1(_07993_),
    .B2(_07988_),
    .Y(_07994_));
 sky130_fd_sc_hd__a21oi_2 _30020_ (.A1(_07988_),
    .A2(_07991_),
    .B1(_07994_),
    .Y(_07995_));
 sky130_fd_sc_hd__o21bai_2 _30021_ (.A1(_07884_),
    .A2(_07885_),
    .B1_N(_07995_),
    .Y(_07996_));
 sky130_fd_sc_hd__a21o_2 _30022_ (.A1(_07878_),
    .A2(_07882_),
    .B1(_07883_),
    .X(_07997_));
 sky130_fd_sc_hd__nand3_2 _30023_ (.A(_07878_),
    .B(_07882_),
    .C(_07883_),
    .Y(_07998_));
 sky130_fd_sc_hd__nand3_2 _30024_ (.A(_07997_),
    .B(_07995_),
    .C(_07998_),
    .Y(_07999_));
 sky130_fd_sc_hd__nand2_2 _30025_ (.A(_07746_),
    .B(_07736_),
    .Y(_08000_));
 sky130_fd_sc_hd__o21ai_2 _30026_ (.A1(_07647_),
    .A2(_08000_),
    .B1(_07739_),
    .Y(_08001_));
 sky130_fd_sc_hd__a21oi_2 _30027_ (.A1(_07996_),
    .A2(_07999_),
    .B1(_08001_),
    .Y(_08002_));
 sky130_fd_sc_hd__nand2_2 _30028_ (.A(_07993_),
    .B(_07988_),
    .Y(_08003_));
 sky130_fd_sc_hd__nand2_2 _30029_ (.A(_08003_),
    .B(_07738_),
    .Y(_08004_));
 sky130_fd_sc_hd__nand2_2 _30030_ (.A(_07991_),
    .B(_07988_),
    .Y(_08005_));
 sky130_fd_sc_hd__nand3_2 _30031_ (.A(_07998_),
    .B(_08004_),
    .C(_08005_),
    .Y(_08006_));
 sky130_fd_sc_hd__o211a_2 _30032_ (.A1(_07884_),
    .A2(_08006_),
    .B1(_07996_),
    .C1(_08001_),
    .X(_08007_));
 sky130_fd_sc_hd__nand2_2 _30033_ (.A(_07746_),
    .B(_07640_),
    .Y(_08008_));
 sky130_fd_sc_hd__o21ai_2 _30034_ (.A1(_07627_),
    .A2(_07621_),
    .B1(_07625_),
    .Y(_08009_));
 sky130_fd_sc_hd__nand2_2 _30035_ (.A(_08008_),
    .B(_08009_),
    .Y(_08010_));
 sky130_fd_sc_hd__nand3b_2 _30036_ (.A_N(_08009_),
    .B(_07746_),
    .C(_07640_),
    .Y(_08011_));
 sky130_fd_sc_hd__nand2_2 _30037_ (.A(_08010_),
    .B(_08011_),
    .Y(_08012_));
 sky130_fd_sc_hd__o21ai_2 _30038_ (.A1(_08002_),
    .A2(_08007_),
    .B1(_08012_),
    .Y(_08013_));
 sky130_fd_sc_hd__nand2_2 _30039_ (.A(_07996_),
    .B(_07999_),
    .Y(_08014_));
 sky130_fd_sc_hd__o21a_2 _30040_ (.A1(_07647_),
    .A2(_08000_),
    .B1(_07739_),
    .X(_08015_));
 sky130_fd_sc_hd__nand2_2 _30041_ (.A(_08014_),
    .B(_08015_),
    .Y(_08016_));
 sky130_fd_sc_hd__nand3_2 _30042_ (.A(_08001_),
    .B(_07996_),
    .C(_07999_),
    .Y(_08017_));
 sky130_fd_sc_hd__inv_2 _30043_ (.A(_08012_),
    .Y(_08018_));
 sky130_fd_sc_hd__nand3_2 _30044_ (.A(_08016_),
    .B(_08017_),
    .C(_08018_),
    .Y(_08019_));
 sky130_fd_sc_hd__nand2_2 _30045_ (.A(_08013_),
    .B(_08019_),
    .Y(_08020_));
 sky130_fd_sc_hd__inv_2 _30046_ (.A(_07748_),
    .Y(_08021_));
 sky130_fd_sc_hd__and2_2 _30047_ (.A(_07753_),
    .B(_07762_),
    .X(_08022_));
 sky130_fd_sc_hd__nor2_2 _30048_ (.A(_08021_),
    .B(_08022_),
    .Y(_08023_));
 sky130_fd_sc_hd__nand2_2 _30049_ (.A(_08020_),
    .B(_08023_),
    .Y(_08024_));
 sky130_fd_sc_hd__inv_2 _30050_ (.A(_07758_),
    .Y(_08025_));
 sky130_fd_sc_hd__a21bo_2 _30051_ (.A1(_07753_),
    .A2(_07762_),
    .B1_N(_07748_),
    .X(_08026_));
 sky130_fd_sc_hd__nand3_2 _30052_ (.A(_08026_),
    .B(_08013_),
    .C(_08019_),
    .Y(_08027_));
 sky130_fd_sc_hd__nand3_2 _30053_ (.A(_08024_),
    .B(_08025_),
    .C(_08027_),
    .Y(_08028_));
 sky130_fd_sc_hd__nand2_2 _30054_ (.A(_08024_),
    .B(_08027_),
    .Y(_08029_));
 sky130_fd_sc_hd__nand2_2 _30055_ (.A(_07771_),
    .B(_07516_),
    .Y(_08030_));
 sky130_fd_sc_hd__nand2_2 _30056_ (.A(_08030_),
    .B(_07764_),
    .Y(_08031_));
 sky130_fd_sc_hd__a21boi_2 _30057_ (.A1(_08029_),
    .A2(_07758_),
    .B1_N(_08031_),
    .Y(_08032_));
 sky130_fd_sc_hd__a21oi_2 _30058_ (.A1(_08013_),
    .A2(_08019_),
    .B1(_08026_),
    .Y(_08033_));
 sky130_fd_sc_hd__o211a_2 _30059_ (.A1(_08021_),
    .A2(_08022_),
    .B1(_08019_),
    .C1(_08013_),
    .X(_08034_));
 sky130_fd_sc_hd__o22ai_2 _30060_ (.A1(_07757_),
    .A2(_07766_),
    .B1(_08033_),
    .B2(_08034_),
    .Y(_08035_));
 sky130_fd_sc_hd__a21oi_2 _30061_ (.A1(_08035_),
    .A2(_08028_),
    .B1(_08031_),
    .Y(_08036_));
 sky130_fd_sc_hd__a21oi_2 _30062_ (.A1(_08028_),
    .A2(_08032_),
    .B1(_08036_),
    .Y(_08037_));
 sky130_fd_sc_hd__a21oi_2 _30063_ (.A1(_07780_),
    .A2(_07781_),
    .B1(_07777_),
    .Y(_08038_));
 sky130_fd_sc_hd__a21oi_2 _30064_ (.A1(_07540_),
    .A2(_07782_),
    .B1(_08038_),
    .Y(_08039_));
 sky130_fd_sc_hd__o22ai_2 _30065_ (.A1(_07779_),
    .A2(_07778_),
    .B1(_07526_),
    .B2(_07774_),
    .Y(_08040_));
 sky130_fd_sc_hd__o2111ai_2 _30066_ (.A1(_07772_),
    .A2(_08040_),
    .B1(_07535_),
    .C1(_07540_),
    .D1(_07776_),
    .Y(_08041_));
 sky130_fd_sc_hd__nor2_2 _30067_ (.A(_08041_),
    .B(_07548_),
    .Y(_08042_));
 sky130_fd_sc_hd__nor2_2 _30068_ (.A(_08039_),
    .B(_08042_),
    .Y(_08043_));
 sky130_fd_sc_hd__xnor2_2 _30069_ (.A(_08037_),
    .B(_08043_),
    .Y(_02641_));
 sky130_fd_sc_hd__a22oi_2 _30070_ (.A1(_05758_),
    .A2(_06957_),
    .B1(_05760_),
    .B2(_06949_),
    .Y(_08044_));
 sky130_fd_sc_hd__inv_2 _30071_ (.A(\pcpi_mul.rs1[16] ),
    .Y(_08045_));
 sky130_fd_sc_hd__nand3_2 _30072_ (.A(_06008_),
    .B(_06334_),
    .C(_19593_),
    .Y(_08046_));
 sky130_fd_sc_hd__nor2_2 _30073_ (.A(_08045_),
    .B(_08046_),
    .Y(_08047_));
 sky130_fd_sc_hd__nand2_2 _30074_ (.A(_05763_),
    .B(_19587_),
    .Y(_08048_));
 sky130_fd_sc_hd__inv_2 _30075_ (.A(_08048_),
    .Y(_08049_));
 sky130_fd_sc_hd__o21ai_2 _30076_ (.A1(_08044_),
    .A2(_08047_),
    .B1(_08049_),
    .Y(_08050_));
 sky130_fd_sc_hd__o21ai_2 _30077_ (.A1(_07941_),
    .A2(_07942_),
    .B1(_07944_),
    .Y(_08051_));
 sky130_fd_sc_hd__nand2_2 _30078_ (.A(_08051_),
    .B(_07947_),
    .Y(_08052_));
 sky130_fd_sc_hd__buf_1 _30079_ (.A(_08045_),
    .X(_08053_));
 sky130_fd_sc_hd__a22o_2 _30080_ (.A1(_05542_),
    .A2(_06373_),
    .B1(_19383_),
    .B2(_06946_),
    .X(_08054_));
 sky130_fd_sc_hd__o211ai_2 _30081_ (.A1(_08053_),
    .A2(_08046_),
    .B1(_08048_),
    .C1(_08054_),
    .Y(_08055_));
 sky130_fd_sc_hd__nand3_2 _30082_ (.A(_08050_),
    .B(_08052_),
    .C(_08055_),
    .Y(_08056_));
 sky130_fd_sc_hd__o21ai_2 _30083_ (.A1(_08044_),
    .A2(_08047_),
    .B1(_08048_),
    .Y(_08057_));
 sky130_fd_sc_hd__o21ai_2 _30084_ (.A1(_07944_),
    .A2(_07940_),
    .B1(_07946_),
    .Y(_08058_));
 sky130_fd_sc_hd__o211ai_2 _30085_ (.A1(_08053_),
    .A2(_08046_),
    .B1(_08049_),
    .C1(_08054_),
    .Y(_08059_));
 sky130_fd_sc_hd__nand3_2 _30086_ (.A(_08057_),
    .B(_08058_),
    .C(_08059_),
    .Y(_08060_));
 sky130_fd_sc_hd__nor2_2 _30087_ (.A(_07796_),
    .B(_07791_),
    .Y(_08061_));
 sky130_fd_sc_hd__o2bb2ai_2 _30088_ (.A1_N(_08056_),
    .A2_N(_08060_),
    .B1(_07789_),
    .B2(_08061_),
    .Y(_08062_));
 sky130_fd_sc_hd__nor2_2 _30089_ (.A(_07789_),
    .B(_08061_),
    .Y(_08063_));
 sky130_fd_sc_hd__nand3_2 _30090_ (.A(_08056_),
    .B(_08060_),
    .C(_08063_),
    .Y(_08064_));
 sky130_fd_sc_hd__nand2_2 _30091_ (.A(_07938_),
    .B(_07949_),
    .Y(_08065_));
 sky130_fd_sc_hd__nand2_2 _30092_ (.A(_08065_),
    .B(_07932_),
    .Y(_08066_));
 sky130_fd_sc_hd__a21oi_2 _30093_ (.A1(_08062_),
    .A2(_08064_),
    .B1(_08066_),
    .Y(_08067_));
 sky130_fd_sc_hd__and3_2 _30094_ (.A(_08057_),
    .B(_08058_),
    .C(_08059_),
    .X(_08068_));
 sky130_fd_sc_hd__nand2_2 _30095_ (.A(_08056_),
    .B(_08063_),
    .Y(_08069_));
 sky130_fd_sc_hd__o211a_2 _30096_ (.A1(_08068_),
    .A2(_08069_),
    .B1(_08062_),
    .C1(_08066_),
    .X(_08070_));
 sky130_fd_sc_hd__nand2_2 _30097_ (.A(_07806_),
    .B(_07809_),
    .Y(_08071_));
 sky130_fd_sc_hd__and2_2 _30098_ (.A(_08071_),
    .B(_07801_),
    .X(_08072_));
 sky130_fd_sc_hd__o21bai_2 _30099_ (.A1(_08067_),
    .A2(_08070_),
    .B1_N(_08072_),
    .Y(_08073_));
 sky130_fd_sc_hd__nand2_2 _30100_ (.A(_07811_),
    .B(_07820_),
    .Y(_08074_));
 sky130_fd_sc_hd__nand2_2 _30101_ (.A(_08074_),
    .B(_07814_),
    .Y(_08075_));
 sky130_fd_sc_hd__a21o_2 _30102_ (.A1(_08062_),
    .A2(_08064_),
    .B1(_08066_),
    .X(_08076_));
 sky130_fd_sc_hd__nand3_2 _30103_ (.A(_08066_),
    .B(_08062_),
    .C(_08064_),
    .Y(_08077_));
 sky130_fd_sc_hd__nand3_2 _30104_ (.A(_08076_),
    .B(_08077_),
    .C(_08072_),
    .Y(_08078_));
 sky130_fd_sc_hd__nand3_2 _30105_ (.A(_08073_),
    .B(_08075_),
    .C(_08078_),
    .Y(_08079_));
 sky130_fd_sc_hd__o21ai_2 _30106_ (.A1(_08067_),
    .A2(_08070_),
    .B1(_08072_),
    .Y(_08080_));
 sky130_fd_sc_hd__a21oi_2 _30107_ (.A1(_07808_),
    .A2(_07810_),
    .B1(_07788_),
    .Y(_08081_));
 sky130_fd_sc_hd__o21ai_2 _30108_ (.A1(_07820_),
    .A2(_08081_),
    .B1(_07811_),
    .Y(_08082_));
 sky130_fd_sc_hd__nand3b_2 _30109_ (.A_N(_08072_),
    .B(_08076_),
    .C(_08077_),
    .Y(_08083_));
 sky130_fd_sc_hd__nand3_2 _30110_ (.A(_08080_),
    .B(_08082_),
    .C(_08083_),
    .Y(_08084_));
 sky130_fd_sc_hd__buf_1 _30111_ (.A(\pcpi_mul.rs1[23] ),
    .X(_08085_));
 sky130_fd_sc_hd__nand2_2 _30112_ (.A(_05192_),
    .B(_08085_),
    .Y(_08086_));
 sky130_fd_sc_hd__a22oi_2 _30113_ (.A1(_05180_),
    .A2(_19584_),
    .B1(_05155_),
    .B2(_07138_),
    .Y(_08087_));
 sky130_fd_sc_hd__nor2_2 _30114_ (.A(_08086_),
    .B(_08087_),
    .Y(_08088_));
 sky130_fd_sc_hd__buf_1 _30115_ (.A(\pcpi_mul.rs1[18] ),
    .X(_08089_));
 sky130_fd_sc_hd__nand2_2 _30116_ (.A(_06731_),
    .B(_08089_),
    .Y(_08090_));
 sky130_fd_sc_hd__nand2_2 _30117_ (.A(_05189_),
    .B(_07138_),
    .Y(_08091_));
 sky130_fd_sc_hd__or2_2 _30118_ (.A(_08090_),
    .B(_08091_),
    .X(_08092_));
 sky130_fd_sc_hd__nand2_2 _30119_ (.A(_08088_),
    .B(_08092_),
    .Y(_08093_));
 sky130_fd_sc_hd__o2bb2ai_2 _30120_ (.A1_N(_07835_),
    .A2_N(_07840_),
    .B1(_07833_),
    .B2(_07834_),
    .Y(_08094_));
 sky130_fd_sc_hd__nor2_2 _30121_ (.A(_08090_),
    .B(_08091_),
    .Y(_08095_));
 sky130_fd_sc_hd__o21ai_2 _30122_ (.A1(_08087_),
    .A2(_08095_),
    .B1(_08086_),
    .Y(_08096_));
 sky130_fd_sc_hd__nand3_2 _30123_ (.A(_08093_),
    .B(_08094_),
    .C(_08096_),
    .Y(_08097_));
 sky130_fd_sc_hd__inv_2 _30124_ (.A(_08087_),
    .Y(_08098_));
 sky130_fd_sc_hd__nand3_2 _30125_ (.A(_08092_),
    .B(_08098_),
    .C(_08086_),
    .Y(_08099_));
 sky130_fd_sc_hd__a2bb2oi_2 _30126_ (.A1_N(_07833_),
    .A2_N(_07834_),
    .B1(_07840_),
    .B2(_07835_),
    .Y(_08100_));
 sky130_fd_sc_hd__o21bai_2 _30127_ (.A1(_08087_),
    .A2(_08095_),
    .B1_N(_08086_),
    .Y(_08101_));
 sky130_fd_sc_hd__nand3_2 _30128_ (.A(_08099_),
    .B(_08100_),
    .C(_08101_),
    .Y(_08102_));
 sky130_fd_sc_hd__buf_1 _30129_ (.A(_07837_),
    .X(_08103_));
 sky130_fd_sc_hd__nand2_2 _30130_ (.A(_05209_),
    .B(_19577_),
    .Y(_08104_));
 sky130_fd_sc_hd__a21o_2 _30131_ (.A1(_05143_),
    .A2(_08103_),
    .B1(_08104_),
    .X(_08105_));
 sky130_fd_sc_hd__nand2_2 _30132_ (.A(_05210_),
    .B(_19573_),
    .Y(_08106_));
 sky130_fd_sc_hd__a21o_2 _30133_ (.A1(_19398_),
    .A2(_07849_),
    .B1(_08106_),
    .X(_08107_));
 sky130_fd_sc_hd__buf_1 _30134_ (.A(_07594_),
    .X(_08108_));
 sky130_fd_sc_hd__nand2_2 _30135_ (.A(_19393_),
    .B(_08108_),
    .Y(_08109_));
 sky130_fd_sc_hd__and3_2 _30136_ (.A(_08105_),
    .B(_08107_),
    .C(_08109_),
    .X(_08110_));
 sky130_fd_sc_hd__a21oi_2 _30137_ (.A1(_08105_),
    .A2(_08107_),
    .B1(_08109_),
    .Y(_08111_));
 sky130_fd_sc_hd__o2bb2ai_2 _30138_ (.A1_N(_08097_),
    .A2_N(_08102_),
    .B1(_08110_),
    .B2(_08111_),
    .Y(_08112_));
 sky130_fd_sc_hd__nor2_2 _30139_ (.A(_08111_),
    .B(_08110_),
    .Y(_08113_));
 sky130_fd_sc_hd__nand3_2 _30140_ (.A(_08113_),
    .B(_08097_),
    .C(_08102_),
    .Y(_08114_));
 sky130_fd_sc_hd__o21ai_2 _30141_ (.A1(_07856_),
    .A2(_07843_),
    .B1(_07863_),
    .Y(_08115_));
 sky130_fd_sc_hd__a21o_2 _30142_ (.A1(_08112_),
    .A2(_08114_),
    .B1(_08115_),
    .X(_08116_));
 sky130_fd_sc_hd__nand3_2 _30143_ (.A(_08115_),
    .B(_08112_),
    .C(_08114_),
    .Y(_08117_));
 sky130_fd_sc_hd__nor2_2 _30144_ (.A(_07846_),
    .B(_07850_),
    .Y(_08118_));
 sky130_fd_sc_hd__a21oi_2 _30145_ (.A1(_07847_),
    .A2(_07851_),
    .B1(_07853_),
    .Y(_08119_));
 sky130_fd_sc_hd__nor2_2 _30146_ (.A(_08118_),
    .B(_08119_),
    .Y(_08120_));
 sky130_fd_sc_hd__inv_2 _30147_ (.A(_08120_),
    .Y(_08121_));
 sky130_fd_sc_hd__a21oi_2 _30148_ (.A1(_08116_),
    .A2(_08117_),
    .B1(_08121_),
    .Y(_08122_));
 sky130_fd_sc_hd__and3_2 _30149_ (.A(_08116_),
    .B(_08121_),
    .C(_08117_),
    .X(_08123_));
 sky130_fd_sc_hd__o2bb2ai_2 _30150_ (.A1_N(_08079_),
    .A2_N(_08084_),
    .B1(_08122_),
    .B2(_08123_),
    .Y(_08124_));
 sky130_fd_sc_hd__a21oi_2 _30151_ (.A1(_08112_),
    .A2(_08114_),
    .B1(_08115_),
    .Y(_08125_));
 sky130_fd_sc_hd__inv_2 _30152_ (.A(_08097_),
    .Y(_08126_));
 sky130_fd_sc_hd__a21o_2 _30153_ (.A1(_08105_),
    .A2(_08107_),
    .B1(_08109_),
    .X(_08127_));
 sky130_fd_sc_hd__nand3b_2 _30154_ (.A_N(_08110_),
    .B(_08102_),
    .C(_08127_),
    .Y(_08128_));
 sky130_fd_sc_hd__o211a_2 _30155_ (.A1(_08126_),
    .A2(_08128_),
    .B1(_08112_),
    .C1(_08115_),
    .X(_08129_));
 sky130_fd_sc_hd__o21ai_2 _30156_ (.A1(_08125_),
    .A2(_08129_),
    .B1(_08121_),
    .Y(_08130_));
 sky130_fd_sc_hd__nand3_2 _30157_ (.A(_08116_),
    .B(_08120_),
    .C(_08117_),
    .Y(_08131_));
 sky130_fd_sc_hd__nand2_2 _30158_ (.A(_08130_),
    .B(_08131_),
    .Y(_08132_));
 sky130_fd_sc_hd__nand3_2 _30159_ (.A(_08132_),
    .B(_08084_),
    .C(_08079_),
    .Y(_08133_));
 sky130_fd_sc_hd__inv_2 _30160_ (.A(_07965_),
    .Y(_08134_));
 sky130_fd_sc_hd__a21oi_2 _30161_ (.A1(_08124_),
    .A2(_08133_),
    .B1(_08134_),
    .Y(_08135_));
 sky130_fd_sc_hd__and3_2 _30162_ (.A(_08080_),
    .B(_08082_),
    .C(_08083_),
    .X(_08136_));
 sky130_fd_sc_hd__nand2_2 _30163_ (.A(_08132_),
    .B(_08079_),
    .Y(_08137_));
 sky130_fd_sc_hd__o211a_2 _30164_ (.A1(_08136_),
    .A2(_08137_),
    .B1(_08134_),
    .C1(_08124_),
    .X(_08138_));
 sky130_fd_sc_hd__a21bo_2 _30165_ (.A1(_07873_),
    .A2(_07822_),
    .B1_N(_07830_),
    .X(_08139_));
 sky130_fd_sc_hd__o21bai_2 _30166_ (.A1(_08135_),
    .A2(_08138_),
    .B1_N(_08139_),
    .Y(_08140_));
 sky130_fd_sc_hd__a21o_2 _30167_ (.A1(_08124_),
    .A2(_08133_),
    .B1(_08134_),
    .X(_08141_));
 sky130_fd_sc_hd__nand3_2 _30168_ (.A(_08124_),
    .B(_08134_),
    .C(_08133_),
    .Y(_08142_));
 sky130_fd_sc_hd__nand3_2 _30169_ (.A(_08141_),
    .B(_08142_),
    .C(_08139_),
    .Y(_08143_));
 sky130_fd_sc_hd__nand2_2 _30170_ (.A(_08140_),
    .B(_08143_),
    .Y(_08144_));
 sky130_fd_sc_hd__nand2_2 _30171_ (.A(_19339_),
    .B(_19635_),
    .Y(_08145_));
 sky130_fd_sc_hd__nand2_2 _30172_ (.A(_19336_),
    .B(_19639_),
    .Y(_08146_));
 sky130_fd_sc_hd__nor2_2 _30173_ (.A(_08145_),
    .B(_08146_),
    .Y(_08147_));
 sky130_fd_sc_hd__and2_2 _30174_ (.A(_08145_),
    .B(_08146_),
    .X(_08148_));
 sky130_fd_sc_hd__nand2_2 _30175_ (.A(\pcpi_mul.rs2[21] ),
    .B(_05248_),
    .Y(_08149_));
 sky130_fd_sc_hd__o21ai_2 _30176_ (.A1(_08147_),
    .A2(_08148_),
    .B1(_08149_),
    .Y(_08150_));
 sky130_fd_sc_hd__or2_2 _30177_ (.A(_08145_),
    .B(_08146_),
    .X(_08151_));
 sky130_fd_sc_hd__inv_2 _30178_ (.A(_08149_),
    .Y(_08152_));
 sky130_fd_sc_hd__nand2_2 _30179_ (.A(_08145_),
    .B(_08146_),
    .Y(_08153_));
 sky130_fd_sc_hd__nand3_2 _30180_ (.A(_08151_),
    .B(_08152_),
    .C(_08153_),
    .Y(_08154_));
 sky130_fd_sc_hd__nand3b_2 _30181_ (.A_N(_07978_),
    .B(_08150_),
    .C(_08154_),
    .Y(_08155_));
 sky130_fd_sc_hd__o21ai_2 _30182_ (.A1(_08147_),
    .A2(_08148_),
    .B1(_08152_),
    .Y(_08156_));
 sky130_fd_sc_hd__nand3_2 _30183_ (.A(_08151_),
    .B(_08149_),
    .C(_08153_),
    .Y(_08157_));
 sky130_fd_sc_hd__nand3_2 _30184_ (.A(_08156_),
    .B(_08157_),
    .C(_07978_),
    .Y(_08158_));
 sky130_fd_sc_hd__buf_1 _30185_ (.A(\pcpi_mul.rs2[19] ),
    .X(_08159_));
 sky130_fd_sc_hd__a22oi_2 _30186_ (.A1(_07903_),
    .A2(_19630_),
    .B1(_08159_),
    .B2(_06629_),
    .Y(_08160_));
 sky130_fd_sc_hd__nand3_2 _30187_ (.A(_07483_),
    .B(_07906_),
    .C(_06447_),
    .Y(_08161_));
 sky130_fd_sc_hd__nor2_2 _30188_ (.A(_06105_),
    .B(_08161_),
    .Y(_08162_));
 sky130_fd_sc_hd__a211o_2 _30189_ (.A1(_19352_),
    .A2(_19626_),
    .B1(_08160_),
    .C1(_08162_),
    .X(_08163_));
 sky130_fd_sc_hd__nand2_2 _30190_ (.A(_07475_),
    .B(_05345_),
    .Y(_08164_));
 sky130_fd_sc_hd__inv_2 _30191_ (.A(_08164_),
    .Y(_08165_));
 sky130_fd_sc_hd__o21ai_2 _30192_ (.A1(_08160_),
    .A2(_08162_),
    .B1(_08165_),
    .Y(_08166_));
 sky130_fd_sc_hd__nand2_2 _30193_ (.A(_08163_),
    .B(_08166_),
    .Y(_08167_));
 sky130_fd_sc_hd__a21o_2 _30194_ (.A1(_08155_),
    .A2(_08158_),
    .B1(_08167_),
    .X(_08168_));
 sky130_fd_sc_hd__nand3_2 _30195_ (.A(_08155_),
    .B(_08167_),
    .C(_08158_),
    .Y(_08169_));
 sky130_fd_sc_hd__nand2_2 _30196_ (.A(_08168_),
    .B(_08169_),
    .Y(_08170_));
 sky130_fd_sc_hd__nor2_2 _30197_ (.A(_07982_),
    .B(_08170_),
    .Y(_08171_));
 sky130_fd_sc_hd__inv_2 _30198_ (.A(_07982_),
    .Y(_08172_));
 sky130_fd_sc_hd__inv_2 _30199_ (.A(_08170_),
    .Y(_08173_));
 sky130_fd_sc_hd__nor2_2 _30200_ (.A(_08172_),
    .B(_08173_),
    .Y(_08174_));
 sky130_fd_sc_hd__nand2_2 _30201_ (.A(_07911_),
    .B(_07912_),
    .Y(_08175_));
 sky130_fd_sc_hd__a22oi_2 _30202_ (.A1(_07416_),
    .A2(_05347_),
    .B1(_07652_),
    .B2(_06808_),
    .Y(_08176_));
 sky130_fd_sc_hd__nand3_2 _30203_ (.A(_06821_),
    .B(_06827_),
    .C(_05342_),
    .Y(_08177_));
 sky130_fd_sc_hd__nor2_2 _30204_ (.A(_06332_),
    .B(_08177_),
    .Y(_08178_));
 sky130_fd_sc_hd__nand2_2 _30205_ (.A(\pcpi_mul.rs2[15] ),
    .B(_05730_),
    .Y(_08179_));
 sky130_fd_sc_hd__o21ai_2 _30206_ (.A1(_08176_),
    .A2(_08178_),
    .B1(_08179_),
    .Y(_08180_));
 sky130_fd_sc_hd__inv_2 _30207_ (.A(_08179_),
    .Y(_08181_));
 sky130_fd_sc_hd__buf_1 _30208_ (.A(_07236_),
    .X(_08182_));
 sky130_fd_sc_hd__a22o_2 _30209_ (.A1(_08182_),
    .A2(_19622_),
    .B1(_19357_),
    .B2(_05426_),
    .X(_08183_));
 sky130_fd_sc_hd__o211ai_2 _30210_ (.A1(_06333_),
    .A2(_08177_),
    .B1(_08181_),
    .C1(_08183_),
    .Y(_08184_));
 sky130_fd_sc_hd__buf_1 _30211_ (.A(_07478_),
    .X(_08185_));
 sky130_fd_sc_hd__nand3b_2 _30212_ (.A_N(_07968_),
    .B(_08185_),
    .C(_05204_),
    .Y(_08186_));
 sky130_fd_sc_hd__o21ai_2 _30213_ (.A1(_07966_),
    .A2(_07967_),
    .B1(_08186_),
    .Y(_08187_));
 sky130_fd_sc_hd__nand3_2 _30214_ (.A(_08180_),
    .B(_08184_),
    .C(_08187_),
    .Y(_08188_));
 sky130_fd_sc_hd__o21ai_2 _30215_ (.A1(_08176_),
    .A2(_08178_),
    .B1(_08181_),
    .Y(_08189_));
 sky130_fd_sc_hd__o21ai_2 _30216_ (.A1(_07968_),
    .A2(_07969_),
    .B1(_07966_),
    .Y(_08190_));
 sky130_fd_sc_hd__nand2_2 _30217_ (.A(_07968_),
    .B(_07969_),
    .Y(_08191_));
 sky130_fd_sc_hd__nand2_2 _30218_ (.A(_08190_),
    .B(_08191_),
    .Y(_08192_));
 sky130_fd_sc_hd__o211ai_2 _30219_ (.A1(_06333_),
    .A2(_08177_),
    .B1(_08179_),
    .C1(_08183_),
    .Y(_08193_));
 sky130_fd_sc_hd__nand3_2 _30220_ (.A(_08189_),
    .B(_08192_),
    .C(_08193_),
    .Y(_08194_));
 sky130_fd_sc_hd__nor2_2 _30221_ (.A(_07892_),
    .B(_07889_),
    .Y(_08195_));
 sky130_fd_sc_hd__o2bb2ai_2 _30222_ (.A1_N(_08188_),
    .A2_N(_08194_),
    .B1(_07887_),
    .B2(_08195_),
    .Y(_08196_));
 sky130_fd_sc_hd__a21oi_2 _30223_ (.A1(_07899_),
    .A2(_07892_),
    .B1(_07889_),
    .Y(_08197_));
 sky130_fd_sc_hd__nand3b_2 _30224_ (.A_N(_08197_),
    .B(_08188_),
    .C(_08194_),
    .Y(_08198_));
 sky130_fd_sc_hd__a22oi_2 _30225_ (.A1(_07901_),
    .A2(_08175_),
    .B1(_08196_),
    .B2(_08198_),
    .Y(_08199_));
 sky130_fd_sc_hd__a31oi_2 _30226_ (.A1(_07893_),
    .A2(_07897_),
    .A3(_07900_),
    .B1(_07912_),
    .Y(_08200_));
 sky130_fd_sc_hd__o211a_2 _30227_ (.A1(_07919_),
    .A2(_08200_),
    .B1(_08198_),
    .C1(_08196_),
    .X(_08201_));
 sky130_fd_sc_hd__a22oi_2 _30228_ (.A1(_06270_),
    .A2(_19613_),
    .B1(_19365_),
    .B2(_06889_),
    .Y(_08202_));
 sky130_fd_sc_hd__nand2_2 _30229_ (.A(_06269_),
    .B(_19612_),
    .Y(_08203_));
 sky130_fd_sc_hd__nand2_2 _30230_ (.A(_06275_),
    .B(_05597_),
    .Y(_08204_));
 sky130_fd_sc_hd__nor2_2 _30231_ (.A(_08203_),
    .B(_08204_),
    .Y(_08205_));
 sky130_fd_sc_hd__nand2_2 _30232_ (.A(_19367_),
    .B(_05910_),
    .Y(_08206_));
 sky130_fd_sc_hd__o21bai_2 _30233_ (.A1(_08202_),
    .A2(_08205_),
    .B1_N(_08206_),
    .Y(_08207_));
 sky130_fd_sc_hd__nand3b_2 _30234_ (.A_N(_08203_),
    .B(_07020_),
    .C(_05733_),
    .Y(_08208_));
 sky130_fd_sc_hd__nand2_2 _30235_ (.A(_08203_),
    .B(_08204_),
    .Y(_08209_));
 sky130_fd_sc_hd__nand3_2 _30236_ (.A(_08208_),
    .B(_08209_),
    .C(_08206_),
    .Y(_08210_));
 sky130_fd_sc_hd__o21ai_2 _30237_ (.A1(_07922_),
    .A2(_07923_),
    .B1(_07925_),
    .Y(_08211_));
 sky130_fd_sc_hd__nand2_2 _30238_ (.A(_08211_),
    .B(_07927_),
    .Y(_08212_));
 sky130_fd_sc_hd__a21o_2 _30239_ (.A1(_08207_),
    .A2(_08210_),
    .B1(_08212_),
    .X(_08213_));
 sky130_fd_sc_hd__nand3_2 _30240_ (.A(_08207_),
    .B(_08210_),
    .C(_08212_),
    .Y(_08214_));
 sky130_fd_sc_hd__nand2_2 _30241_ (.A(_08213_),
    .B(_08214_),
    .Y(_08215_));
 sky130_fd_sc_hd__a22oi_2 _30242_ (.A1(_05956_),
    .A2(_06732_),
    .B1(_19373_),
    .B2(_07311_),
    .Y(_08216_));
 sky130_fd_sc_hd__nand2_2 _30243_ (.A(_05955_),
    .B(_05896_),
    .Y(_08217_));
 sky130_fd_sc_hd__buf_1 _30244_ (.A(\pcpi_mul.rs1[13] ),
    .X(_08218_));
 sky130_fd_sc_hd__nand2_2 _30245_ (.A(_05802_),
    .B(_08218_),
    .Y(_08219_));
 sky130_fd_sc_hd__nor2_2 _30246_ (.A(_08217_),
    .B(_08219_),
    .Y(_08220_));
 sky130_fd_sc_hd__nand2_2 _30247_ (.A(_05672_),
    .B(_06205_),
    .Y(_08221_));
 sky130_fd_sc_hd__inv_2 _30248_ (.A(_08221_),
    .Y(_08222_));
 sky130_fd_sc_hd__o21ai_2 _30249_ (.A1(_08216_),
    .A2(_08220_),
    .B1(_08222_),
    .Y(_08223_));
 sky130_fd_sc_hd__nand3b_2 _30250_ (.A_N(_08217_),
    .B(_05670_),
    .C(_19600_),
    .Y(_08224_));
 sky130_fd_sc_hd__nand2_2 _30251_ (.A(_08217_),
    .B(_08219_),
    .Y(_08225_));
 sky130_fd_sc_hd__nand3_2 _30252_ (.A(_08224_),
    .B(_08225_),
    .C(_08221_),
    .Y(_08226_));
 sky130_fd_sc_hd__nand2_2 _30253_ (.A(_08223_),
    .B(_08226_),
    .Y(_08227_));
 sky130_fd_sc_hd__inv_2 _30254_ (.A(_08227_),
    .Y(_08228_));
 sky130_fd_sc_hd__nand2_2 _30255_ (.A(_08215_),
    .B(_08228_),
    .Y(_08229_));
 sky130_fd_sc_hd__nand3_2 _30256_ (.A(_08213_),
    .B(_08214_),
    .C(_08227_),
    .Y(_08230_));
 sky130_fd_sc_hd__nand2_2 _30257_ (.A(_08229_),
    .B(_08230_),
    .Y(_08231_));
 sky130_fd_sc_hd__o21ai_2 _30258_ (.A1(_08199_),
    .A2(_08201_),
    .B1(_08231_),
    .Y(_08232_));
 sky130_fd_sc_hd__nand2_2 _30259_ (.A(_07920_),
    .B(_07911_),
    .Y(_08233_));
 sky130_fd_sc_hd__a21o_2 _30260_ (.A1(_08196_),
    .A2(_08198_),
    .B1(_08233_),
    .X(_08234_));
 sky130_fd_sc_hd__nand2_2 _30261_ (.A(_08215_),
    .B(_08227_),
    .Y(_08235_));
 sky130_fd_sc_hd__nand3_2 _30262_ (.A(_08228_),
    .B(_08213_),
    .C(_08214_),
    .Y(_08236_));
 sky130_fd_sc_hd__nand2_2 _30263_ (.A(_08235_),
    .B(_08236_),
    .Y(_08237_));
 sky130_fd_sc_hd__nand3_2 _30264_ (.A(_08233_),
    .B(_08196_),
    .C(_08198_),
    .Y(_08238_));
 sky130_fd_sc_hd__nand3_2 _30265_ (.A(_08234_),
    .B(_08237_),
    .C(_08238_),
    .Y(_08239_));
 sky130_fd_sc_hd__nand3_2 _30266_ (.A(_08232_),
    .B(_07986_),
    .C(_08239_),
    .Y(_08240_));
 sky130_fd_sc_hd__nor2_2 _30267_ (.A(_08227_),
    .B(_08215_),
    .Y(_08241_));
 sky130_fd_sc_hd__a21oi_2 _30268_ (.A1(_08213_),
    .A2(_08214_),
    .B1(_08228_),
    .Y(_08242_));
 sky130_fd_sc_hd__o22ai_2 _30269_ (.A1(_08241_),
    .A2(_08242_),
    .B1(_08199_),
    .B2(_08201_),
    .Y(_08243_));
 sky130_fd_sc_hd__nand3_2 _30270_ (.A(_08234_),
    .B(_08231_),
    .C(_08238_),
    .Y(_08244_));
 sky130_fd_sc_hd__nand3_2 _30271_ (.A(_08243_),
    .B(_08244_),
    .C(_07985_),
    .Y(_08245_));
 sky130_fd_sc_hd__o21ai_2 _30272_ (.A1(_07918_),
    .A2(_07958_),
    .B1(_07959_),
    .Y(_08246_));
 sky130_fd_sc_hd__a21oi_2 _30273_ (.A1(_08240_),
    .A2(_08245_),
    .B1(_08246_),
    .Y(_08247_));
 sky130_fd_sc_hd__nor2_2 _30274_ (.A(_07918_),
    .B(_07958_),
    .Y(_08248_));
 sky130_fd_sc_hd__o211a_2 _30275_ (.A1(_07921_),
    .A2(_08248_),
    .B1(_08245_),
    .C1(_08240_),
    .X(_08249_));
 sky130_fd_sc_hd__o22ai_2 _30276_ (.A1(_08171_),
    .A2(_08174_),
    .B1(_08247_),
    .B2(_08249_),
    .Y(_08250_));
 sky130_fd_sc_hd__nor2_2 _30277_ (.A(_08172_),
    .B(_08170_),
    .Y(_08251_));
 sky130_fd_sc_hd__nor2_2 _30278_ (.A(_07982_),
    .B(_08173_),
    .Y(_08252_));
 sky130_fd_sc_hd__nor2_2 _30279_ (.A(_08251_),
    .B(_08252_),
    .Y(_08253_));
 sky130_fd_sc_hd__nand2_2 _30280_ (.A(_08240_),
    .B(_08245_),
    .Y(_08254_));
 sky130_fd_sc_hd__a21oi_2 _30281_ (.A1(_07956_),
    .A2(_07952_),
    .B1(_07921_),
    .Y(_08255_));
 sky130_fd_sc_hd__nand2_2 _30282_ (.A(_08254_),
    .B(_08255_),
    .Y(_08256_));
 sky130_fd_sc_hd__nand3_2 _30283_ (.A(_08240_),
    .B(_08245_),
    .C(_08246_),
    .Y(_08257_));
 sky130_fd_sc_hd__nand3b_2 _30284_ (.A_N(_08253_),
    .B(_08256_),
    .C(_08257_),
    .Y(_08258_));
 sky130_fd_sc_hd__o2bb2ai_2 _30285_ (.A1_N(_08250_),
    .A2_N(_08258_),
    .B1(_07990_),
    .B2(_07989_),
    .Y(_08259_));
 sky130_fd_sc_hd__inv_2 _30286_ (.A(_07988_),
    .Y(_08260_));
 sky130_fd_sc_hd__nand3_2 _30287_ (.A(_08250_),
    .B(_08258_),
    .C(_08260_),
    .Y(_08261_));
 sky130_fd_sc_hd__nand3_2 _30288_ (.A(_08144_),
    .B(_08259_),
    .C(_08261_),
    .Y(_08262_));
 sky130_fd_sc_hd__a21oi_2 _30289_ (.A1(_08250_),
    .A2(_08258_),
    .B1(_08260_),
    .Y(_08263_));
 sky130_fd_sc_hd__o2bb2ai_2 _30290_ (.A1_N(_08255_),
    .A2_N(_08254_),
    .B1(_08251_),
    .B2(_08252_),
    .Y(_08264_));
 sky130_fd_sc_hd__o211a_2 _30291_ (.A1(_08249_),
    .A2(_08264_),
    .B1(_08260_),
    .C1(_08250_),
    .X(_08265_));
 sky130_fd_sc_hd__o211ai_2 _30292_ (.A1(_08263_),
    .A2(_08265_),
    .B1(_08143_),
    .C1(_08140_),
    .Y(_08266_));
 sky130_fd_sc_hd__inv_2 _30293_ (.A(_08005_),
    .Y(_08267_));
 sky130_fd_sc_hd__a31oi_2 _30294_ (.A1(_07997_),
    .A2(_08004_),
    .A3(_07998_),
    .B1(_08267_),
    .Y(_08268_));
 sky130_fd_sc_hd__nand3_2 _30295_ (.A(_08262_),
    .B(_08266_),
    .C(_08268_),
    .Y(_08269_));
 sky130_fd_sc_hd__o2bb2ai_2 _30296_ (.A1_N(_08143_),
    .A2_N(_08140_),
    .B1(_08263_),
    .B2(_08265_),
    .Y(_08270_));
 sky130_fd_sc_hd__nand2_2 _30297_ (.A(_08142_),
    .B(_08139_),
    .Y(_08271_));
 sky130_fd_sc_hd__o2111ai_2 _30298_ (.A1(_08135_),
    .A2(_08271_),
    .B1(_08261_),
    .C1(_08259_),
    .D1(_08140_),
    .Y(_08272_));
 sky130_fd_sc_hd__o22ai_2 _30299_ (.A1(_07738_),
    .A2(_08003_),
    .B1(_07884_),
    .B2(_08006_),
    .Y(_08273_));
 sky130_fd_sc_hd__nand3_2 _30300_ (.A(_08270_),
    .B(_08272_),
    .C(_08273_),
    .Y(_08274_));
 sky130_fd_sc_hd__nand2_2 _30301_ (.A(_08269_),
    .B(_08274_),
    .Y(_08275_));
 sky130_fd_sc_hd__nand2_2 _30302_ (.A(_07998_),
    .B(_07882_),
    .Y(_08276_));
 sky130_fd_sc_hd__inv_2 _30303_ (.A(_07870_),
    .Y(_08277_));
 sky130_fd_sc_hd__nand2_2 _30304_ (.A(_08277_),
    .B(_07865_),
    .Y(_08278_));
 sky130_fd_sc_hd__nand2_2 _30305_ (.A(_08276_),
    .B(_08278_),
    .Y(_08279_));
 sky130_fd_sc_hd__inv_2 _30306_ (.A(_08278_),
    .Y(_08280_));
 sky130_fd_sc_hd__nand3_2 _30307_ (.A(_07998_),
    .B(_07882_),
    .C(_08280_),
    .Y(_08281_));
 sky130_fd_sc_hd__and2_2 _30308_ (.A(_08279_),
    .B(_08281_),
    .X(_08282_));
 sky130_fd_sc_hd__nand2_2 _30309_ (.A(_08275_),
    .B(_08282_),
    .Y(_08283_));
 sky130_fd_sc_hd__a21oi_2 _30310_ (.A1(_08016_),
    .A2(_08018_),
    .B1(_08007_),
    .Y(_08284_));
 sky130_fd_sc_hd__nand2_2 _30311_ (.A(_08279_),
    .B(_08281_),
    .Y(_08285_));
 sky130_fd_sc_hd__nand3_2 _30312_ (.A(_08269_),
    .B(_08274_),
    .C(_08285_),
    .Y(_08286_));
 sky130_fd_sc_hd__nand3_2 _30313_ (.A(_08283_),
    .B(_08284_),
    .C(_08286_),
    .Y(_08287_));
 sky130_fd_sc_hd__nand2_2 _30314_ (.A(_08275_),
    .B(_08285_),
    .Y(_08288_));
 sky130_fd_sc_hd__o21ai_2 _30315_ (.A1(_08012_),
    .A2(_08002_),
    .B1(_08017_),
    .Y(_08289_));
 sky130_fd_sc_hd__nand3_2 _30316_ (.A(_08269_),
    .B(_08274_),
    .C(_08282_),
    .Y(_08290_));
 sky130_fd_sc_hd__nand3_2 _30317_ (.A(_08288_),
    .B(_08289_),
    .C(_08290_),
    .Y(_08291_));
 sky130_fd_sc_hd__nand2_2 _30318_ (.A(_08287_),
    .B(_08291_),
    .Y(_08292_));
 sky130_fd_sc_hd__nor2_2 _30319_ (.A(_08010_),
    .B(_08292_),
    .Y(_08293_));
 sky130_fd_sc_hd__nand2_2 _30320_ (.A(_08292_),
    .B(_08010_),
    .Y(_08294_));
 sky130_fd_sc_hd__o21ai_2 _30321_ (.A1(_07758_),
    .A2(_08033_),
    .B1(_08027_),
    .Y(_08295_));
 sky130_fd_sc_hd__nand2_2 _30322_ (.A(_08294_),
    .B(_08295_),
    .Y(_08296_));
 sky130_fd_sc_hd__nand3_2 _30323_ (.A(_08287_),
    .B(_08291_),
    .C(_08010_),
    .Y(_08297_));
 sky130_fd_sc_hd__inv_2 _30324_ (.A(_08010_),
    .Y(_08298_));
 sky130_fd_sc_hd__nand2_2 _30325_ (.A(_08292_),
    .B(_08298_),
    .Y(_08299_));
 sky130_fd_sc_hd__o2111ai_2 _30326_ (.A1(_07758_),
    .A2(_08033_),
    .B1(_08027_),
    .C1(_08297_),
    .D1(_08299_),
    .Y(_08300_));
 sky130_fd_sc_hd__o21a_2 _30327_ (.A1(_08293_),
    .A2(_08296_),
    .B1(_08300_),
    .X(_08301_));
 sky130_fd_sc_hd__nand3_2 _30328_ (.A(_08035_),
    .B(_08028_),
    .C(_08031_),
    .Y(_08302_));
 sky130_fd_sc_hd__o21ai_2 _30329_ (.A1(_08036_),
    .A2(_08043_),
    .B1(_08302_),
    .Y(_08303_));
 sky130_fd_sc_hd__xor2_2 _30330_ (.A(_08301_),
    .B(_08303_),
    .X(_02642_));
 sky130_fd_sc_hd__nand3_2 _30331_ (.A(_08140_),
    .B(_08259_),
    .C(_08143_),
    .Y(_08304_));
 sky130_fd_sc_hd__nand2_2 _30332_ (.A(_08304_),
    .B(_08261_),
    .Y(_08305_));
 sky130_fd_sc_hd__nor3_2 _30333_ (.A(_08253_),
    .B(_08247_),
    .C(_08249_),
    .Y(_08306_));
 sky130_fd_sc_hd__nand2_2 _30334_ (.A(_06624_),
    .B(_06497_),
    .Y(_08307_));
 sky130_fd_sc_hd__nand2_2 _30335_ (.A(_07015_),
    .B(_06539_),
    .Y(_08308_));
 sky130_fd_sc_hd__nor2_2 _30336_ (.A(_08307_),
    .B(_08308_),
    .Y(_08309_));
 sky130_fd_sc_hd__nand2_2 _30337_ (.A(_06117_),
    .B(_05896_),
    .Y(_08310_));
 sky130_fd_sc_hd__inv_2 _30338_ (.A(_08310_),
    .Y(_08311_));
 sky130_fd_sc_hd__nand2_2 _30339_ (.A(_08307_),
    .B(_08308_),
    .Y(_08312_));
 sky130_fd_sc_hd__nand2_2 _30340_ (.A(_08311_),
    .B(_08312_),
    .Y(_08313_));
 sky130_fd_sc_hd__o21ai_2 _30341_ (.A1(_08203_),
    .A2(_08204_),
    .B1(_08206_),
    .Y(_08314_));
 sky130_fd_sc_hd__buf_1 _30342_ (.A(_19362_),
    .X(_08315_));
 sky130_fd_sc_hd__a22oi_2 _30343_ (.A1(_08315_),
    .A2(_19609_),
    .B1(_07934_),
    .B2(_06540_),
    .Y(_08316_));
 sky130_fd_sc_hd__o21ai_2 _30344_ (.A1(_08316_),
    .A2(_08309_),
    .B1(_08310_),
    .Y(_08317_));
 sky130_fd_sc_hd__o2111ai_2 _30345_ (.A1(_08309_),
    .A2(_08313_),
    .B1(_08209_),
    .C1(_08314_),
    .D1(_08317_),
    .Y(_08318_));
 sky130_fd_sc_hd__o21ai_2 _30346_ (.A1(_08316_),
    .A2(_08309_),
    .B1(_08311_),
    .Y(_08319_));
 sky130_fd_sc_hd__buf_1 _30347_ (.A(_06272_),
    .X(_08320_));
 sky130_fd_sc_hd__nand3b_2 _30348_ (.A_N(_08307_),
    .B(_08320_),
    .C(_05911_),
    .Y(_08321_));
 sky130_fd_sc_hd__nand3_2 _30349_ (.A(_08321_),
    .B(_08312_),
    .C(_08310_),
    .Y(_08322_));
 sky130_fd_sc_hd__nand2_2 _30350_ (.A(_08314_),
    .B(_08209_),
    .Y(_08323_));
 sky130_fd_sc_hd__nand3_2 _30351_ (.A(_08319_),
    .B(_08322_),
    .C(_08323_),
    .Y(_08324_));
 sky130_fd_sc_hd__a22oi_2 _30352_ (.A1(_06500_),
    .A2(_06724_),
    .B1(_06433_),
    .B2(_07143_),
    .Y(_08325_));
 sky130_fd_sc_hd__nand2_2 _30353_ (.A(_06430_),
    .B(_08218_),
    .Y(_08326_));
 sky130_fd_sc_hd__nand2_2 _30354_ (.A(_06258_),
    .B(_06206_),
    .Y(_08327_));
 sky130_fd_sc_hd__nor2_2 _30355_ (.A(_08326_),
    .B(_08327_),
    .Y(_08328_));
 sky130_fd_sc_hd__nand2_2 _30356_ (.A(_06616_),
    .B(_19594_),
    .Y(_08329_));
 sky130_fd_sc_hd__o21bai_2 _30357_ (.A1(_08325_),
    .A2(_08328_),
    .B1_N(_08329_),
    .Y(_08330_));
 sky130_fd_sc_hd__buf_1 _30358_ (.A(_05958_),
    .X(_08331_));
 sky130_fd_sc_hd__nand3b_2 _30359_ (.A_N(_08326_),
    .B(_08331_),
    .C(_19597_),
    .Y(_08332_));
 sky130_fd_sc_hd__nand2_2 _30360_ (.A(_08326_),
    .B(_08327_),
    .Y(_08333_));
 sky130_fd_sc_hd__nand3_2 _30361_ (.A(_08332_),
    .B(_08333_),
    .C(_08329_),
    .Y(_08334_));
 sky130_fd_sc_hd__nand2_2 _30362_ (.A(_08330_),
    .B(_08334_),
    .Y(_08335_));
 sky130_fd_sc_hd__and3_2 _30363_ (.A(_08318_),
    .B(_08324_),
    .C(_08335_),
    .X(_08336_));
 sky130_fd_sc_hd__a21oi_2 _30364_ (.A1(_08318_),
    .A2(_08324_),
    .B1(_08335_),
    .Y(_08337_));
 sky130_fd_sc_hd__nand2_2 _30365_ (.A(_08188_),
    .B(_08197_),
    .Y(_08338_));
 sky130_fd_sc_hd__a22oi_2 _30366_ (.A1(_07886_),
    .A2(_05505_),
    .B1(_06828_),
    .B2(_05613_),
    .Y(_08339_));
 sky130_fd_sc_hd__nand3_2 _30367_ (.A(_07416_),
    .B(_07417_),
    .C(_06808_),
    .Y(_08340_));
 sky130_fd_sc_hd__nor2_2 _30368_ (.A(_05731_),
    .B(_08340_),
    .Y(_08341_));
 sky130_fd_sc_hd__and2_2 _30369_ (.A(_07890_),
    .B(_19613_),
    .X(_08342_));
 sky130_fd_sc_hd__o21bai_2 _30370_ (.A1(_08339_),
    .A2(_08341_),
    .B1_N(_08342_),
    .Y(_08343_));
 sky130_fd_sc_hd__o22ai_2 _30371_ (.A1(_05850_),
    .A2(_08161_),
    .B1(_08164_),
    .B2(_08160_),
    .Y(_08344_));
 sky130_fd_sc_hd__buf_1 _30372_ (.A(_06823_),
    .X(_08345_));
 sky130_fd_sc_hd__a22o_2 _30373_ (.A1(_07898_),
    .A2(_19619_),
    .B1(_08345_),
    .B2(_19616_),
    .X(_08346_));
 sky130_fd_sc_hd__o211ai_2 _30374_ (.A1(_05732_),
    .A2(_08340_),
    .B1(_08342_),
    .C1(_08346_),
    .Y(_08347_));
 sky130_fd_sc_hd__nand3_2 _30375_ (.A(_08343_),
    .B(_08344_),
    .C(_08347_),
    .Y(_08348_));
 sky130_fd_sc_hd__o21ai_2 _30376_ (.A1(_08339_),
    .A2(_08341_),
    .B1(_08342_),
    .Y(_08349_));
 sky130_fd_sc_hd__a22o_2 _30377_ (.A1(_19347_),
    .A2(_05330_),
    .B1(_08159_),
    .B2(_06501_),
    .X(_08350_));
 sky130_fd_sc_hd__a2bb2oi_2 _30378_ (.A1_N(_05850_),
    .A2_N(_08161_),
    .B1(_08165_),
    .B2(_08350_),
    .Y(_08351_));
 sky130_fd_sc_hd__buf_1 _30379_ (.A(_06831_),
    .X(_08352_));
 sky130_fd_sc_hd__o221ai_2 _30380_ (.A1(_08352_),
    .A2(_06505_),
    .B1(_05732_),
    .B2(_08340_),
    .C1(_08346_),
    .Y(_08353_));
 sky130_fd_sc_hd__nand3_2 _30381_ (.A(_08349_),
    .B(_08351_),
    .C(_08353_),
    .Y(_08354_));
 sky130_fd_sc_hd__nor2_2 _30382_ (.A(_08181_),
    .B(_08178_),
    .Y(_08355_));
 sky130_fd_sc_hd__o2bb2ai_2 _30383_ (.A1_N(_08348_),
    .A2_N(_08354_),
    .B1(_08176_),
    .B2(_08355_),
    .Y(_08356_));
 sky130_fd_sc_hd__nor2_2 _30384_ (.A(_08176_),
    .B(_08355_),
    .Y(_08357_));
 sky130_fd_sc_hd__nand3_2 _30385_ (.A(_08354_),
    .B(_08348_),
    .C(_08357_),
    .Y(_08358_));
 sky130_fd_sc_hd__a22oi_2 _30386_ (.A1(_08194_),
    .A2(_08338_),
    .B1(_08356_),
    .B2(_08358_),
    .Y(_08359_));
 sky130_fd_sc_hd__and3_2 _30387_ (.A(_08180_),
    .B(_08187_),
    .C(_08184_),
    .X(_08360_));
 sky130_fd_sc_hd__a31oi_2 _30388_ (.A1(_08189_),
    .A2(_08192_),
    .A3(_08193_),
    .B1(_08197_),
    .Y(_08361_));
 sky130_fd_sc_hd__o211a_2 _30389_ (.A1(_08360_),
    .A2(_08361_),
    .B1(_08358_),
    .C1(_08356_),
    .X(_08362_));
 sky130_fd_sc_hd__o22ai_2 _30390_ (.A1(_08336_),
    .A2(_08337_),
    .B1(_08359_),
    .B2(_08362_),
    .Y(_08363_));
 sky130_fd_sc_hd__nor2_2 _30391_ (.A(_08337_),
    .B(_08336_),
    .Y(_08364_));
 sky130_fd_sc_hd__inv_2 _30392_ (.A(_08194_),
    .Y(_08365_));
 sky130_fd_sc_hd__and2_2 _30393_ (.A(_08188_),
    .B(_08197_),
    .X(_08366_));
 sky130_fd_sc_hd__o2bb2ai_2 _30394_ (.A1_N(_08358_),
    .A2_N(_08356_),
    .B1(_08365_),
    .B2(_08366_),
    .Y(_08367_));
 sky130_fd_sc_hd__o211ai_2 _30395_ (.A1(_08361_),
    .A2(_08360_),
    .B1(_08358_),
    .C1(_08356_),
    .Y(_08368_));
 sky130_fd_sc_hd__nand3_2 _30396_ (.A(_08364_),
    .B(_08367_),
    .C(_08368_),
    .Y(_08369_));
 sky130_fd_sc_hd__nand3_2 _30397_ (.A(_08363_),
    .B(_08369_),
    .C(_08171_),
    .Y(_08370_));
 sky130_fd_sc_hd__o21ai_2 _30398_ (.A1(_08359_),
    .A2(_08362_),
    .B1(_08364_),
    .Y(_08371_));
 sky130_fd_sc_hd__nand3_2 _30399_ (.A(_08172_),
    .B(_08168_),
    .C(_08169_),
    .Y(_08372_));
 sky130_fd_sc_hd__and2_2 _30400_ (.A(_08324_),
    .B(_08335_),
    .X(_08373_));
 sky130_fd_sc_hd__a21o_2 _30401_ (.A1(_08373_),
    .A2(_08318_),
    .B1(_08337_),
    .X(_08374_));
 sky130_fd_sc_hd__nand3_2 _30402_ (.A(_08374_),
    .B(_08367_),
    .C(_08368_),
    .Y(_08375_));
 sky130_fd_sc_hd__nand3_2 _30403_ (.A(_08371_),
    .B(_08372_),
    .C(_08375_),
    .Y(_08376_));
 sky130_fd_sc_hd__nor2_2 _30404_ (.A(_08201_),
    .B(_08237_),
    .Y(_08377_));
 sky130_fd_sc_hd__o2bb2ai_2 _30405_ (.A1_N(_08370_),
    .A2_N(_08376_),
    .B1(_08199_),
    .B2(_08377_),
    .Y(_08378_));
 sky130_fd_sc_hd__o21ai_2 _30406_ (.A1(_08199_),
    .A2(_08231_),
    .B1(_08238_),
    .Y(_08379_));
 sky130_fd_sc_hd__nand3_2 _30407_ (.A(_08376_),
    .B(_08370_),
    .C(_08379_),
    .Y(_08380_));
 sky130_fd_sc_hd__a21oi_2 _30408_ (.A1(_08152_),
    .A2(_08153_),
    .B1(_08147_),
    .Y(_08381_));
 sky130_fd_sc_hd__buf_1 _30409_ (.A(\pcpi_mul.rs2[23] ),
    .X(_08382_));
 sky130_fd_sc_hd__buf_1 _30410_ (.A(_19339_),
    .X(_08383_));
 sky130_fd_sc_hd__a22oi_2 _30411_ (.A1(_08382_),
    .A2(_05804_),
    .B1(_08383_),
    .B2(_19633_),
    .Y(_08384_));
 sky130_fd_sc_hd__buf_1 _30412_ (.A(\pcpi_mul.rs2[23] ),
    .X(_08385_));
 sky130_fd_sc_hd__buf_1 _30413_ (.A(\pcpi_mul.rs2[22] ),
    .X(_08386_));
 sky130_fd_sc_hd__and4_2 _30414_ (.A(_08385_),
    .B(_08386_),
    .C(_05545_),
    .D(_07904_),
    .X(_08387_));
 sky130_fd_sc_hd__buf_1 _30415_ (.A(\pcpi_mul.rs2[21] ),
    .X(_08388_));
 sky130_fd_sc_hd__nand2_2 _30416_ (.A(_08388_),
    .B(_06792_),
    .Y(_08389_));
 sky130_fd_sc_hd__o21ai_2 _30417_ (.A1(_08384_),
    .A2(_08387_),
    .B1(_08389_),
    .Y(_08390_));
 sky130_fd_sc_hd__buf_1 _30418_ (.A(\pcpi_mul.rs2[23] ),
    .X(_08391_));
 sky130_fd_sc_hd__nand2_2 _30419_ (.A(_08391_),
    .B(_05543_),
    .Y(_08392_));
 sky130_fd_sc_hd__buf_1 _30420_ (.A(_05323_),
    .X(_08393_));
 sky130_fd_sc_hd__nand3b_2 _30421_ (.A_N(_08392_),
    .B(_19340_),
    .C(_08393_),
    .Y(_08394_));
 sky130_fd_sc_hd__inv_2 _30422_ (.A(_08389_),
    .Y(_08395_));
 sky130_fd_sc_hd__buf_1 _30423_ (.A(\pcpi_mul.rs2[23] ),
    .X(_08396_));
 sky130_fd_sc_hd__a22o_2 _30424_ (.A1(_08396_),
    .A2(_19636_),
    .B1(_08383_),
    .B2(_19633_),
    .X(_08397_));
 sky130_fd_sc_hd__nand3_2 _30425_ (.A(_08394_),
    .B(_08395_),
    .C(_08397_),
    .Y(_08398_));
 sky130_fd_sc_hd__nand3b_2 _30426_ (.A_N(_08381_),
    .B(_08390_),
    .C(_08398_),
    .Y(_08399_));
 sky130_fd_sc_hd__o21ai_2 _30427_ (.A1(_08384_),
    .A2(_08387_),
    .B1(_08395_),
    .Y(_08400_));
 sky130_fd_sc_hd__nand3_2 _30428_ (.A(_08394_),
    .B(_08389_),
    .C(_08397_),
    .Y(_08401_));
 sky130_fd_sc_hd__nand3_2 _30429_ (.A(_08400_),
    .B(_08401_),
    .C(_08381_),
    .Y(_08402_));
 sky130_fd_sc_hd__a22oi_2 _30430_ (.A1(_07894_),
    .A2(_05338_),
    .B1(_08159_),
    .B2(_05765_),
    .Y(_08403_));
 sky130_fd_sc_hd__nand2_2 _30431_ (.A(_19346_),
    .B(_05158_),
    .Y(_08404_));
 sky130_fd_sc_hd__nand2_2 _30432_ (.A(_19349_),
    .B(_05340_),
    .Y(_08405_));
 sky130_fd_sc_hd__nor2_2 _30433_ (.A(_08404_),
    .B(_08405_),
    .Y(_08406_));
 sky130_fd_sc_hd__buf_1 _30434_ (.A(\pcpi_mul.rs2[18] ),
    .X(_08407_));
 sky130_fd_sc_hd__nand2_2 _30435_ (.A(_08407_),
    .B(_06614_),
    .Y(_08408_));
 sky130_fd_sc_hd__o21bai_2 _30436_ (.A1(_08403_),
    .A2(_08406_),
    .B1_N(_08408_),
    .Y(_08409_));
 sky130_fd_sc_hd__nand3b_2 _30437_ (.A_N(_08404_),
    .B(_19350_),
    .C(_05341_),
    .Y(_08410_));
 sky130_fd_sc_hd__nand2_2 _30438_ (.A(_08404_),
    .B(_08405_),
    .Y(_08411_));
 sky130_fd_sc_hd__nand3_2 _30439_ (.A(_08410_),
    .B(_08411_),
    .C(_08408_),
    .Y(_08412_));
 sky130_fd_sc_hd__nand2_2 _30440_ (.A(_08409_),
    .B(_08412_),
    .Y(_08413_));
 sky130_fd_sc_hd__a21o_2 _30441_ (.A1(_08399_),
    .A2(_08402_),
    .B1(_08413_),
    .X(_08414_));
 sky130_fd_sc_hd__nand3_2 _30442_ (.A(_08399_),
    .B(_08402_),
    .C(_08413_),
    .Y(_08415_));
 sky130_fd_sc_hd__nand2_2 _30443_ (.A(_08414_),
    .B(_08415_),
    .Y(_08416_));
 sky130_fd_sc_hd__nand2_2 _30444_ (.A(_08167_),
    .B(_08158_),
    .Y(_08417_));
 sky130_fd_sc_hd__and2_2 _30445_ (.A(_08417_),
    .B(_08155_),
    .X(_08418_));
 sky130_fd_sc_hd__nand2_2 _30446_ (.A(_08416_),
    .B(_08418_),
    .Y(_08419_));
 sky130_fd_sc_hd__nand2_2 _30447_ (.A(_08417_),
    .B(_08155_),
    .Y(_08420_));
 sky130_fd_sc_hd__nand3_2 _30448_ (.A(_08420_),
    .B(_08414_),
    .C(_08415_),
    .Y(_08421_));
 sky130_fd_sc_hd__buf_1 _30449_ (.A(_08421_),
    .X(_08422_));
 sky130_fd_sc_hd__inv_2 _30450_ (.A(\pcpi_mul.rs2[24] ),
    .Y(_08423_));
 sky130_fd_sc_hd__buf_1 _30451_ (.A(_08423_),
    .X(_08424_));
 sky130_fd_sc_hd__nor2_2 _30452_ (.A(_08424_),
    .B(_04839_),
    .Y(_08425_));
 sky130_fd_sc_hd__a21oi_2 _30453_ (.A1(_08419_),
    .A2(_08422_),
    .B1(_08425_),
    .Y(_08426_));
 sky130_fd_sc_hd__inv_2 _30454_ (.A(_08425_),
    .Y(_08427_));
 sky130_fd_sc_hd__a21oi_2 _30455_ (.A1(_08414_),
    .A2(_08415_),
    .B1(_08420_),
    .Y(_08428_));
 sky130_fd_sc_hd__nor3b_2 _30456_ (.A(_08427_),
    .B(_08428_),
    .C_N(_08422_),
    .Y(_08429_));
 sky130_fd_sc_hd__nor2_2 _30457_ (.A(_08426_),
    .B(_08429_),
    .Y(_08430_));
 sky130_fd_sc_hd__nand3_2 _30458_ (.A(_08378_),
    .B(_08380_),
    .C(_08430_),
    .Y(_08431_));
 sky130_fd_sc_hd__o2bb2ai_2 _30459_ (.A1_N(_08380_),
    .A2_N(_08378_),
    .B1(_08426_),
    .B2(_08429_),
    .Y(_08432_));
 sky130_fd_sc_hd__nand3_2 _30460_ (.A(_08306_),
    .B(_08431_),
    .C(_08432_),
    .Y(_08433_));
 sky130_fd_sc_hd__inv_2 _30461_ (.A(_08426_),
    .Y(_08434_));
 sky130_fd_sc_hd__nand3_2 _30462_ (.A(_08419_),
    .B(_08425_),
    .C(_08422_),
    .Y(_08435_));
 sky130_fd_sc_hd__a22oi_2 _30463_ (.A1(_08434_),
    .A2(_08435_),
    .B1(_08378_),
    .B2(_08380_),
    .Y(_08436_));
 sky130_fd_sc_hd__and3_2 _30464_ (.A(_08363_),
    .B(_08171_),
    .C(_08369_),
    .X(_08437_));
 sky130_fd_sc_hd__nand2_2 _30465_ (.A(_08376_),
    .B(_08379_),
    .Y(_08438_));
 sky130_fd_sc_hd__o211a_2 _30466_ (.A1(_08437_),
    .A2(_08438_),
    .B1(_08430_),
    .C1(_08378_),
    .X(_08439_));
 sky130_fd_sc_hd__o22ai_2 _30467_ (.A1(_08249_),
    .A2(_08264_),
    .B1(_08436_),
    .B2(_08439_),
    .Y(_08440_));
 sky130_fd_sc_hd__buf_1 _30468_ (.A(_08440_),
    .X(_08441_));
 sky130_fd_sc_hd__a22oi_2 _30469_ (.A1(_05542_),
    .A2(_06949_),
    .B1(_05445_),
    .B2(_06951_),
    .Y(_08442_));
 sky130_fd_sc_hd__and4_2 _30470_ (.A(_05758_),
    .B(_05641_),
    .C(_19587_),
    .D(_06949_),
    .X(_08443_));
 sky130_fd_sc_hd__nand2_2 _30471_ (.A(_05763_),
    .B(_19584_),
    .Y(_08444_));
 sky130_fd_sc_hd__o21ai_2 _30472_ (.A1(_08442_),
    .A2(_08443_),
    .B1(_08444_),
    .Y(_08445_));
 sky130_fd_sc_hd__nand2_2 _30473_ (.A(_05639_),
    .B(_07360_),
    .Y(_08446_));
 sky130_fd_sc_hd__buf_1 _30474_ (.A(_19587_),
    .X(_08447_));
 sky130_fd_sc_hd__nand3b_2 _30475_ (.A_N(_08446_),
    .B(_06896_),
    .C(_08447_),
    .Y(_08448_));
 sky130_fd_sc_hd__inv_2 _30476_ (.A(_08444_),
    .Y(_08449_));
 sky130_fd_sc_hd__a22o_2 _30477_ (.A1(_05542_),
    .A2(_06542_),
    .B1(_19383_),
    .B2(_06951_),
    .X(_08450_));
 sky130_fd_sc_hd__nand3_2 _30478_ (.A(_08448_),
    .B(_08449_),
    .C(_08450_),
    .Y(_08451_));
 sky130_fd_sc_hd__o21ai_2 _30479_ (.A1(_08221_),
    .A2(_08216_),
    .B1(_08224_),
    .Y(_08452_));
 sky130_fd_sc_hd__and3_2 _30480_ (.A(_08445_),
    .B(_08451_),
    .C(_08452_),
    .X(_08453_));
 sky130_fd_sc_hd__o21ai_2 _30481_ (.A1(_08442_),
    .A2(_08443_),
    .B1(_08449_),
    .Y(_08454_));
 sky130_fd_sc_hd__nand3_2 _30482_ (.A(_08448_),
    .B(_08444_),
    .C(_08450_),
    .Y(_08455_));
 sky130_fd_sc_hd__a21oi_2 _30483_ (.A1(_08222_),
    .A2(_08225_),
    .B1(_08220_),
    .Y(_08456_));
 sky130_fd_sc_hd__nand3_2 _30484_ (.A(_08454_),
    .B(_08455_),
    .C(_08456_),
    .Y(_08457_));
 sky130_fd_sc_hd__nor2_2 _30485_ (.A(_08049_),
    .B(_08047_),
    .Y(_08458_));
 sky130_fd_sc_hd__nor2_2 _30486_ (.A(_08044_),
    .B(_08458_),
    .Y(_08459_));
 sky130_fd_sc_hd__nand2_2 _30487_ (.A(_08457_),
    .B(_08459_),
    .Y(_08460_));
 sky130_fd_sc_hd__nand3_2 _30488_ (.A(_08445_),
    .B(_08451_),
    .C(_08452_),
    .Y(_08461_));
 sky130_fd_sc_hd__o2bb2ai_2 _30489_ (.A1_N(_08461_),
    .A2_N(_08457_),
    .B1(_08044_),
    .B2(_08458_),
    .Y(_08462_));
 sky130_fd_sc_hd__nand2_2 _30490_ (.A(_08214_),
    .B(_08227_),
    .Y(_08463_));
 sky130_fd_sc_hd__nand2_2 _30491_ (.A(_08463_),
    .B(_08213_),
    .Y(_08464_));
 sky130_fd_sc_hd__o211a_2 _30492_ (.A1(_08453_),
    .A2(_08460_),
    .B1(_08462_),
    .C1(_08464_),
    .X(_08465_));
 sky130_fd_sc_hd__a21oi_2 _30493_ (.A1(_08461_),
    .A2(_08457_),
    .B1(_08459_),
    .Y(_08466_));
 sky130_fd_sc_hd__nor2_2 _30494_ (.A(_08048_),
    .B(_08044_),
    .Y(_08467_));
 sky130_fd_sc_hd__o211a_2 _30495_ (.A1(_08047_),
    .A2(_08467_),
    .B1(_08461_),
    .C1(_08457_),
    .X(_08468_));
 sky130_fd_sc_hd__o21bai_2 _30496_ (.A1(_08466_),
    .A2(_08468_),
    .B1_N(_08464_),
    .Y(_08469_));
 sky130_fd_sc_hd__nand2_2 _30497_ (.A(_08069_),
    .B(_08060_),
    .Y(_08470_));
 sky130_fd_sc_hd__nand2_2 _30498_ (.A(_08469_),
    .B(_08470_),
    .Y(_08471_));
 sky130_fd_sc_hd__o21ai_2 _30499_ (.A1(_08072_),
    .A2(_08067_),
    .B1(_08077_),
    .Y(_08472_));
 sky130_fd_sc_hd__nand3_2 _30500_ (.A(_08461_),
    .B(_08457_),
    .C(_08459_),
    .Y(_08473_));
 sky130_fd_sc_hd__a21oi_2 _30501_ (.A1(_08462_),
    .A2(_08473_),
    .B1(_08464_),
    .Y(_08474_));
 sky130_fd_sc_hd__inv_2 _30502_ (.A(_08470_),
    .Y(_08475_));
 sky130_fd_sc_hd__o21ai_2 _30503_ (.A1(_08474_),
    .A2(_08465_),
    .B1(_08475_),
    .Y(_08476_));
 sky130_fd_sc_hd__o211ai_2 _30504_ (.A1(_08465_),
    .A2(_08471_),
    .B1(_08472_),
    .C1(_08476_),
    .Y(_08477_));
 sky130_fd_sc_hd__o21ai_2 _30505_ (.A1(_08474_),
    .A2(_08465_),
    .B1(_08470_),
    .Y(_08478_));
 sky130_fd_sc_hd__nand2_2 _30506_ (.A(_08077_),
    .B(_08072_),
    .Y(_08479_));
 sky130_fd_sc_hd__nand2_2 _30507_ (.A(_08479_),
    .B(_08076_),
    .Y(_08480_));
 sky130_fd_sc_hd__nand3_2 _30508_ (.A(_08464_),
    .B(_08462_),
    .C(_08473_),
    .Y(_08481_));
 sky130_fd_sc_hd__nand3_2 _30509_ (.A(_08469_),
    .B(_08475_),
    .C(_08481_),
    .Y(_08482_));
 sky130_fd_sc_hd__nand3_2 _30510_ (.A(_08478_),
    .B(_08480_),
    .C(_08482_),
    .Y(_08483_));
 sky130_fd_sc_hd__nand2_2 _30511_ (.A(_08477_),
    .B(_08483_),
    .Y(_08484_));
 sky130_fd_sc_hd__and4_2 _30512_ (.A(_06731_),
    .B(_05891_),
    .C(_07358_),
    .D(_07377_),
    .X(_08485_));
 sky130_fd_sc_hd__a22o_2 _30513_ (.A1(_06199_),
    .A2(_07593_),
    .B1(_19391_),
    .B2(_07590_),
    .X(_08486_));
 sky130_fd_sc_hd__inv_2 _30514_ (.A(\pcpi_mul.rs1[24] ),
    .Y(_08487_));
 sky130_fd_sc_hd__nor2_2 _30515_ (.A(_04835_),
    .B(_08487_),
    .Y(_08488_));
 sky130_fd_sc_hd__nand3b_2 _30516_ (.A_N(_08485_),
    .B(_08486_),
    .C(_08488_),
    .Y(_08489_));
 sky130_fd_sc_hd__buf_1 _30517_ (.A(_07377_),
    .X(_08490_));
 sky130_fd_sc_hd__a22oi_2 _30518_ (.A1(_05712_),
    .A2(_08490_),
    .B1(_05892_),
    .B2(_08108_),
    .Y(_08491_));
 sky130_fd_sc_hd__o21bai_2 _30519_ (.A1(_08491_),
    .A2(_08485_),
    .B1_N(_08488_),
    .Y(_08492_));
 sky130_fd_sc_hd__o21ai_2 _30520_ (.A1(_08086_),
    .A2(_08087_),
    .B1(_08092_),
    .Y(_08493_));
 sky130_fd_sc_hd__a21oi_2 _30521_ (.A1(_08489_),
    .A2(_08492_),
    .B1(_08493_),
    .Y(_08494_));
 sky130_fd_sc_hd__o211a_2 _30522_ (.A1(_08095_),
    .A2(_08088_),
    .B1(_08492_),
    .C1(_08489_),
    .X(_08495_));
 sky130_fd_sc_hd__buf_1 _30523_ (.A(_08085_),
    .X(_08496_));
 sky130_fd_sc_hd__buf_1 _30524_ (.A(\pcpi_mul.rs1[22] ),
    .X(_08497_));
 sky130_fd_sc_hd__nand2_2 _30525_ (.A(_05203_),
    .B(_08497_),
    .Y(_08498_));
 sky130_fd_sc_hd__a21o_2 _30526_ (.A1(_05909_),
    .A2(_08496_),
    .B1(_08498_),
    .X(_08499_));
 sky130_fd_sc_hd__nand2_2 _30527_ (.A(_05143_),
    .B(_19570_),
    .Y(_08500_));
 sky130_fd_sc_hd__a21o_2 _30528_ (.A1(_05736_),
    .A2(_19574_),
    .B1(_08500_),
    .X(_08501_));
 sky130_fd_sc_hd__nand2_2 _30529_ (.A(_05115_),
    .B(_07845_),
    .Y(_08502_));
 sky130_fd_sc_hd__a21o_2 _30530_ (.A1(_08499_),
    .A2(_08501_),
    .B1(_08502_),
    .X(_08503_));
 sky130_fd_sc_hd__nand3_2 _30531_ (.A(_08499_),
    .B(_08501_),
    .C(_08502_),
    .Y(_08504_));
 sky130_fd_sc_hd__nand2_2 _30532_ (.A(_08503_),
    .B(_08504_),
    .Y(_08505_));
 sky130_fd_sc_hd__o21ai_2 _30533_ (.A1(_08494_),
    .A2(_08495_),
    .B1(_08505_),
    .Y(_08506_));
 sky130_fd_sc_hd__nand2_2 _30534_ (.A(_08128_),
    .B(_08097_),
    .Y(_08507_));
 sky130_fd_sc_hd__and2_2 _30535_ (.A(_08503_),
    .B(_08504_),
    .X(_08508_));
 sky130_fd_sc_hd__nand2_2 _30536_ (.A(_08489_),
    .B(_08492_),
    .Y(_08509_));
 sky130_fd_sc_hd__nor2_2 _30537_ (.A(_08095_),
    .B(_08088_),
    .Y(_08510_));
 sky130_fd_sc_hd__nand2_2 _30538_ (.A(_08509_),
    .B(_08510_),
    .Y(_08511_));
 sky130_fd_sc_hd__nand3_2 _30539_ (.A(_08489_),
    .B(_08493_),
    .C(_08492_),
    .Y(_08512_));
 sky130_fd_sc_hd__nand3_2 _30540_ (.A(_08508_),
    .B(_08511_),
    .C(_08512_),
    .Y(_08513_));
 sky130_fd_sc_hd__nand3_2 _30541_ (.A(_08506_),
    .B(_08507_),
    .C(_08513_),
    .Y(_08514_));
 sky130_fd_sc_hd__a21oi_2 _30542_ (.A1(_08113_),
    .A2(_08102_),
    .B1(_08126_),
    .Y(_08515_));
 sky130_fd_sc_hd__o21ai_2 _30543_ (.A1(_08494_),
    .A2(_08495_),
    .B1(_08508_),
    .Y(_08516_));
 sky130_fd_sc_hd__nand3_2 _30544_ (.A(_08511_),
    .B(_08505_),
    .C(_08512_),
    .Y(_08517_));
 sky130_fd_sc_hd__nor2_2 _30545_ (.A(_08104_),
    .B(_08106_),
    .Y(_08518_));
 sky130_fd_sc_hd__nor2_2 _30546_ (.A(_08518_),
    .B(_08111_),
    .Y(_08519_));
 sky130_fd_sc_hd__a31oi_2 _30547_ (.A1(_08515_),
    .A2(_08516_),
    .A3(_08517_),
    .B1(_08519_),
    .Y(_08520_));
 sky130_fd_sc_hd__nand3_2 _30548_ (.A(_08515_),
    .B(_08516_),
    .C(_08517_),
    .Y(_08521_));
 sky130_fd_sc_hd__inv_2 _30549_ (.A(_08519_),
    .Y(_08522_));
 sky130_fd_sc_hd__a21oi_2 _30550_ (.A1(_08521_),
    .A2(_08514_),
    .B1(_08522_),
    .Y(_08523_));
 sky130_fd_sc_hd__a21oi_2 _30551_ (.A1(_08514_),
    .A2(_08520_),
    .B1(_08523_),
    .Y(_08524_));
 sky130_fd_sc_hd__nand2_2 _30552_ (.A(_08484_),
    .B(_08524_),
    .Y(_08525_));
 sky130_fd_sc_hd__a21boi_2 _30553_ (.A1(_08245_),
    .A2(_08246_),
    .B1_N(_08240_),
    .Y(_08526_));
 sky130_fd_sc_hd__and3_2 _30554_ (.A(_08521_),
    .B(_08514_),
    .C(_08522_),
    .X(_08527_));
 sky130_fd_sc_hd__o211ai_2 _30555_ (.A1(_08523_),
    .A2(_08527_),
    .B1(_08483_),
    .C1(_08477_),
    .Y(_08528_));
 sky130_fd_sc_hd__nand3_2 _30556_ (.A(_08525_),
    .B(_08526_),
    .C(_08528_),
    .Y(_08529_));
 sky130_fd_sc_hd__o2bb2ai_2 _30557_ (.A1_N(_08483_),
    .A2_N(_08477_),
    .B1(_08527_),
    .B2(_08523_),
    .Y(_08530_));
 sky130_fd_sc_hd__nand3_2 _30558_ (.A(_08524_),
    .B(_08483_),
    .C(_08477_),
    .Y(_08531_));
 sky130_fd_sc_hd__nand2_2 _30559_ (.A(_08245_),
    .B(_08246_),
    .Y(_08532_));
 sky130_fd_sc_hd__nand2_2 _30560_ (.A(_08532_),
    .B(_08240_),
    .Y(_08533_));
 sky130_fd_sc_hd__nand3_2 _30561_ (.A(_08530_),
    .B(_08531_),
    .C(_08533_),
    .Y(_08534_));
 sky130_fd_sc_hd__nand2_2 _30562_ (.A(_08137_),
    .B(_08084_),
    .Y(_08535_));
 sky130_fd_sc_hd__a21oi_2 _30563_ (.A1(_08529_),
    .A2(_08534_),
    .B1(_08535_),
    .Y(_08536_));
 sky130_fd_sc_hd__and3_2 _30564_ (.A(_08529_),
    .B(_08534_),
    .C(_08535_),
    .X(_08537_));
 sky130_fd_sc_hd__o2bb2ai_2 _30565_ (.A1_N(_08433_),
    .A2_N(_08441_),
    .B1(_08536_),
    .B2(_08537_),
    .Y(_08538_));
 sky130_fd_sc_hd__a21oi_2 _30566_ (.A1(_08525_),
    .A2(_08528_),
    .B1(_08526_),
    .Y(_08539_));
 sky130_fd_sc_hd__nand2_2 _30567_ (.A(_08529_),
    .B(_08535_),
    .Y(_08540_));
 sky130_fd_sc_hd__a21o_2 _30568_ (.A1(_08529_),
    .A2(_08534_),
    .B1(_08535_),
    .X(_08541_));
 sky130_fd_sc_hd__o2111ai_2 _30569_ (.A1(_08539_),
    .A2(_08540_),
    .B1(_08433_),
    .C1(_08441_),
    .D1(_08541_),
    .Y(_08542_));
 sky130_fd_sc_hd__nand3_2 _30570_ (.A(_08305_),
    .B(_08538_),
    .C(_08542_),
    .Y(_08543_));
 sky130_fd_sc_hd__a31oi_2 _30571_ (.A1(_08140_),
    .A2(_08259_),
    .A3(_08143_),
    .B1(_08265_),
    .Y(_08544_));
 sky130_fd_sc_hd__o211ai_2 _30572_ (.A1(_08536_),
    .A2(_08537_),
    .B1(_08433_),
    .C1(_08441_),
    .Y(_08545_));
 sky130_fd_sc_hd__nand2_2 _30573_ (.A(_08441_),
    .B(_08433_),
    .Y(_08546_));
 sky130_fd_sc_hd__nand3_2 _30574_ (.A(_08529_),
    .B(_08534_),
    .C(_08535_),
    .Y(_08547_));
 sky130_fd_sc_hd__nand3_2 _30575_ (.A(_08546_),
    .B(_08541_),
    .C(_08547_),
    .Y(_08548_));
 sky130_fd_sc_hd__nand3_2 _30576_ (.A(_08544_),
    .B(_08545_),
    .C(_08548_),
    .Y(_08549_));
 sky130_fd_sc_hd__nand2_2 _30577_ (.A(_08543_),
    .B(_08549_),
    .Y(_08550_));
 sky130_fd_sc_hd__nand2_2 _30578_ (.A(_08143_),
    .B(_08142_),
    .Y(_08551_));
 sky130_fd_sc_hd__a21oi_2 _30579_ (.A1(_08116_),
    .A2(_08121_),
    .B1(_08129_),
    .Y(_08552_));
 sky130_fd_sc_hd__nand2_2 _30580_ (.A(_08551_),
    .B(_08552_),
    .Y(_08553_));
 sky130_fd_sc_hd__a211o_2 _30581_ (.A1(_08141_),
    .A2(_08139_),
    .B1(_08138_),
    .C1(_08552_),
    .X(_08554_));
 sky130_fd_sc_hd__and2_2 _30582_ (.A(_08553_),
    .B(_08554_),
    .X(_08555_));
 sky130_fd_sc_hd__nand2_2 _30583_ (.A(_08550_),
    .B(_08555_),
    .Y(_08556_));
 sky130_fd_sc_hd__a21oi_2 _30584_ (.A1(_08270_),
    .A2(_08272_),
    .B1(_08273_),
    .Y(_08557_));
 sky130_fd_sc_hd__o21ai_2 _30585_ (.A1(_08285_),
    .A2(_08557_),
    .B1(_08274_),
    .Y(_08558_));
 sky130_fd_sc_hd__nand2_2 _30586_ (.A(_08553_),
    .B(_08554_),
    .Y(_08559_));
 sky130_fd_sc_hd__nand3_2 _30587_ (.A(_08543_),
    .B(_08549_),
    .C(_08559_),
    .Y(_08560_));
 sky130_fd_sc_hd__nand3_2 _30588_ (.A(_08556_),
    .B(_08558_),
    .C(_08560_),
    .Y(_08561_));
 sky130_fd_sc_hd__inv_2 _30589_ (.A(_08553_),
    .Y(_08562_));
 sky130_fd_sc_hd__inv_2 _30590_ (.A(_08554_),
    .Y(_08563_));
 sky130_fd_sc_hd__o2bb2ai_2 _30591_ (.A1_N(_08543_),
    .A2_N(_08549_),
    .B1(_08562_),
    .B2(_08563_),
    .Y(_08564_));
 sky130_fd_sc_hd__a21boi_2 _30592_ (.A1(_08269_),
    .A2(_08282_),
    .B1_N(_08274_),
    .Y(_08565_));
 sky130_fd_sc_hd__nand3_2 _30593_ (.A(_08555_),
    .B(_08543_),
    .C(_08549_),
    .Y(_08566_));
 sky130_fd_sc_hd__nand3_2 _30594_ (.A(_08564_),
    .B(_08565_),
    .C(_08566_),
    .Y(_08567_));
 sky130_fd_sc_hd__a21o_2 _30595_ (.A1(_08561_),
    .A2(_08567_),
    .B1(_08279_),
    .X(_08568_));
 sky130_fd_sc_hd__a21boi_2 _30596_ (.A1(_08298_),
    .A2(_08287_),
    .B1_N(_08291_),
    .Y(_08569_));
 sky130_fd_sc_hd__nand3_2 _30597_ (.A(_08561_),
    .B(_08567_),
    .C(_08279_),
    .Y(_08570_));
 sky130_fd_sc_hd__nand3_2 _30598_ (.A(_08568_),
    .B(_08569_),
    .C(_08570_),
    .Y(_08571_));
 sky130_fd_sc_hd__inv_2 _30599_ (.A(_08276_),
    .Y(_08572_));
 sky130_fd_sc_hd__o2bb2ai_2 _30600_ (.A1_N(_08561_),
    .A2_N(_08567_),
    .B1(_08280_),
    .B2(_08572_),
    .Y(_08573_));
 sky130_fd_sc_hd__inv_2 _30601_ (.A(_08290_),
    .Y(_08574_));
 sky130_fd_sc_hd__nand2_2 _30602_ (.A(_08288_),
    .B(_08289_),
    .Y(_08575_));
 sky130_fd_sc_hd__o2bb2ai_2 _30603_ (.A1_N(_08298_),
    .A2_N(_08287_),
    .B1(_08574_),
    .B2(_08575_),
    .Y(_08576_));
 sky130_fd_sc_hd__inv_2 _30604_ (.A(_08279_),
    .Y(_08577_));
 sky130_fd_sc_hd__nand3_2 _30605_ (.A(_08561_),
    .B(_08567_),
    .C(_08577_),
    .Y(_08578_));
 sky130_fd_sc_hd__nand3_2 _30606_ (.A(_08573_),
    .B(_08576_),
    .C(_08578_),
    .Y(_08579_));
 sky130_fd_sc_hd__and2_2 _30607_ (.A(_08571_),
    .B(_08579_),
    .X(_08580_));
 sky130_fd_sc_hd__o2111a_2 _30608_ (.A1(_07772_),
    .A2(_08040_),
    .B1(_07535_),
    .C1(_07540_),
    .D1(_07776_),
    .X(_08581_));
 sky130_fd_sc_hd__nand3_2 _30609_ (.A(_08581_),
    .B(_08037_),
    .C(_08301_),
    .Y(_08582_));
 sky130_fd_sc_hd__or3_2 _30610_ (.A(_07544_),
    .B(_08582_),
    .C(_06491_),
    .X(_08583_));
 sky130_fd_sc_hd__o2111a_2 _30611_ (.A1(_08020_),
    .A2(_08023_),
    .B1(_08297_),
    .C1(_08028_),
    .D1(_08299_),
    .X(_08584_));
 sky130_fd_sc_hd__o22ai_2 _30612_ (.A1(_08293_),
    .A2(_08296_),
    .B1(_08302_),
    .B2(_08584_),
    .Y(_08585_));
 sky130_fd_sc_hd__a31oi_2 _30613_ (.A1(_08037_),
    .A2(_08301_),
    .A3(_08039_),
    .B1(_08585_),
    .Y(_08586_));
 sky130_fd_sc_hd__o21ai_2 _30614_ (.A1(_08582_),
    .A2(_07547_),
    .B1(_08586_),
    .Y(_08587_));
 sky130_fd_sc_hd__inv_2 _30615_ (.A(_08587_),
    .Y(_08588_));
 sky130_fd_sc_hd__nand2_2 _30616_ (.A(_08583_),
    .B(_08588_),
    .Y(_08589_));
 sky130_fd_sc_hd__nor2_2 _30617_ (.A(_08580_),
    .B(_08589_),
    .Y(_08590_));
 sky130_fd_sc_hd__and2_2 _30618_ (.A(_08589_),
    .B(_08580_),
    .X(_08591_));
 sky130_fd_sc_hd__nor2_2 _30619_ (.A(_08590_),
    .B(_08591_),
    .Y(_02643_));
 sky130_fd_sc_hd__a21oi_2 _30620_ (.A1(_08564_),
    .A2(_08566_),
    .B1(_08565_),
    .Y(_08592_));
 sky130_fd_sc_hd__a21o_2 _30621_ (.A1(_08577_),
    .A2(_08567_),
    .B1(_08592_),
    .X(_08593_));
 sky130_fd_sc_hd__nand3_2 _30622_ (.A(_08541_),
    .B(_08440_),
    .C(_08547_),
    .Y(_08594_));
 sky130_fd_sc_hd__nand2_2 _30623_ (.A(_08594_),
    .B(_08433_),
    .Y(_08595_));
 sky130_fd_sc_hd__buf_1 _30624_ (.A(_19584_),
    .X(_08596_));
 sky130_fd_sc_hd__a22oi_2 _30625_ (.A1(_05851_),
    .A2(_06728_),
    .B1(_06508_),
    .B2(_08596_),
    .Y(_08597_));
 sky130_fd_sc_hd__inv_2 _30626_ (.A(\pcpi_mul.rs1[18] ),
    .Y(_08598_));
 sky130_fd_sc_hd__nand3_2 _30627_ (.A(_05758_),
    .B(_05641_),
    .C(_06944_),
    .Y(_08599_));
 sky130_fd_sc_hd__nor2_2 _30628_ (.A(_08598_),
    .B(_08599_),
    .Y(_08600_));
 sky130_fd_sc_hd__nand2_2 _30629_ (.A(_06496_),
    .B(_07138_),
    .Y(_08601_));
 sky130_fd_sc_hd__o21ai_2 _30630_ (.A1(_08597_),
    .A2(_08600_),
    .B1(_08601_),
    .Y(_08602_));
 sky130_fd_sc_hd__o21ai_2 _30631_ (.A1(_08329_),
    .A2(_08325_),
    .B1(_08332_),
    .Y(_08603_));
 sky130_fd_sc_hd__buf_1 _30632_ (.A(_08598_),
    .X(_08604_));
 sky130_fd_sc_hd__inv_2 _30633_ (.A(_08601_),
    .Y(_08605_));
 sky130_fd_sc_hd__a22o_2 _30634_ (.A1(_05857_),
    .A2(_06728_),
    .B1(_06896_),
    .B2(_08596_),
    .X(_08606_));
 sky130_fd_sc_hd__o211ai_2 _30635_ (.A1(_08604_),
    .A2(_08599_),
    .B1(_08605_),
    .C1(_08606_),
    .Y(_08607_));
 sky130_fd_sc_hd__nand3_2 _30636_ (.A(_08602_),
    .B(_08603_),
    .C(_08607_),
    .Y(_08608_));
 sky130_fd_sc_hd__o21ai_2 _30637_ (.A1(_08597_),
    .A2(_08600_),
    .B1(_08605_),
    .Y(_08609_));
 sky130_fd_sc_hd__a31oi_2 _30638_ (.A1(_08333_),
    .A2(_06020_),
    .A3(_19595_),
    .B1(_08328_),
    .Y(_08610_));
 sky130_fd_sc_hd__buf_1 _30639_ (.A(_08598_),
    .X(_08611_));
 sky130_fd_sc_hd__o211ai_2 _30640_ (.A1(_08611_),
    .A2(_08599_),
    .B1(_08601_),
    .C1(_08606_),
    .Y(_08612_));
 sky130_fd_sc_hd__nand3_2 _30641_ (.A(_08609_),
    .B(_08610_),
    .C(_08612_),
    .Y(_08613_));
 sky130_fd_sc_hd__nor2_2 _30642_ (.A(_08449_),
    .B(_08443_),
    .Y(_08614_));
 sky130_fd_sc_hd__o2bb2ai_2 _30643_ (.A1_N(_08608_),
    .A2_N(_08613_),
    .B1(_08442_),
    .B2(_08614_),
    .Y(_08615_));
 sky130_fd_sc_hd__nor2_2 _30644_ (.A(_08442_),
    .B(_08614_),
    .Y(_08616_));
 sky130_fd_sc_hd__nand3_2 _30645_ (.A(_08613_),
    .B(_08608_),
    .C(_08616_),
    .Y(_08617_));
 sky130_fd_sc_hd__nand2_2 _30646_ (.A(_08324_),
    .B(_08335_),
    .Y(_08618_));
 sky130_fd_sc_hd__nand2_2 _30647_ (.A(_08618_),
    .B(_08318_),
    .Y(_08619_));
 sky130_fd_sc_hd__a21oi_2 _30648_ (.A1(_08615_),
    .A2(_08617_),
    .B1(_08619_),
    .Y(_08620_));
 sky130_fd_sc_hd__nand2_2 _30649_ (.A(_08613_),
    .B(_08616_),
    .Y(_08621_));
 sky130_fd_sc_hd__inv_2 _30650_ (.A(_08608_),
    .Y(_08622_));
 sky130_fd_sc_hd__o211a_2 _30651_ (.A1(_08621_),
    .A2(_08622_),
    .B1(_08615_),
    .C1(_08619_),
    .X(_08623_));
 sky130_fd_sc_hd__nand2_2 _30652_ (.A(_08460_),
    .B(_08461_),
    .Y(_08624_));
 sky130_fd_sc_hd__o21ai_2 _30653_ (.A1(_08620_),
    .A2(_08623_),
    .B1(_08624_),
    .Y(_08625_));
 sky130_fd_sc_hd__nand2_2 _30654_ (.A(_08464_),
    .B(_08462_),
    .Y(_08626_));
 sky130_fd_sc_hd__a2bb2oi_2 _30655_ (.A1_N(_08468_),
    .A2_N(_08626_),
    .B1(_08470_),
    .B2(_08469_),
    .Y(_08627_));
 sky130_fd_sc_hd__a21o_2 _30656_ (.A1(_08615_),
    .A2(_08617_),
    .B1(_08619_),
    .X(_08628_));
 sky130_fd_sc_hd__nand3_2 _30657_ (.A(_08619_),
    .B(_08615_),
    .C(_08617_),
    .Y(_08629_));
 sky130_fd_sc_hd__inv_2 _30658_ (.A(_08624_),
    .Y(_08630_));
 sky130_fd_sc_hd__nand3_2 _30659_ (.A(_08628_),
    .B(_08629_),
    .C(_08630_),
    .Y(_08631_));
 sky130_fd_sc_hd__nand3_2 _30660_ (.A(_08625_),
    .B(_08627_),
    .C(_08631_),
    .Y(_08632_));
 sky130_fd_sc_hd__inv_2 _30661_ (.A(_08457_),
    .Y(_08633_));
 sky130_fd_sc_hd__nor2_2 _30662_ (.A(_08459_),
    .B(_08453_),
    .Y(_08634_));
 sky130_fd_sc_hd__o22ai_2 _30663_ (.A1(_08633_),
    .A2(_08634_),
    .B1(_08620_),
    .B2(_08623_),
    .Y(_08635_));
 sky130_fd_sc_hd__o21ai_2 _30664_ (.A1(_08475_),
    .A2(_08474_),
    .B1(_08481_),
    .Y(_08636_));
 sky130_fd_sc_hd__nand3_2 _30665_ (.A(_08628_),
    .B(_08629_),
    .C(_08624_),
    .Y(_08637_));
 sky130_fd_sc_hd__nand3_2 _30666_ (.A(_08635_),
    .B(_08636_),
    .C(_08637_),
    .Y(_08638_));
 sky130_fd_sc_hd__nand2_2 _30667_ (.A(_08632_),
    .B(_08638_),
    .Y(_08639_));
 sky130_fd_sc_hd__o21ai_2 _30668_ (.A1(_08505_),
    .A2(_08494_),
    .B1(_08512_),
    .Y(_08640_));
 sky130_fd_sc_hd__a21o_2 _30669_ (.A1(_08488_),
    .A2(_08486_),
    .B1(_08485_),
    .X(_08641_));
 sky130_fd_sc_hd__nand2_2 _30670_ (.A(_06731_),
    .B(_07594_),
    .Y(_08642_));
 sky130_fd_sc_hd__nand2_2 _30671_ (.A(_05891_),
    .B(_19577_),
    .Y(_08643_));
 sky130_fd_sc_hd__or2_2 _30672_ (.A(_08642_),
    .B(_08643_),
    .X(_08644_));
 sky130_fd_sc_hd__buf_1 _30673_ (.A(\pcpi_mul.rs1[25] ),
    .X(_08645_));
 sky130_fd_sc_hd__nand2_2 _30674_ (.A(_05192_),
    .B(_08645_),
    .Y(_08646_));
 sky130_fd_sc_hd__inv_2 _30675_ (.A(_08646_),
    .Y(_08647_));
 sky130_fd_sc_hd__nand2_2 _30676_ (.A(_08642_),
    .B(_08643_),
    .Y(_08648_));
 sky130_fd_sc_hd__nand3_2 _30677_ (.A(_08644_),
    .B(_08647_),
    .C(_08648_),
    .Y(_08649_));
 sky130_fd_sc_hd__buf_1 _30678_ (.A(_07594_),
    .X(_08650_));
 sky130_fd_sc_hd__buf_1 _30679_ (.A(_07605_),
    .X(_08651_));
 sky130_fd_sc_hd__a22oi_2 _30680_ (.A1(_06735_),
    .A2(_08650_),
    .B1(_05403_),
    .B2(_08651_),
    .Y(_08652_));
 sky130_fd_sc_hd__nor2_2 _30681_ (.A(_08642_),
    .B(_08643_),
    .Y(_08653_));
 sky130_fd_sc_hd__o21ai_2 _30682_ (.A1(_08652_),
    .A2(_08653_),
    .B1(_08646_),
    .Y(_08654_));
 sky130_fd_sc_hd__nand3_2 _30683_ (.A(_08641_),
    .B(_08649_),
    .C(_08654_),
    .Y(_08655_));
 sky130_fd_sc_hd__nand3_2 _30684_ (.A(_08644_),
    .B(_08646_),
    .C(_08648_),
    .Y(_08656_));
 sky130_fd_sc_hd__a21oi_2 _30685_ (.A1(_08488_),
    .A2(_08486_),
    .B1(_08485_),
    .Y(_08657_));
 sky130_fd_sc_hd__o21ai_2 _30686_ (.A1(_08652_),
    .A2(_08653_),
    .B1(_08647_),
    .Y(_08658_));
 sky130_fd_sc_hd__nand3_2 _30687_ (.A(_08656_),
    .B(_08657_),
    .C(_08658_),
    .Y(_08659_));
 sky130_fd_sc_hd__nand2_2 _30688_ (.A(_08655_),
    .B(_08659_),
    .Y(_08660_));
 sky130_fd_sc_hd__buf_1 _30689_ (.A(\pcpi_mul.rs1[24] ),
    .X(_08661_));
 sky130_fd_sc_hd__buf_1 _30690_ (.A(_08661_),
    .X(_08662_));
 sky130_fd_sc_hd__a22oi_2 _30691_ (.A1(_06072_),
    .A2(_08496_),
    .B1(_19401_),
    .B2(_08662_),
    .Y(_08663_));
 sky130_fd_sc_hd__buf_1 _30692_ (.A(\pcpi_mul.rs1[24] ),
    .X(_08664_));
 sky130_fd_sc_hd__and4_2 _30693_ (.A(_05123_),
    .B(_05909_),
    .C(_08664_),
    .D(_08496_),
    .X(_08665_));
 sky130_fd_sc_hd__nor2_2 _30694_ (.A(_08663_),
    .B(_08665_),
    .Y(_08666_));
 sky130_fd_sc_hd__inv_2 _30695_ (.A(_07837_),
    .Y(_08667_));
 sky130_fd_sc_hd__nor2_2 _30696_ (.A(_05149_),
    .B(_08667_),
    .Y(_08668_));
 sky130_fd_sc_hd__nand2_2 _30697_ (.A(_08666_),
    .B(_08668_),
    .Y(_08669_));
 sky130_fd_sc_hd__inv_2 _30698_ (.A(_08668_),
    .Y(_08670_));
 sky130_fd_sc_hd__o21ai_2 _30699_ (.A1(_08663_),
    .A2(_08665_),
    .B1(_08670_),
    .Y(_08671_));
 sky130_fd_sc_hd__nand2_2 _30700_ (.A(_08669_),
    .B(_08671_),
    .Y(_08672_));
 sky130_fd_sc_hd__nand2_2 _30701_ (.A(_08660_),
    .B(_08672_),
    .Y(_08673_));
 sky130_fd_sc_hd__nand2_2 _30702_ (.A(_08666_),
    .B(_08670_),
    .Y(_08674_));
 sky130_fd_sc_hd__o21ai_2 _30703_ (.A1(_08663_),
    .A2(_08665_),
    .B1(_08668_),
    .Y(_08675_));
 sky130_fd_sc_hd__nand2_2 _30704_ (.A(_08674_),
    .B(_08675_),
    .Y(_08676_));
 sky130_fd_sc_hd__nand3_2 _30705_ (.A(_08676_),
    .B(_08655_),
    .C(_08659_),
    .Y(_08677_));
 sky130_fd_sc_hd__nand3_2 _30706_ (.A(_08640_),
    .B(_08673_),
    .C(_08677_),
    .Y(_08678_));
 sky130_fd_sc_hd__inv_2 _30707_ (.A(_08678_),
    .Y(_08679_));
 sky130_fd_sc_hd__nand3_2 _30708_ (.A(_08672_),
    .B(_08655_),
    .C(_08659_),
    .Y(_08680_));
 sky130_fd_sc_hd__nand2_2 _30709_ (.A(_08660_),
    .B(_08676_),
    .Y(_08681_));
 sky130_fd_sc_hd__o2111ai_2 _30710_ (.A1(_08505_),
    .A2(_08494_),
    .B1(_08512_),
    .C1(_08680_),
    .D1(_08681_),
    .Y(_08682_));
 sky130_fd_sc_hd__nor2_2 _30711_ (.A(_08498_),
    .B(_08500_),
    .Y(_08683_));
 sky130_fd_sc_hd__a21oi_2 _30712_ (.A1(_08499_),
    .A2(_08501_),
    .B1(_08502_),
    .Y(_08684_));
 sky130_fd_sc_hd__nor2_2 _30713_ (.A(_08683_),
    .B(_08684_),
    .Y(_08685_));
 sky130_fd_sc_hd__inv_2 _30714_ (.A(_08685_),
    .Y(_08686_));
 sky130_fd_sc_hd__nand2_2 _30715_ (.A(_08682_),
    .B(_08686_),
    .Y(_08687_));
 sky130_fd_sc_hd__nand2_2 _30716_ (.A(_08682_),
    .B(_08678_),
    .Y(_08688_));
 sky130_fd_sc_hd__nand2_2 _30717_ (.A(_08688_),
    .B(_08685_),
    .Y(_08689_));
 sky130_fd_sc_hd__o21ai_2 _30718_ (.A1(_08679_),
    .A2(_08687_),
    .B1(_08689_),
    .Y(_08690_));
 sky130_fd_sc_hd__nand2_2 _30719_ (.A(_08639_),
    .B(_08690_),
    .Y(_08691_));
 sky130_fd_sc_hd__nand2_2 _30720_ (.A(_08438_),
    .B(_08370_),
    .Y(_08692_));
 sky130_fd_sc_hd__nand2_2 _30721_ (.A(_08688_),
    .B(_08686_),
    .Y(_08693_));
 sky130_fd_sc_hd__nand3_2 _30722_ (.A(_08682_),
    .B(_08678_),
    .C(_08685_),
    .Y(_08694_));
 sky130_fd_sc_hd__nand2_2 _30723_ (.A(_08693_),
    .B(_08694_),
    .Y(_08695_));
 sky130_fd_sc_hd__nand3_2 _30724_ (.A(_08695_),
    .B(_08632_),
    .C(_08638_),
    .Y(_08696_));
 sky130_fd_sc_hd__nand3_2 _30725_ (.A(_08691_),
    .B(_08692_),
    .C(_08696_),
    .Y(_08697_));
 sky130_fd_sc_hd__buf_1 _30726_ (.A(_08697_),
    .X(_08698_));
 sky130_fd_sc_hd__inv_2 _30727_ (.A(_08694_),
    .Y(_08699_));
 sky130_fd_sc_hd__and2_2 _30728_ (.A(_08688_),
    .B(_08686_),
    .X(_08700_));
 sky130_fd_sc_hd__o2bb2ai_2 _30729_ (.A1_N(_08638_),
    .A2_N(_08632_),
    .B1(_08699_),
    .B2(_08700_),
    .Y(_08701_));
 sky130_fd_sc_hd__nand2_2 _30730_ (.A(_08367_),
    .B(_08368_),
    .Y(_08702_));
 sky130_fd_sc_hd__a21oi_2 _30731_ (.A1(_08702_),
    .A2(_08374_),
    .B1(_08372_),
    .Y(_08703_));
 sky130_fd_sc_hd__a22oi_2 _30732_ (.A1(_08703_),
    .A2(_08369_),
    .B1(_08376_),
    .B2(_08379_),
    .Y(_08704_));
 sky130_fd_sc_hd__nand3_2 _30733_ (.A(_08690_),
    .B(_08632_),
    .C(_08638_),
    .Y(_08705_));
 sky130_fd_sc_hd__nand3_2 _30734_ (.A(_08701_),
    .B(_08704_),
    .C(_08705_),
    .Y(_08706_));
 sky130_fd_sc_hd__inv_2 _30735_ (.A(_08477_),
    .Y(_08707_));
 sky130_fd_sc_hd__a21o_2 _30736_ (.A1(_08524_),
    .A2(_08483_),
    .B1(_08707_),
    .X(_08708_));
 sky130_fd_sc_hd__a21oi_2 _30737_ (.A1(_08698_),
    .A2(_08706_),
    .B1(_08708_),
    .Y(_08709_));
 sky130_fd_sc_hd__and2_2 _30738_ (.A(_08524_),
    .B(_08483_),
    .X(_08710_));
 sky130_fd_sc_hd__o211a_2 _30739_ (.A1(_08707_),
    .A2(_08710_),
    .B1(_08706_),
    .C1(_08697_),
    .X(_08711_));
 sky130_fd_sc_hd__a22oi_2 _30740_ (.A1(_08182_),
    .A2(_05506_),
    .B1(_07652_),
    .B2(_06492_),
    .Y(_08712_));
 sky130_fd_sc_hd__nand3_2 _30741_ (.A(_07416_),
    .B(_06827_),
    .C(_05408_),
    .Y(_08713_));
 sky130_fd_sc_hd__nor2_2 _30742_ (.A(_06494_),
    .B(_08713_),
    .Y(_08714_));
 sky130_fd_sc_hd__nand2_2 _30743_ (.A(_07890_),
    .B(_06497_),
    .Y(_08715_));
 sky130_fd_sc_hd__inv_2 _30744_ (.A(_08715_),
    .Y(_08716_));
 sky130_fd_sc_hd__o21ai_2 _30745_ (.A1(_08712_),
    .A2(_08714_),
    .B1(_08716_),
    .Y(_08717_));
 sky130_fd_sc_hd__a31oi_2 _30746_ (.A1(_08411_),
    .A2(_19352_),
    .A3(_19623_),
    .B1(_08406_),
    .Y(_08718_));
 sky130_fd_sc_hd__a22o_2 _30747_ (.A1(_08182_),
    .A2(_06162_),
    .B1(_19357_),
    .B2(_06492_),
    .X(_08719_));
 sky130_fd_sc_hd__o211ai_2 _30748_ (.A1(_06494_),
    .A2(_08713_),
    .B1(_08715_),
    .C1(_08719_),
    .Y(_08720_));
 sky130_fd_sc_hd__nand3_2 _30749_ (.A(_08717_),
    .B(_08718_),
    .C(_08720_),
    .Y(_08721_));
 sky130_fd_sc_hd__o21ai_2 _30750_ (.A1(_08712_),
    .A2(_08714_),
    .B1(_08715_),
    .Y(_08722_));
 sky130_fd_sc_hd__o21ai_2 _30751_ (.A1(_08408_),
    .A2(_08403_),
    .B1(_08410_),
    .Y(_08723_));
 sky130_fd_sc_hd__o211ai_2 _30752_ (.A1(_06505_),
    .A2(_08713_),
    .B1(_08716_),
    .C1(_08719_),
    .Y(_08724_));
 sky130_fd_sc_hd__nand3_2 _30753_ (.A(_08722_),
    .B(_08723_),
    .C(_08724_),
    .Y(_08725_));
 sky130_fd_sc_hd__a21o_2 _30754_ (.A1(_08346_),
    .A2(_08342_),
    .B1(_08341_),
    .X(_08726_));
 sky130_fd_sc_hd__a21oi_2 _30755_ (.A1(_08721_),
    .A2(_08725_),
    .B1(_08726_),
    .Y(_08727_));
 sky130_fd_sc_hd__nand3_2 _30756_ (.A(_08721_),
    .B(_08725_),
    .C(_08726_),
    .Y(_08728_));
 sky130_fd_sc_hd__o21ai_2 _30757_ (.A1(_08176_),
    .A2(_08355_),
    .B1(_08348_),
    .Y(_08729_));
 sky130_fd_sc_hd__nand3_2 _30758_ (.A(_08728_),
    .B(_08354_),
    .C(_08729_),
    .Y(_08730_));
 sky130_fd_sc_hd__nor2_2 _30759_ (.A(_08727_),
    .B(_08730_),
    .Y(_08731_));
 sky130_fd_sc_hd__nand2_2 _30760_ (.A(_08721_),
    .B(_08725_),
    .Y(_08732_));
 sky130_fd_sc_hd__a21oi_2 _30761_ (.A1(_08346_),
    .A2(_08342_),
    .B1(_08341_),
    .Y(_08733_));
 sky130_fd_sc_hd__nand2_2 _30762_ (.A(_08732_),
    .B(_08733_),
    .Y(_08734_));
 sky130_fd_sc_hd__nand2_2 _30763_ (.A(_08354_),
    .B(_08357_),
    .Y(_08735_));
 sky130_fd_sc_hd__nand2_2 _30764_ (.A(_08735_),
    .B(_08348_),
    .Y(_08736_));
 sky130_fd_sc_hd__a21oi_2 _30765_ (.A1(_08734_),
    .A2(_08728_),
    .B1(_08736_),
    .Y(_08737_));
 sky130_fd_sc_hd__and4_2 _30766_ (.A(_06441_),
    .B(_19365_),
    .C(_06732_),
    .D(_06369_),
    .X(_08738_));
 sky130_fd_sc_hd__a22o_2 _30767_ (.A1(_07012_),
    .A2(_05717_),
    .B1(_07020_),
    .B2(_07939_),
    .X(_08739_));
 sky130_fd_sc_hd__nand2_2 _30768_ (.A(_19367_),
    .B(_19599_),
    .Y(_08740_));
 sky130_fd_sc_hd__inv_2 _30769_ (.A(_08740_),
    .Y(_08741_));
 sky130_fd_sc_hd__nand2_2 _30770_ (.A(_08739_),
    .B(_08741_),
    .Y(_08742_));
 sky130_fd_sc_hd__a22oi_2 _30771_ (.A1(_19363_),
    .A2(_19606_),
    .B1(_06276_),
    .B2(_05897_),
    .Y(_08743_));
 sky130_fd_sc_hd__o21ai_2 _30772_ (.A1(_08743_),
    .A2(_08738_),
    .B1(_08740_),
    .Y(_08744_));
 sky130_fd_sc_hd__nand2_2 _30773_ (.A(_08313_),
    .B(_08321_),
    .Y(_08745_));
 sky130_fd_sc_hd__o211ai_2 _30774_ (.A1(_08738_),
    .A2(_08742_),
    .B1(_08744_),
    .C1(_08745_),
    .Y(_08746_));
 sky130_fd_sc_hd__o21ai_2 _30775_ (.A1(_08743_),
    .A2(_08738_),
    .B1(_08741_),
    .Y(_08747_));
 sky130_fd_sc_hd__nand2_2 _30776_ (.A(_06441_),
    .B(_05910_),
    .Y(_08748_));
 sky130_fd_sc_hd__nand3b_2 _30777_ (.A_N(_08748_),
    .B(_07934_),
    .C(_19603_),
    .Y(_08749_));
 sky130_fd_sc_hd__nand3_2 _30778_ (.A(_08749_),
    .B(_08740_),
    .C(_08739_),
    .Y(_08750_));
 sky130_fd_sc_hd__a21oi_2 _30779_ (.A1(_08311_),
    .A2(_08312_),
    .B1(_08309_),
    .Y(_08751_));
 sky130_fd_sc_hd__nand3_2 _30780_ (.A(_08747_),
    .B(_08750_),
    .C(_08751_),
    .Y(_08752_));
 sky130_fd_sc_hd__nand2_2 _30781_ (.A(_08746_),
    .B(_08752_),
    .Y(_08753_));
 sky130_fd_sc_hd__a22oi_2 _30782_ (.A1(_06256_),
    .A2(_06206_),
    .B1(_05670_),
    .B2(_06560_),
    .Y(_08754_));
 sky130_fd_sc_hd__and4_2 _30783_ (.A(_19370_),
    .B(_05802_),
    .C(_06957_),
    .D(_19596_),
    .X(_08755_));
 sky130_fd_sc_hd__nand2_2 _30784_ (.A(_19375_),
    .B(_07360_),
    .Y(_08756_));
 sky130_fd_sc_hd__inv_2 _30785_ (.A(_08756_),
    .Y(_08757_));
 sky130_fd_sc_hd__o21ai_2 _30786_ (.A1(_08754_),
    .A2(_08755_),
    .B1(_08757_),
    .Y(_08758_));
 sky130_fd_sc_hd__nand2_2 _30787_ (.A(_19370_),
    .B(_19596_),
    .Y(_08759_));
 sky130_fd_sc_hd__nand3b_2 _30788_ (.A_N(_08759_),
    .B(_05803_),
    .C(_07798_),
    .Y(_08760_));
 sky130_fd_sc_hd__buf_1 _30789_ (.A(_06205_),
    .X(_08761_));
 sky130_fd_sc_hd__a22o_2 _30790_ (.A1(_07203_),
    .A2(_08761_),
    .B1(_19373_),
    .B2(_06373_),
    .X(_08762_));
 sky130_fd_sc_hd__nand3_2 _30791_ (.A(_08760_),
    .B(_08756_),
    .C(_08762_),
    .Y(_08763_));
 sky130_fd_sc_hd__nand2_2 _30792_ (.A(_08758_),
    .B(_08763_),
    .Y(_08764_));
 sky130_fd_sc_hd__nand2_2 _30793_ (.A(_08753_),
    .B(_08764_),
    .Y(_08765_));
 sky130_fd_sc_hd__inv_2 _30794_ (.A(_08764_),
    .Y(_08766_));
 sky130_fd_sc_hd__nand3_2 _30795_ (.A(_08766_),
    .B(_08746_),
    .C(_08752_),
    .Y(_08767_));
 sky130_fd_sc_hd__nand2_2 _30796_ (.A(_08765_),
    .B(_08767_),
    .Y(_08768_));
 sky130_fd_sc_hd__o21ai_2 _30797_ (.A1(_08731_),
    .A2(_08737_),
    .B1(_08768_),
    .Y(_08769_));
 sky130_fd_sc_hd__a21o_2 _30798_ (.A1(_08734_),
    .A2(_08728_),
    .B1(_08736_),
    .X(_08770_));
 sky130_fd_sc_hd__nand3_2 _30799_ (.A(_08734_),
    .B(_08736_),
    .C(_08728_),
    .Y(_08771_));
 sky130_fd_sc_hd__nand2_2 _30800_ (.A(_08753_),
    .B(_08766_),
    .Y(_08772_));
 sky130_fd_sc_hd__nand3_2 _30801_ (.A(_08746_),
    .B(_08752_),
    .C(_08764_),
    .Y(_08773_));
 sky130_fd_sc_hd__nand2_2 _30802_ (.A(_08772_),
    .B(_08773_),
    .Y(_08774_));
 sky130_fd_sc_hd__nand3_2 _30803_ (.A(_08770_),
    .B(_08771_),
    .C(_08774_),
    .Y(_08775_));
 sky130_fd_sc_hd__nand3_2 _30804_ (.A(_08769_),
    .B(_08422_),
    .C(_08775_),
    .Y(_08776_));
 sky130_fd_sc_hd__inv_2 _30805_ (.A(_08773_),
    .Y(_08777_));
 sky130_fd_sc_hd__inv_2 _30806_ (.A(_08772_),
    .Y(_08778_));
 sky130_fd_sc_hd__o22ai_2 _30807_ (.A1(_08777_),
    .A2(_08778_),
    .B1(_08731_),
    .B2(_08737_),
    .Y(_08779_));
 sky130_fd_sc_hd__inv_2 _30808_ (.A(_08421_),
    .Y(_08780_));
 sky130_fd_sc_hd__nand3_2 _30809_ (.A(_08770_),
    .B(_08771_),
    .C(_08768_),
    .Y(_08781_));
 sky130_fd_sc_hd__nand3_2 _30810_ (.A(_08779_),
    .B(_08780_),
    .C(_08781_),
    .Y(_08782_));
 sky130_fd_sc_hd__o21ai_2 _30811_ (.A1(_08359_),
    .A2(_08374_),
    .B1(_08368_),
    .Y(_08783_));
 sky130_fd_sc_hd__a21oi_2 _30812_ (.A1(_08776_),
    .A2(_08782_),
    .B1(_08783_),
    .Y(_08784_));
 sky130_fd_sc_hd__and3_2 _30813_ (.A(_08776_),
    .B(_08782_),
    .C(_08783_),
    .X(_08785_));
 sky130_fd_sc_hd__nand2_2 _30814_ (.A(_08419_),
    .B(_08422_),
    .Y(_08786_));
 sky130_fd_sc_hd__and4_2 _30815_ (.A(_19332_),
    .B(_19334_),
    .C(_19637_),
    .D(_19641_),
    .X(_08787_));
 sky130_fd_sc_hd__inv_2 _30816_ (.A(_08787_),
    .Y(_08788_));
 sky130_fd_sc_hd__a22o_2 _30817_ (.A1(_19332_),
    .A2(_19642_),
    .B1(_19335_),
    .B2(_19638_),
    .X(_08789_));
 sky130_fd_sc_hd__buf_1 _30818_ (.A(_19336_),
    .X(_08790_));
 sky130_fd_sc_hd__buf_1 _30819_ (.A(\pcpi_mul.rs2[22] ),
    .X(_08791_));
 sky130_fd_sc_hd__a22oi_2 _30820_ (.A1(_08790_),
    .A2(_08393_),
    .B1(_08791_),
    .B2(_05204_),
    .Y(_08792_));
 sky130_fd_sc_hd__and4_2 _30821_ (.A(_08396_),
    .B(_07974_),
    .C(_05330_),
    .D(_19633_),
    .X(_08793_));
 sky130_fd_sc_hd__nand2_2 _30822_ (.A(_19342_),
    .B(_19627_),
    .Y(_08794_));
 sky130_fd_sc_hd__inv_2 _30823_ (.A(_08794_),
    .Y(_08795_));
 sky130_fd_sc_hd__o21ai_2 _30824_ (.A1(_08792_),
    .A2(_08793_),
    .B1(_08795_),
    .Y(_08796_));
 sky130_fd_sc_hd__a21oi_2 _30825_ (.A1(_08397_),
    .A2(_08395_),
    .B1(_08387_),
    .Y(_08797_));
 sky130_fd_sc_hd__nand2_2 _30826_ (.A(_08385_),
    .B(_05545_),
    .Y(_08798_));
 sky130_fd_sc_hd__buf_1 _30827_ (.A(_08386_),
    .X(_08799_));
 sky130_fd_sc_hd__nand3b_2 _30828_ (.A_N(_08798_),
    .B(_08799_),
    .C(_06622_),
    .Y(_08800_));
 sky130_fd_sc_hd__a22o_2 _30829_ (.A1(_08790_),
    .A2(_19633_),
    .B1(_08791_),
    .B2(_05204_),
    .X(_08801_));
 sky130_fd_sc_hd__nand3_2 _30830_ (.A(_08800_),
    .B(_08801_),
    .C(_08794_),
    .Y(_08802_));
 sky130_fd_sc_hd__nand3_2 _30831_ (.A(_08796_),
    .B(_08797_),
    .C(_08802_),
    .Y(_08803_));
 sky130_fd_sc_hd__o21ai_2 _30832_ (.A1(_08792_),
    .A2(_08793_),
    .B1(_08794_),
    .Y(_08804_));
 sky130_fd_sc_hd__nand3_2 _30833_ (.A(_08800_),
    .B(_08801_),
    .C(_08795_),
    .Y(_08805_));
 sky130_fd_sc_hd__o21ai_2 _30834_ (.A1(_08389_),
    .A2(_08384_),
    .B1(_08394_),
    .Y(_08806_));
 sky130_fd_sc_hd__nand3_2 _30835_ (.A(_08804_),
    .B(_08805_),
    .C(_08806_),
    .Y(_08807_));
 sky130_fd_sc_hd__buf_1 _30836_ (.A(_07722_),
    .X(_08808_));
 sky130_fd_sc_hd__buf_1 _30837_ (.A(_19349_),
    .X(_08809_));
 sky130_fd_sc_hd__a22oi_2 _30838_ (.A1(_08808_),
    .A2(_19626_),
    .B1(_08809_),
    .B2(_19623_),
    .Y(_08810_));
 sky130_fd_sc_hd__nand2_2 _30839_ (.A(_07722_),
    .B(_05194_),
    .Y(_08811_));
 sky130_fd_sc_hd__nand2_2 _30840_ (.A(_08159_),
    .B(_06614_),
    .Y(_08812_));
 sky130_fd_sc_hd__nor2_2 _30841_ (.A(_08811_),
    .B(_08812_),
    .Y(_08813_));
 sky130_fd_sc_hd__nand2_2 _30842_ (.A(_08407_),
    .B(_05421_),
    .Y(_08814_));
 sky130_fd_sc_hd__o21bai_2 _30843_ (.A1(_08810_),
    .A2(_08813_),
    .B1_N(_08814_),
    .Y(_08815_));
 sky130_fd_sc_hd__buf_1 _30844_ (.A(_07723_),
    .X(_08816_));
 sky130_fd_sc_hd__nand3b_2 _30845_ (.A_N(_08811_),
    .B(_08816_),
    .C(_19623_),
    .Y(_08817_));
 sky130_fd_sc_hd__nand2_2 _30846_ (.A(_08811_),
    .B(_08812_),
    .Y(_08818_));
 sky130_fd_sc_hd__nand3_2 _30847_ (.A(_08817_),
    .B(_08814_),
    .C(_08818_),
    .Y(_08819_));
 sky130_fd_sc_hd__nand2_2 _30848_ (.A(_08815_),
    .B(_08819_),
    .Y(_08820_));
 sky130_fd_sc_hd__a21o_2 _30849_ (.A1(_08803_),
    .A2(_08807_),
    .B1(_08820_),
    .X(_08821_));
 sky130_fd_sc_hd__nand3_2 _30850_ (.A(_08803_),
    .B(_08807_),
    .C(_08820_),
    .Y(_08822_));
 sky130_fd_sc_hd__nand2_2 _30851_ (.A(_08402_),
    .B(_08413_),
    .Y(_08823_));
 sky130_fd_sc_hd__nand2_2 _30852_ (.A(_08823_),
    .B(_08399_),
    .Y(_08824_));
 sky130_fd_sc_hd__a21o_2 _30853_ (.A1(_08821_),
    .A2(_08822_),
    .B1(_08824_),
    .X(_08825_));
 sky130_fd_sc_hd__nand3_2 _30854_ (.A(_08821_),
    .B(_08824_),
    .C(_08822_),
    .Y(_08826_));
 sky130_fd_sc_hd__a22oi_2 _30855_ (.A1(_08788_),
    .A2(_08789_),
    .B1(_08825_),
    .B2(_08826_),
    .Y(_08827_));
 sky130_fd_sc_hd__nand2_2 _30856_ (.A(_08788_),
    .B(_08789_),
    .Y(_08828_));
 sky130_fd_sc_hd__a21oi_2 _30857_ (.A1(_08821_),
    .A2(_08822_),
    .B1(_08824_),
    .Y(_08829_));
 sky130_fd_sc_hd__and3_2 _30858_ (.A(_08821_),
    .B(_08824_),
    .C(_08822_),
    .X(_08830_));
 sky130_fd_sc_hd__nor3_2 _30859_ (.A(_08828_),
    .B(_08829_),
    .C(_08830_),
    .Y(_08831_));
 sky130_fd_sc_hd__o22ai_2 _30860_ (.A1(_08427_),
    .A2(_08786_),
    .B1(_08827_),
    .B2(_08831_),
    .Y(_08832_));
 sky130_fd_sc_hd__o21ai_2 _30861_ (.A1(_08829_),
    .A2(_08830_),
    .B1(_08828_),
    .Y(_08833_));
 sky130_fd_sc_hd__nand3b_2 _30862_ (.A_N(_08828_),
    .B(_08825_),
    .C(_08826_),
    .Y(_08834_));
 sky130_fd_sc_hd__nand3_2 _30863_ (.A(_08429_),
    .B(_08833_),
    .C(_08834_),
    .Y(_08835_));
 sky130_fd_sc_hd__nand2_2 _30864_ (.A(_08832_),
    .B(_08835_),
    .Y(_08836_));
 sky130_fd_sc_hd__o21bai_2 _30865_ (.A1(_08784_),
    .A2(_08785_),
    .B1_N(_08836_),
    .Y(_08837_));
 sky130_fd_sc_hd__a21o_2 _30866_ (.A1(_08776_),
    .A2(_08782_),
    .B1(_08783_),
    .X(_08838_));
 sky130_fd_sc_hd__nand3_2 _30867_ (.A(_08776_),
    .B(_08782_),
    .C(_08783_),
    .Y(_08839_));
 sky130_fd_sc_hd__nand3_2 _30868_ (.A(_08838_),
    .B(_08836_),
    .C(_08839_),
    .Y(_08840_));
 sky130_fd_sc_hd__nand3_2 _30869_ (.A(_08837_),
    .B(_08431_),
    .C(_08840_),
    .Y(_08841_));
 sky130_fd_sc_hd__a21oi_2 _30870_ (.A1(_08833_),
    .A2(_08834_),
    .B1(_08429_),
    .Y(_08842_));
 sky130_fd_sc_hd__nand2_2 _30871_ (.A(_08833_),
    .B(_08834_),
    .Y(_08843_));
 sky130_fd_sc_hd__nor2_2 _30872_ (.A(_08435_),
    .B(_08843_),
    .Y(_08844_));
 sky130_fd_sc_hd__o22ai_2 _30873_ (.A1(_08842_),
    .A2(_08844_),
    .B1(_08784_),
    .B2(_08785_),
    .Y(_08845_));
 sky130_fd_sc_hd__nand2_2 _30874_ (.A(_08429_),
    .B(_08833_),
    .Y(_08846_));
 sky130_fd_sc_hd__o2111ai_2 _30875_ (.A1(_08831_),
    .A2(_08846_),
    .B1(_08832_),
    .C1(_08839_),
    .D1(_08838_),
    .Y(_08847_));
 sky130_fd_sc_hd__nand3_2 _30876_ (.A(_08845_),
    .B(_08847_),
    .C(_08439_),
    .Y(_08848_));
 sky130_fd_sc_hd__nand2_2 _30877_ (.A(_08841_),
    .B(_08848_),
    .Y(_08849_));
 sky130_fd_sc_hd__o21ai_2 _30878_ (.A1(_08709_),
    .A2(_08711_),
    .B1(_08849_),
    .Y(_08850_));
 sky130_fd_sc_hd__nand2_2 _30879_ (.A(_08708_),
    .B(_08706_),
    .Y(_08851_));
 sky130_fd_sc_hd__inv_2 _30880_ (.A(_08698_),
    .Y(_08852_));
 sky130_fd_sc_hd__nand2_2 _30881_ (.A(_08698_),
    .B(_08706_),
    .Y(_08853_));
 sky130_fd_sc_hd__nor2_2 _30882_ (.A(_08707_),
    .B(_08710_),
    .Y(_08854_));
 sky130_fd_sc_hd__nand2_2 _30883_ (.A(_08853_),
    .B(_08854_),
    .Y(_08855_));
 sky130_fd_sc_hd__o2111ai_2 _30884_ (.A1(_08851_),
    .A2(_08852_),
    .B1(_08848_),
    .C1(_08841_),
    .D1(_08855_),
    .Y(_08856_));
 sky130_fd_sc_hd__nand3_2 _30885_ (.A(_08595_),
    .B(_08850_),
    .C(_08856_),
    .Y(_08857_));
 sky130_fd_sc_hd__nor3_2 _30886_ (.A(_08258_),
    .B(_08436_),
    .C(_08439_),
    .Y(_08858_));
 sky130_fd_sc_hd__a31oi_2 _30887_ (.A1(_08541_),
    .A2(_08441_),
    .A3(_08547_),
    .B1(_08858_),
    .Y(_08859_));
 sky130_fd_sc_hd__o211ai_2 _30888_ (.A1(_08709_),
    .A2(_08711_),
    .B1(_08841_),
    .C1(_08848_),
    .Y(_08860_));
 sky130_fd_sc_hd__nand3_2 _30889_ (.A(_08698_),
    .B(_08708_),
    .C(_08706_),
    .Y(_08861_));
 sky130_fd_sc_hd__nand3_2 _30890_ (.A(_08849_),
    .B(_08855_),
    .C(_08861_),
    .Y(_08862_));
 sky130_fd_sc_hd__nand3_2 _30891_ (.A(_08859_),
    .B(_08860_),
    .C(_08862_),
    .Y(_08863_));
 sky130_fd_sc_hd__and2b_2 _30892_ (.A_N(_08520_),
    .B(_08514_),
    .X(_08864_));
 sky130_fd_sc_hd__a21oi_2 _30893_ (.A1(_08540_),
    .A2(_08534_),
    .B1(_08864_),
    .Y(_08865_));
 sky130_fd_sc_hd__and3_2 _30894_ (.A(_08540_),
    .B(_08534_),
    .C(_08864_),
    .X(_08866_));
 sky130_fd_sc_hd__nor2_2 _30895_ (.A(_08865_),
    .B(_08866_),
    .Y(_08867_));
 sky130_fd_sc_hd__inv_2 _30896_ (.A(_08867_),
    .Y(_08868_));
 sky130_fd_sc_hd__a21o_2 _30897_ (.A1(_08857_),
    .A2(_08863_),
    .B1(_08868_),
    .X(_08869_));
 sky130_fd_sc_hd__nand3_2 _30898_ (.A(_08441_),
    .B(_08547_),
    .C(_08433_),
    .Y(_08870_));
 sky130_fd_sc_hd__a2bb2oi_2 _30899_ (.A1_N(_08536_),
    .A2_N(_08870_),
    .B1(_08261_),
    .B2(_08304_),
    .Y(_08871_));
 sky130_fd_sc_hd__a22oi_2 _30900_ (.A1(_08871_),
    .A2(_08538_),
    .B1(_08549_),
    .B2(_08559_),
    .Y(_08872_));
 sky130_fd_sc_hd__nand3_2 _30901_ (.A(_08868_),
    .B(_08857_),
    .C(_08863_),
    .Y(_08873_));
 sky130_fd_sc_hd__nand3_2 _30902_ (.A(_08869_),
    .B(_08872_),
    .C(_08873_),
    .Y(_08874_));
 sky130_fd_sc_hd__nand2_2 _30903_ (.A(_08538_),
    .B(_08542_),
    .Y(_08875_));
 sky130_fd_sc_hd__nor2_2 _30904_ (.A(_08544_),
    .B(_08875_),
    .Y(_08876_));
 sky130_fd_sc_hd__a22oi_2 _30905_ (.A1(_08553_),
    .A2(_08554_),
    .B1(_08875_),
    .B2(_08544_),
    .Y(_08877_));
 sky130_fd_sc_hd__nand3_2 _30906_ (.A(_08857_),
    .B(_08863_),
    .C(_08867_),
    .Y(_08878_));
 sky130_fd_sc_hd__o2bb2ai_2 _30907_ (.A1_N(_08863_),
    .A2_N(_08857_),
    .B1(_08865_),
    .B2(_08866_),
    .Y(_08879_));
 sky130_fd_sc_hd__o211ai_2 _30908_ (.A1(_08876_),
    .A2(_08877_),
    .B1(_08878_),
    .C1(_08879_),
    .Y(_08880_));
 sky130_fd_sc_hd__nand2_2 _30909_ (.A(_08874_),
    .B(_08880_),
    .Y(_08881_));
 sky130_fd_sc_hd__inv_2 _30910_ (.A(_08551_),
    .Y(_08882_));
 sky130_fd_sc_hd__nor2_2 _30911_ (.A(_08552_),
    .B(_08882_),
    .Y(_08883_));
 sky130_fd_sc_hd__inv_2 _30912_ (.A(_08883_),
    .Y(_08884_));
 sky130_fd_sc_hd__nand2_2 _30913_ (.A(_08881_),
    .B(_08884_),
    .Y(_08885_));
 sky130_fd_sc_hd__nand3_2 _30914_ (.A(_08874_),
    .B(_08880_),
    .C(_08883_),
    .Y(_08886_));
 sky130_fd_sc_hd__nand3_2 _30915_ (.A(_08593_),
    .B(_08885_),
    .C(_08886_),
    .Y(_08887_));
 sky130_fd_sc_hd__nand2_2 _30916_ (.A(_08881_),
    .B(_08883_),
    .Y(_08888_));
 sky130_fd_sc_hd__a21oi_2 _30917_ (.A1(_08543_),
    .A2(_08549_),
    .B1(_08559_),
    .Y(_08889_));
 sky130_fd_sc_hd__and3_2 _30918_ (.A(_08270_),
    .B(_08272_),
    .C(_08273_),
    .X(_08890_));
 sky130_fd_sc_hd__a31oi_2 _30919_ (.A1(_08262_),
    .A2(_08266_),
    .A3(_08268_),
    .B1(_08285_),
    .Y(_08891_));
 sky130_fd_sc_hd__o21ai_2 _30920_ (.A1(_08890_),
    .A2(_08891_),
    .B1(_08560_),
    .Y(_08892_));
 sky130_fd_sc_hd__a2bb2oi_2 _30921_ (.A1_N(_08889_),
    .A2_N(_08892_),
    .B1(_08577_),
    .B2(_08567_),
    .Y(_08893_));
 sky130_fd_sc_hd__nand3_2 _30922_ (.A(_08874_),
    .B(_08880_),
    .C(_08884_),
    .Y(_08894_));
 sky130_fd_sc_hd__nand3_2 _30923_ (.A(_08888_),
    .B(_08893_),
    .C(_08894_),
    .Y(_08895_));
 sky130_fd_sc_hd__and2_2 _30924_ (.A(_08887_),
    .B(_08895_),
    .X(_08896_));
 sky130_fd_sc_hd__and2b_2 _30925_ (.A_N(_08591_),
    .B(_08579_),
    .X(_08897_));
 sky130_fd_sc_hd__xnor2_2 _30926_ (.A(_08896_),
    .B(_08897_),
    .Y(_02644_));
 sky130_fd_sc_hd__and2_2 _30927_ (.A(_08687_),
    .B(_08678_),
    .X(_08898_));
 sky130_fd_sc_hd__a21o_2 _30928_ (.A1(_08851_),
    .A2(_08698_),
    .B1(_08898_),
    .X(_08899_));
 sky130_fd_sc_hd__inv_2 _30929_ (.A(_08899_),
    .Y(_08900_));
 sky130_fd_sc_hd__and3_2 _30930_ (.A(_08851_),
    .B(_08698_),
    .C(_08898_),
    .X(_08901_));
 sky130_fd_sc_hd__nand2_2 _30931_ (.A(_06735_),
    .B(_08651_),
    .Y(_08902_));
 sky130_fd_sc_hd__nand2_2 _30932_ (.A(_05721_),
    .B(_08103_),
    .Y(_08903_));
 sky130_fd_sc_hd__nor2_2 _30933_ (.A(_08902_),
    .B(_08903_),
    .Y(_08904_));
 sky130_fd_sc_hd__buf_1 _30934_ (.A(\pcpi_mul.rs1[26] ),
    .X(_08905_));
 sky130_fd_sc_hd__nand2_2 _30935_ (.A(_06057_),
    .B(_08905_),
    .Y(_08906_));
 sky130_fd_sc_hd__inv_2 _30936_ (.A(_08906_),
    .Y(_08907_));
 sky130_fd_sc_hd__nand2_2 _30937_ (.A(_08902_),
    .B(_08903_),
    .Y(_08908_));
 sky130_fd_sc_hd__nand2_2 _30938_ (.A(_08907_),
    .B(_08908_),
    .Y(_08909_));
 sky130_fd_sc_hd__buf_1 _30939_ (.A(_08497_),
    .X(_08910_));
 sky130_fd_sc_hd__a22oi_2 _30940_ (.A1(_19389_),
    .A2(_19579_),
    .B1(_19392_),
    .B2(_08910_),
    .Y(_08911_));
 sky130_fd_sc_hd__o21ai_2 _30941_ (.A1(_08911_),
    .A2(_08904_),
    .B1(_08906_),
    .Y(_08912_));
 sky130_fd_sc_hd__a21o_2 _30942_ (.A1(_08647_),
    .A2(_08648_),
    .B1(_08653_),
    .X(_08913_));
 sky130_fd_sc_hd__o211ai_2 _30943_ (.A1(_08904_),
    .A2(_08909_),
    .B1(_08912_),
    .C1(_08913_),
    .Y(_08914_));
 sky130_fd_sc_hd__or2_2 _30944_ (.A(_08902_),
    .B(_08903_),
    .X(_08915_));
 sky130_fd_sc_hd__nand3_2 _30945_ (.A(_08915_),
    .B(_08908_),
    .C(_08906_),
    .Y(_08916_));
 sky130_fd_sc_hd__a21oi_2 _30946_ (.A1(_08647_),
    .A2(_08648_),
    .B1(_08653_),
    .Y(_08917_));
 sky130_fd_sc_hd__o21ai_2 _30947_ (.A1(_08911_),
    .A2(_08904_),
    .B1(_08907_),
    .Y(_08918_));
 sky130_fd_sc_hd__nand3_2 _30948_ (.A(_08916_),
    .B(_08917_),
    .C(_08918_),
    .Y(_08919_));
 sky130_fd_sc_hd__buf_1 _30949_ (.A(\pcpi_mul.rs1[25] ),
    .X(_08920_));
 sky130_fd_sc_hd__buf_1 _30950_ (.A(_08920_),
    .X(_08921_));
 sky130_fd_sc_hd__buf_1 _30951_ (.A(_08661_),
    .X(_08922_));
 sky130_fd_sc_hd__nand2_2 _30952_ (.A(_06219_),
    .B(_08922_),
    .Y(_08923_));
 sky130_fd_sc_hd__a21o_2 _30953_ (.A1(_19402_),
    .A2(_08921_),
    .B1(_08923_),
    .X(_08924_));
 sky130_fd_sc_hd__nand2_2 _30954_ (.A(_06220_),
    .B(_19565_),
    .Y(_08925_));
 sky130_fd_sc_hd__a21o_2 _30955_ (.A1(_19399_),
    .A2(_19568_),
    .B1(_08925_),
    .X(_08926_));
 sky130_fd_sc_hd__nand2_2 _30956_ (.A(_05116_),
    .B(_19572_),
    .Y(_08927_));
 sky130_fd_sc_hd__and3_2 _30957_ (.A(_08924_),
    .B(_08926_),
    .C(_08927_),
    .X(_08928_));
 sky130_fd_sc_hd__a21oi_2 _30958_ (.A1(_08924_),
    .A2(_08926_),
    .B1(_08927_),
    .Y(_08929_));
 sky130_fd_sc_hd__o2bb2ai_2 _30959_ (.A1_N(_08914_),
    .A2_N(_08919_),
    .B1(_08928_),
    .B2(_08929_),
    .Y(_08930_));
 sky130_fd_sc_hd__nor2_2 _30960_ (.A(_08929_),
    .B(_08928_),
    .Y(_08931_));
 sky130_fd_sc_hd__nand3_2 _30961_ (.A(_08931_),
    .B(_08919_),
    .C(_08914_),
    .Y(_08932_));
 sky130_fd_sc_hd__nand2_2 _30962_ (.A(_08676_),
    .B(_08659_),
    .Y(_08933_));
 sky130_fd_sc_hd__nand2_2 _30963_ (.A(_08933_),
    .B(_08655_),
    .Y(_08934_));
 sky130_fd_sc_hd__a21oi_2 _30964_ (.A1(_08930_),
    .A2(_08932_),
    .B1(_08934_),
    .Y(_08935_));
 sky130_fd_sc_hd__and3_2 _30965_ (.A(_08934_),
    .B(_08930_),
    .C(_08932_),
    .X(_08936_));
 sky130_fd_sc_hd__inv_2 _30966_ (.A(_08669_),
    .Y(_08937_));
 sky130_fd_sc_hd__nor2_2 _30967_ (.A(_08665_),
    .B(_08937_),
    .Y(_08938_));
 sky130_fd_sc_hd__inv_2 _30968_ (.A(_08938_),
    .Y(_08939_));
 sky130_fd_sc_hd__o21ai_2 _30969_ (.A1(_08935_),
    .A2(_08936_),
    .B1(_08939_),
    .Y(_08940_));
 sky130_fd_sc_hd__a21o_2 _30970_ (.A1(_08930_),
    .A2(_08932_),
    .B1(_08934_),
    .X(_08941_));
 sky130_fd_sc_hd__nand3_2 _30971_ (.A(_08934_),
    .B(_08932_),
    .C(_08930_),
    .Y(_08942_));
 sky130_fd_sc_hd__nand3_2 _30972_ (.A(_08941_),
    .B(_08938_),
    .C(_08942_),
    .Y(_08943_));
 sky130_fd_sc_hd__nand2_2 _30973_ (.A(_08940_),
    .B(_08943_),
    .Y(_08944_));
 sky130_fd_sc_hd__a22oi_2 _30974_ (.A1(_19381_),
    .A2(_19586_),
    .B1(_19384_),
    .B2(_19583_),
    .Y(_08945_));
 sky130_fd_sc_hd__inv_2 _30975_ (.A(\pcpi_mul.rs1[19] ),
    .Y(_08946_));
 sky130_fd_sc_hd__buf_1 _30976_ (.A(_08946_),
    .X(_08947_));
 sky130_fd_sc_hd__buf_1 _30977_ (.A(_05448_),
    .X(_08948_));
 sky130_fd_sc_hd__buf_1 _30978_ (.A(_05641_),
    .X(_08949_));
 sky130_fd_sc_hd__buf_1 _30979_ (.A(_08089_),
    .X(_08950_));
 sky130_fd_sc_hd__nand3_2 _30980_ (.A(_08948_),
    .B(_08949_),
    .C(_08950_),
    .Y(_08951_));
 sky130_fd_sc_hd__nor2_2 _30981_ (.A(_08947_),
    .B(_08951_),
    .Y(_08952_));
 sky130_fd_sc_hd__buf_1 _30982_ (.A(_06496_),
    .X(_08953_));
 sky130_fd_sc_hd__nand2_2 _30983_ (.A(_08953_),
    .B(_19580_),
    .Y(_08954_));
 sky130_fd_sc_hd__o21ai_2 _30984_ (.A1(_08945_),
    .A2(_08952_),
    .B1(_08954_),
    .Y(_08955_));
 sky130_fd_sc_hd__o21ai_2 _30985_ (.A1(_08756_),
    .A2(_08754_),
    .B1(_08760_),
    .Y(_08956_));
 sky130_fd_sc_hd__buf_1 _30986_ (.A(_08947_),
    .X(_08957_));
 sky130_fd_sc_hd__inv_2 _30987_ (.A(_08954_),
    .Y(_08958_));
 sky130_fd_sc_hd__buf_1 _30988_ (.A(_08596_),
    .X(_08959_));
 sky130_fd_sc_hd__a22o_2 _30989_ (.A1(_19381_),
    .A2(_08959_),
    .B1(_19384_),
    .B2(_07852_),
    .X(_08960_));
 sky130_fd_sc_hd__o211ai_2 _30990_ (.A1(_08957_),
    .A2(_08951_),
    .B1(_08958_),
    .C1(_08960_),
    .Y(_08961_));
 sky130_fd_sc_hd__nand3_2 _30991_ (.A(_08955_),
    .B(_08956_),
    .C(_08961_),
    .Y(_08962_));
 sky130_fd_sc_hd__o21ai_2 _30992_ (.A1(_08945_),
    .A2(_08952_),
    .B1(_08958_),
    .Y(_08963_));
 sky130_fd_sc_hd__a21oi_2 _30993_ (.A1(_08762_),
    .A2(_08757_),
    .B1(_08755_),
    .Y(_08964_));
 sky130_fd_sc_hd__o211ai_2 _30994_ (.A1(_08957_),
    .A2(_08951_),
    .B1(_08954_),
    .C1(_08960_),
    .Y(_08965_));
 sky130_fd_sc_hd__nand3_2 _30995_ (.A(_08963_),
    .B(_08964_),
    .C(_08965_),
    .Y(_08966_));
 sky130_fd_sc_hd__nor2_2 _30996_ (.A(_08605_),
    .B(_08600_),
    .Y(_08967_));
 sky130_fd_sc_hd__o2bb2ai_2 _30997_ (.A1_N(_08962_),
    .A2_N(_08966_),
    .B1(_08597_),
    .B2(_08967_),
    .Y(_08968_));
 sky130_fd_sc_hd__nor2_2 _30998_ (.A(_08597_),
    .B(_08967_),
    .Y(_08969_));
 sky130_fd_sc_hd__nand3_2 _30999_ (.A(_08966_),
    .B(_08962_),
    .C(_08969_),
    .Y(_08970_));
 sky130_fd_sc_hd__nand2_2 _31000_ (.A(_08752_),
    .B(_08764_),
    .Y(_08971_));
 sky130_fd_sc_hd__nand2_2 _31001_ (.A(_08971_),
    .B(_08746_),
    .Y(_08972_));
 sky130_fd_sc_hd__a21oi_2 _31002_ (.A1(_08968_),
    .A2(_08970_),
    .B1(_08972_),
    .Y(_08973_));
 sky130_fd_sc_hd__nand2_2 _31003_ (.A(_08966_),
    .B(_08969_),
    .Y(_08974_));
 sky130_fd_sc_hd__inv_2 _31004_ (.A(_08962_),
    .Y(_08975_));
 sky130_fd_sc_hd__o211a_2 _31005_ (.A1(_08974_),
    .A2(_08975_),
    .B1(_08968_),
    .C1(_08972_),
    .X(_08976_));
 sky130_fd_sc_hd__nand2_2 _31006_ (.A(_08621_),
    .B(_08608_),
    .Y(_08977_));
 sky130_fd_sc_hd__inv_2 _31007_ (.A(_08977_),
    .Y(_08978_));
 sky130_fd_sc_hd__o21ai_2 _31008_ (.A1(_08973_),
    .A2(_08976_),
    .B1(_08978_),
    .Y(_08979_));
 sky130_fd_sc_hd__a21o_2 _31009_ (.A1(_08968_),
    .A2(_08970_),
    .B1(_08972_),
    .X(_08980_));
 sky130_fd_sc_hd__nand3_2 _31010_ (.A(_08972_),
    .B(_08968_),
    .C(_08970_),
    .Y(_08981_));
 sky130_fd_sc_hd__nand3_2 _31011_ (.A(_08980_),
    .B(_08981_),
    .C(_08977_),
    .Y(_08982_));
 sky130_fd_sc_hd__o21ai_2 _31012_ (.A1(_08630_),
    .A2(_08620_),
    .B1(_08629_),
    .Y(_08983_));
 sky130_fd_sc_hd__nand3_2 _31013_ (.A(_08979_),
    .B(_08982_),
    .C(_08983_),
    .Y(_08984_));
 sky130_fd_sc_hd__o21ai_2 _31014_ (.A1(_08973_),
    .A2(_08976_),
    .B1(_08977_),
    .Y(_08985_));
 sky130_fd_sc_hd__nand3_2 _31015_ (.A(_08980_),
    .B(_08981_),
    .C(_08978_),
    .Y(_08986_));
 sky130_fd_sc_hd__nand2_2 _31016_ (.A(_08629_),
    .B(_08630_),
    .Y(_08987_));
 sky130_fd_sc_hd__nand2_2 _31017_ (.A(_08987_),
    .B(_08628_),
    .Y(_08988_));
 sky130_fd_sc_hd__nand3_2 _31018_ (.A(_08985_),
    .B(_08986_),
    .C(_08988_),
    .Y(_08989_));
 sky130_fd_sc_hd__nand3_2 _31019_ (.A(_08944_),
    .B(_08984_),
    .C(_08989_),
    .Y(_08990_));
 sky130_fd_sc_hd__a21oi_2 _31020_ (.A1(_08941_),
    .A2(_08942_),
    .B1(_08939_),
    .Y(_08991_));
 sky130_fd_sc_hd__and3_2 _31021_ (.A(_08941_),
    .B(_08939_),
    .C(_08942_),
    .X(_08992_));
 sky130_fd_sc_hd__o2bb2ai_2 _31022_ (.A1_N(_08984_),
    .A2_N(_08989_),
    .B1(_08991_),
    .B2(_08992_),
    .Y(_08993_));
 sky130_fd_sc_hd__inv_2 _31023_ (.A(_08776_),
    .Y(_08994_));
 sky130_fd_sc_hd__a21oi_2 _31024_ (.A1(_08364_),
    .A2(_08367_),
    .B1(_08362_),
    .Y(_08995_));
 sky130_fd_sc_hd__and2_2 _31025_ (.A(_08782_),
    .B(_08995_),
    .X(_08996_));
 sky130_fd_sc_hd__o2bb2ai_2 _31026_ (.A1_N(_08990_),
    .A2_N(_08993_),
    .B1(_08994_),
    .B2(_08996_),
    .Y(_08997_));
 sky130_fd_sc_hd__and3_2 _31027_ (.A(_08779_),
    .B(_08781_),
    .C(_08780_),
    .X(_08998_));
 sky130_fd_sc_hd__a31oi_2 _31028_ (.A1(_08769_),
    .A2(_08775_),
    .A3(_08422_),
    .B1(_08995_),
    .Y(_08999_));
 sky130_fd_sc_hd__o211ai_2 _31029_ (.A1(_08998_),
    .A2(_08999_),
    .B1(_08990_),
    .C1(_08993_),
    .Y(_09000_));
 sky130_fd_sc_hd__a21bo_2 _31030_ (.A1(_08632_),
    .A2(_08695_),
    .B1_N(_08638_),
    .X(_09001_));
 sky130_fd_sc_hd__nand3_2 _31031_ (.A(_08997_),
    .B(_09000_),
    .C(_09001_),
    .Y(_09002_));
 sky130_fd_sc_hd__nand2_2 _31032_ (.A(_08782_),
    .B(_08995_),
    .Y(_09003_));
 sky130_fd_sc_hd__a22oi_2 _31033_ (.A1(_08776_),
    .A2(_09003_),
    .B1(_08993_),
    .B2(_08990_),
    .Y(_09004_));
 sky130_fd_sc_hd__o211a_2 _31034_ (.A1(_08998_),
    .A2(_08999_),
    .B1(_08990_),
    .C1(_08993_),
    .X(_09005_));
 sky130_fd_sc_hd__o21bai_2 _31035_ (.A1(_09004_),
    .A2(_09005_),
    .B1_N(_09001_),
    .Y(_09006_));
 sky130_fd_sc_hd__nand2_2 _31036_ (.A(_08725_),
    .B(_08733_),
    .Y(_09007_));
 sky130_fd_sc_hd__buf_1 _31037_ (.A(_19354_),
    .X(_09008_));
 sky130_fd_sc_hd__buf_1 _31038_ (.A(_07417_),
    .X(_09009_));
 sky130_fd_sc_hd__buf_1 _31039_ (.A(_05598_),
    .X(_09010_));
 sky130_fd_sc_hd__a22oi_2 _31040_ (.A1(_09008_),
    .A2(_19614_),
    .B1(_09009_),
    .B2(_09010_),
    .Y(_09011_));
 sky130_fd_sc_hd__buf_1 _31041_ (.A(_06694_),
    .X(_09012_));
 sky130_fd_sc_hd__nand3_2 _31042_ (.A(_07898_),
    .B(_19357_),
    .C(_07210_),
    .Y(_09013_));
 sky130_fd_sc_hd__nor2_2 _31043_ (.A(_09012_),
    .B(_09013_),
    .Y(_09014_));
 sky130_fd_sc_hd__nand2_2 _31044_ (.A(_19359_),
    .B(_06369_),
    .Y(_09015_));
 sky130_fd_sc_hd__o21ai_2 _31045_ (.A1(_09011_),
    .A2(_09014_),
    .B1(_09015_),
    .Y(_09016_));
 sky130_fd_sc_hd__inv_2 _31046_ (.A(_09015_),
    .Y(_09017_));
 sky130_fd_sc_hd__buf_1 _31047_ (.A(_07236_),
    .X(_09018_));
 sky130_fd_sc_hd__buf_1 _31048_ (.A(_06823_),
    .X(_09019_));
 sky130_fd_sc_hd__a22o_2 _31049_ (.A1(_09018_),
    .A2(_05737_),
    .B1(_09019_),
    .B2(_05738_),
    .X(_09020_));
 sky130_fd_sc_hd__o211ai_2 _31050_ (.A1(_09012_),
    .A2(_09013_),
    .B1(_09017_),
    .C1(_09020_),
    .Y(_09021_));
 sky130_fd_sc_hd__o21ai_2 _31051_ (.A1(_08814_),
    .A2(_08810_),
    .B1(_08817_),
    .Y(_09022_));
 sky130_fd_sc_hd__nand3_2 _31052_ (.A(_09016_),
    .B(_09021_),
    .C(_09022_),
    .Y(_09023_));
 sky130_fd_sc_hd__o21ai_2 _31053_ (.A1(_09011_),
    .A2(_09014_),
    .B1(_09017_),
    .Y(_09024_));
 sky130_fd_sc_hd__o21ai_2 _31054_ (.A1(_08811_),
    .A2(_08812_),
    .B1(_08814_),
    .Y(_09025_));
 sky130_fd_sc_hd__nand2_2 _31055_ (.A(_09025_),
    .B(_08818_),
    .Y(_09026_));
 sky130_fd_sc_hd__o211ai_2 _31056_ (.A1(_09012_),
    .A2(_09013_),
    .B1(_09015_),
    .C1(_09020_),
    .Y(_09027_));
 sky130_fd_sc_hd__nand3_2 _31057_ (.A(_09024_),
    .B(_09026_),
    .C(_09027_),
    .Y(_09028_));
 sky130_fd_sc_hd__nor2_2 _31058_ (.A(_08716_),
    .B(_08714_),
    .Y(_09029_));
 sky130_fd_sc_hd__o2bb2ai_2 _31059_ (.A1_N(_09023_),
    .A2_N(_09028_),
    .B1(_08712_),
    .B2(_09029_),
    .Y(_09030_));
 sky130_fd_sc_hd__nor2_2 _31060_ (.A(_08712_),
    .B(_09029_),
    .Y(_09031_));
 sky130_fd_sc_hd__nand3_2 _31061_ (.A(_09023_),
    .B(_09028_),
    .C(_09031_),
    .Y(_09032_));
 sky130_fd_sc_hd__a22oi_2 _31062_ (.A1(_08721_),
    .A2(_09007_),
    .B1(_09030_),
    .B2(_09032_),
    .Y(_09033_));
 sky130_fd_sc_hd__and3_2 _31063_ (.A(_08722_),
    .B(_08723_),
    .C(_08724_),
    .X(_09034_));
 sky130_fd_sc_hd__a31oi_2 _31064_ (.A1(_08717_),
    .A2(_08718_),
    .A3(_08720_),
    .B1(_08733_),
    .Y(_09035_));
 sky130_fd_sc_hd__o211a_2 _31065_ (.A1(_09034_),
    .A2(_09035_),
    .B1(_09032_),
    .C1(_09030_),
    .X(_09036_));
 sky130_fd_sc_hd__a22oi_2 _31066_ (.A1(_08315_),
    .A2(_19603_),
    .B1(_08320_),
    .B2(_06059_),
    .Y(_09037_));
 sky130_fd_sc_hd__and4_2 _31067_ (.A(_08315_),
    .B(_06276_),
    .C(_06724_),
    .D(_06538_),
    .X(_09038_));
 sky130_fd_sc_hd__nand2_2 _31068_ (.A(_06446_),
    .B(_06206_),
    .Y(_09039_));
 sky130_fd_sc_hd__inv_2 _31069_ (.A(_09039_),
    .Y(_09040_));
 sky130_fd_sc_hd__o21ai_2 _31070_ (.A1(_09037_),
    .A2(_09038_),
    .B1(_09040_),
    .Y(_09041_));
 sky130_fd_sc_hd__nand2_2 _31071_ (.A(_07012_),
    .B(_07939_),
    .Y(_09042_));
 sky130_fd_sc_hd__nand3b_2 _31072_ (.A_N(_09042_),
    .B(_06115_),
    .C(_06736_),
    .Y(_09043_));
 sky130_fd_sc_hd__a22o_2 _31073_ (.A1(_08315_),
    .A2(_06726_),
    .B1(_07934_),
    .B2(_06059_),
    .X(_09044_));
 sky130_fd_sc_hd__nand3_2 _31074_ (.A(_09043_),
    .B(_09039_),
    .C(_09044_),
    .Y(_09045_));
 sky130_fd_sc_hd__nand2_2 _31075_ (.A(_09041_),
    .B(_09045_),
    .Y(_09046_));
 sky130_fd_sc_hd__nand2_2 _31076_ (.A(_08742_),
    .B(_08749_),
    .Y(_09047_));
 sky130_fd_sc_hd__nand2_2 _31077_ (.A(_09046_),
    .B(_09047_),
    .Y(_09048_));
 sky130_fd_sc_hd__o2111ai_2 _31078_ (.A1(_08740_),
    .A2(_08743_),
    .B1(_08749_),
    .C1(_09045_),
    .D1(_09041_),
    .Y(_09049_));
 sky130_fd_sc_hd__a22oi_2 _31079_ (.A1(_05801_),
    .A2(_07798_),
    .B1(_08331_),
    .B2(_06950_),
    .Y(_09050_));
 sky130_fd_sc_hd__buf_1 _31080_ (.A(_06430_),
    .X(_09051_));
 sky130_fd_sc_hd__and4_2 _31081_ (.A(_09051_),
    .B(_06433_),
    .C(_19590_),
    .D(_06748_),
    .X(_09052_));
 sky130_fd_sc_hd__nand2_2 _31082_ (.A(_19376_),
    .B(_08447_),
    .Y(_09053_));
 sky130_fd_sc_hd__o21bai_2 _31083_ (.A1(_09050_),
    .A2(_09052_),
    .B1_N(_09053_),
    .Y(_09054_));
 sky130_fd_sc_hd__inv_2 _31084_ (.A(_09054_),
    .Y(_09055_));
 sky130_fd_sc_hd__nand2_2 _31085_ (.A(_06256_),
    .B(_06560_),
    .Y(_09056_));
 sky130_fd_sc_hd__nand3b_2 _31086_ (.A_N(_09056_),
    .B(_05808_),
    .C(_06750_),
    .Y(_09057_));
 sky130_fd_sc_hd__a22o_2 _31087_ (.A1(_05801_),
    .A2(_07798_),
    .B1(_08331_),
    .B2(_06950_),
    .X(_09058_));
 sky130_fd_sc_hd__nand3_2 _31088_ (.A(_09057_),
    .B(_09053_),
    .C(_09058_),
    .Y(_09059_));
 sky130_fd_sc_hd__inv_2 _31089_ (.A(_09059_),
    .Y(_09060_));
 sky130_fd_sc_hd__o2bb2ai_2 _31090_ (.A1_N(_09048_),
    .A2_N(_09049_),
    .B1(_09055_),
    .B2(_09060_),
    .Y(_09061_));
 sky130_fd_sc_hd__nand2_2 _31091_ (.A(_09054_),
    .B(_09059_),
    .Y(_09062_));
 sky130_fd_sc_hd__inv_2 _31092_ (.A(_09062_),
    .Y(_09063_));
 sky130_fd_sc_hd__nand3_2 _31093_ (.A(_09063_),
    .B(_09048_),
    .C(_09049_),
    .Y(_09064_));
 sky130_fd_sc_hd__nand2_2 _31094_ (.A(_09061_),
    .B(_09064_),
    .Y(_09065_));
 sky130_fd_sc_hd__o21ai_2 _31095_ (.A1(_09033_),
    .A2(_09036_),
    .B1(_09065_),
    .Y(_09066_));
 sky130_fd_sc_hd__a21oi_2 _31096_ (.A1(_09048_),
    .A2(_09049_),
    .B1(_09062_),
    .Y(_09067_));
 sky130_fd_sc_hd__nand3_2 _31097_ (.A(_09048_),
    .B(_09062_),
    .C(_09049_),
    .Y(_09068_));
 sky130_fd_sc_hd__inv_2 _31098_ (.A(_09068_),
    .Y(_09069_));
 sky130_fd_sc_hd__o211ai_2 _31099_ (.A1(_09034_),
    .A2(_09035_),
    .B1(_09032_),
    .C1(_09030_),
    .Y(_09070_));
 sky130_fd_sc_hd__nand2_2 _31100_ (.A(_09030_),
    .B(_09032_),
    .Y(_09071_));
 sky130_fd_sc_hd__nand2_2 _31101_ (.A(_09007_),
    .B(_08721_),
    .Y(_09072_));
 sky130_fd_sc_hd__nand2_2 _31102_ (.A(_09071_),
    .B(_09072_),
    .Y(_09073_));
 sky130_fd_sc_hd__o211ai_2 _31103_ (.A1(_09067_),
    .A2(_09069_),
    .B1(_09070_),
    .C1(_09073_),
    .Y(_09074_));
 sky130_fd_sc_hd__nand3_2 _31104_ (.A(_09066_),
    .B(_09074_),
    .C(_08826_),
    .Y(_09075_));
 sky130_fd_sc_hd__o22ai_2 _31105_ (.A1(_09067_),
    .A2(_09069_),
    .B1(_09033_),
    .B2(_09036_),
    .Y(_09076_));
 sky130_fd_sc_hd__nand3_2 _31106_ (.A(_09073_),
    .B(_09065_),
    .C(_09070_),
    .Y(_09077_));
 sky130_fd_sc_hd__nand3_2 _31107_ (.A(_09076_),
    .B(_08830_),
    .C(_09077_),
    .Y(_09078_));
 sky130_fd_sc_hd__nor2_2 _31108_ (.A(_08768_),
    .B(_08731_),
    .Y(_09079_));
 sky130_fd_sc_hd__nor2_2 _31109_ (.A(_08737_),
    .B(_09079_),
    .Y(_09080_));
 sky130_fd_sc_hd__nand3_2 _31110_ (.A(_09075_),
    .B(_09078_),
    .C(_09080_),
    .Y(_09081_));
 sky130_fd_sc_hd__o2bb2ai_2 _31111_ (.A1_N(_09078_),
    .A2_N(_09075_),
    .B1(_08737_),
    .B2(_09079_),
    .Y(_09082_));
 sky130_fd_sc_hd__nor2_2 _31112_ (.A(_08828_),
    .B(_08829_),
    .Y(_09083_));
 sky130_fd_sc_hd__and4_2 _31113_ (.A(_08396_),
    .B(_08386_),
    .C(_06629_),
    .D(_05330_),
    .X(_09084_));
 sky130_fd_sc_hd__a22o_2 _31114_ (.A1(_08396_),
    .A2(_05204_),
    .B1(_08383_),
    .B2(_06501_),
    .X(_09085_));
 sky130_fd_sc_hd__nand2_2 _31115_ (.A(_08388_),
    .B(_05184_),
    .Y(_09086_));
 sky130_fd_sc_hd__inv_2 _31116_ (.A(_09086_),
    .Y(_09087_));
 sky130_fd_sc_hd__nand2_2 _31117_ (.A(_09085_),
    .B(_09087_),
    .Y(_09088_));
 sky130_fd_sc_hd__o21ai_2 _31118_ (.A1(_08794_),
    .A2(_08792_),
    .B1(_08800_),
    .Y(_09089_));
 sky130_fd_sc_hd__a22oi_2 _31119_ (.A1(_08385_),
    .A2(_05330_),
    .B1(_07974_),
    .B2(_06629_),
    .Y(_09090_));
 sky130_fd_sc_hd__o21ai_2 _31120_ (.A1(_09090_),
    .A2(_09084_),
    .B1(_09086_),
    .Y(_09091_));
 sky130_fd_sc_hd__o211ai_2 _31121_ (.A1(_09084_),
    .A2(_09088_),
    .B1(_09089_),
    .C1(_09091_),
    .Y(_09092_));
 sky130_fd_sc_hd__o21ai_2 _31122_ (.A1(_09090_),
    .A2(_09084_),
    .B1(_09087_),
    .Y(_09093_));
 sky130_fd_sc_hd__buf_1 _31123_ (.A(\pcpi_mul.rs2[23] ),
    .X(_09094_));
 sky130_fd_sc_hd__nand2_2 _31124_ (.A(_09094_),
    .B(_06447_),
    .Y(_09095_));
 sky130_fd_sc_hd__nand3b_2 _31125_ (.A_N(_09095_),
    .B(_19340_),
    .C(_05207_),
    .Y(_09096_));
 sky130_fd_sc_hd__nand3_2 _31126_ (.A(_09096_),
    .B(_09086_),
    .C(_09085_),
    .Y(_09097_));
 sky130_fd_sc_hd__nand3b_2 _31127_ (.A_N(_09089_),
    .B(_09093_),
    .C(_09097_),
    .Y(_09098_));
 sky130_fd_sc_hd__nand2_2 _31128_ (.A(_07894_),
    .B(_06606_),
    .Y(_09099_));
 sky130_fd_sc_hd__nand3b_2 _31129_ (.A_N(_09099_),
    .B(_08809_),
    .C(_05713_),
    .Y(_09100_));
 sky130_fd_sc_hd__buf_1 _31130_ (.A(_07480_),
    .X(_09101_));
 sky130_fd_sc_hd__a22o_2 _31131_ (.A1(_09101_),
    .A2(_05343_),
    .B1(_08185_),
    .B2(_05421_),
    .X(_09102_));
 sky130_fd_sc_hd__nand2_2 _31132_ (.A(_07475_),
    .B(_06507_),
    .Y(_09103_));
 sky130_fd_sc_hd__inv_2 _31133_ (.A(_09103_),
    .Y(_09104_));
 sky130_fd_sc_hd__a21oi_2 _31134_ (.A1(_09100_),
    .A2(_09102_),
    .B1(_09104_),
    .Y(_09105_));
 sky130_fd_sc_hd__and3_2 _31135_ (.A(_09100_),
    .B(_09102_),
    .C(_09104_),
    .X(_09106_));
 sky130_fd_sc_hd__nor2_2 _31136_ (.A(_09105_),
    .B(_09106_),
    .Y(_09107_));
 sky130_fd_sc_hd__a21o_2 _31137_ (.A1(_09092_),
    .A2(_09098_),
    .B1(_09107_),
    .X(_09108_));
 sky130_fd_sc_hd__nand2_2 _31138_ (.A(_08803_),
    .B(_08820_),
    .Y(_09109_));
 sky130_fd_sc_hd__nand2_2 _31139_ (.A(_09109_),
    .B(_08807_),
    .Y(_09110_));
 sky130_fd_sc_hd__nand3_2 _31140_ (.A(_09107_),
    .B(_09092_),
    .C(_09098_),
    .Y(_09111_));
 sky130_fd_sc_hd__nand3_2 _31141_ (.A(_09108_),
    .B(_09110_),
    .C(_09111_),
    .Y(_09112_));
 sky130_fd_sc_hd__inv_2 _31142_ (.A(_08803_),
    .Y(_09113_));
 sky130_fd_sc_hd__and3_2 _31143_ (.A(_08807_),
    .B(_08815_),
    .C(_08819_),
    .X(_09114_));
 sky130_fd_sc_hd__a2bb2oi_2 _31144_ (.A1_N(_09105_),
    .A2_N(_09106_),
    .B1(_09092_),
    .B2(_09098_),
    .Y(_09115_));
 sky130_fd_sc_hd__a21oi_2 _31145_ (.A1(_09100_),
    .A2(_09102_),
    .B1(_09103_),
    .Y(_09116_));
 sky130_fd_sc_hd__and3_2 _31146_ (.A(_09100_),
    .B(_09102_),
    .C(_09103_),
    .X(_09117_));
 sky130_fd_sc_hd__o211a_2 _31147_ (.A1(_09116_),
    .A2(_09117_),
    .B1(_09092_),
    .C1(_09098_),
    .X(_09118_));
 sky130_fd_sc_hd__o22ai_2 _31148_ (.A1(_09113_),
    .A2(_09114_),
    .B1(_09115_),
    .B2(_09118_),
    .Y(_09119_));
 sky130_fd_sc_hd__buf_2 _31149_ (.A(\pcpi_mul.rs2[25] ),
    .X(_09120_));
 sky130_fd_sc_hd__nand2_2 _31150_ (.A(_09120_),
    .B(_05543_),
    .Y(_09121_));
 sky130_fd_sc_hd__nand2_2 _31151_ (.A(_19327_),
    .B(_05188_),
    .Y(_09122_));
 sky130_fd_sc_hd__nor2_2 _31152_ (.A(_09121_),
    .B(_09122_),
    .Y(_09123_));
 sky130_fd_sc_hd__and2_2 _31153_ (.A(_09121_),
    .B(_09122_),
    .X(_09124_));
 sky130_fd_sc_hd__nor2_2 _31154_ (.A(_08423_),
    .B(_05101_),
    .Y(_09125_));
 sky130_fd_sc_hd__o21bai_2 _31155_ (.A1(_09123_),
    .A2(_09124_),
    .B1_N(_09125_),
    .Y(_09126_));
 sky130_fd_sc_hd__nand2_2 _31156_ (.A(_09121_),
    .B(_09122_),
    .Y(_09127_));
 sky130_fd_sc_hd__nand3b_2 _31157_ (.A_N(_09123_),
    .B(_09127_),
    .C(_09125_),
    .Y(_09128_));
 sky130_fd_sc_hd__and3_2 _31158_ (.A(_09126_),
    .B(_09128_),
    .C(_08787_),
    .X(_09129_));
 sky130_fd_sc_hd__and2_2 _31159_ (.A(_09126_),
    .B(_09128_),
    .X(_09130_));
 sky130_fd_sc_hd__nor2_2 _31160_ (.A(_08787_),
    .B(_09130_),
    .Y(_09131_));
 sky130_fd_sc_hd__o2bb2ai_2 _31161_ (.A1_N(_09112_),
    .A2_N(_09119_),
    .B1(_09129_),
    .B2(_09131_),
    .Y(_09132_));
 sky130_fd_sc_hd__nor2_2 _31162_ (.A(_09129_),
    .B(_09131_),
    .Y(_09133_));
 sky130_fd_sc_hd__nand3_2 _31163_ (.A(_09119_),
    .B(_09112_),
    .C(_09133_),
    .Y(_09134_));
 sky130_fd_sc_hd__a22oi_2 _31164_ (.A1(_09083_),
    .A2(_08826_),
    .B1(_09132_),
    .B2(_09134_),
    .Y(_09135_));
 sky130_fd_sc_hd__nand3_2 _31165_ (.A(_08831_),
    .B(_09132_),
    .C(_09134_),
    .Y(_09136_));
 sky130_fd_sc_hd__inv_2 _31166_ (.A(_09136_),
    .Y(_09137_));
 sky130_fd_sc_hd__o2bb2ai_2 _31167_ (.A1_N(_09081_),
    .A2_N(_09082_),
    .B1(_09135_),
    .B2(_09137_),
    .Y(_09138_));
 sky130_fd_sc_hd__and3_2 _31168_ (.A(_09119_),
    .B(_09112_),
    .C(_09133_),
    .X(_09139_));
 sky130_fd_sc_hd__nand2_2 _31169_ (.A(_08831_),
    .B(_09132_),
    .Y(_09140_));
 sky130_fd_sc_hd__a21oi_2 _31170_ (.A1(_09119_),
    .A2(_09112_),
    .B1(_09133_),
    .Y(_09141_));
 sky130_fd_sc_hd__o21ai_2 _31171_ (.A1(_09141_),
    .A2(_09139_),
    .B1(_08834_),
    .Y(_09142_));
 sky130_fd_sc_hd__o2111ai_2 _31172_ (.A1(_09139_),
    .A2(_09140_),
    .B1(_09142_),
    .C1(_09081_),
    .D1(_09082_),
    .Y(_09143_));
 sky130_fd_sc_hd__nand2_2 _31173_ (.A(_08839_),
    .B(_08832_),
    .Y(_09144_));
 sky130_fd_sc_hd__o22ai_2 _31174_ (.A1(_08435_),
    .A2(_08843_),
    .B1(_08784_),
    .B2(_09144_),
    .Y(_09145_));
 sky130_fd_sc_hd__a21oi_2 _31175_ (.A1(_09138_),
    .A2(_09143_),
    .B1(_09145_),
    .Y(_09146_));
 sky130_fd_sc_hd__a21oi_2 _31176_ (.A1(_09075_),
    .A2(_09078_),
    .B1(_09080_),
    .Y(_09147_));
 sky130_fd_sc_hd__nand3_2 _31177_ (.A(_09081_),
    .B(_09142_),
    .C(_09136_),
    .Y(_09148_));
 sky130_fd_sc_hd__o211a_2 _31178_ (.A1(_09147_),
    .A2(_09148_),
    .B1(_09138_),
    .C1(_09145_),
    .X(_09149_));
 sky130_fd_sc_hd__o2bb2ai_2 _31179_ (.A1_N(_09002_),
    .A2_N(_09006_),
    .B1(_09146_),
    .B2(_09149_),
    .Y(_09150_));
 sky130_fd_sc_hd__nand2_2 _31180_ (.A(_08997_),
    .B(_09001_),
    .Y(_09151_));
 sky130_fd_sc_hd__a22oi_2 _31181_ (.A1(_09142_),
    .A2(_09136_),
    .B1(_09082_),
    .B2(_09081_),
    .Y(_09152_));
 sky130_fd_sc_hd__nor2_2 _31182_ (.A(_09147_),
    .B(_09148_),
    .Y(_09153_));
 sky130_fd_sc_hd__a31oi_2 _31183_ (.A1(_08838_),
    .A2(_08832_),
    .A3(_08839_),
    .B1(_08844_),
    .Y(_09154_));
 sky130_fd_sc_hd__o21ai_2 _31184_ (.A1(_09152_),
    .A2(_09153_),
    .B1(_09154_),
    .Y(_09155_));
 sky130_fd_sc_hd__nand3_2 _31185_ (.A(_09145_),
    .B(_09138_),
    .C(_09143_),
    .Y(_09156_));
 sky130_fd_sc_hd__o2111ai_2 _31186_ (.A1(_09005_),
    .A2(_09151_),
    .B1(_09155_),
    .C1(_09156_),
    .D1(_09006_),
    .Y(_09157_));
 sky130_fd_sc_hd__a21oi_2 _31187_ (.A1(_08837_),
    .A2(_08840_),
    .B1(_08431_),
    .Y(_09158_));
 sky130_fd_sc_hd__a31o_2 _31188_ (.A1(_08855_),
    .A2(_08841_),
    .A3(_08861_),
    .B1(_09158_),
    .X(_09159_));
 sky130_fd_sc_hd__a21oi_2 _31189_ (.A1(_09150_),
    .A2(_09157_),
    .B1(_09159_),
    .Y(_09160_));
 sky130_fd_sc_hd__a31oi_2 _31190_ (.A1(_08855_),
    .A2(_08841_),
    .A3(_08861_),
    .B1(_09158_),
    .Y(_09161_));
 sky130_fd_sc_hd__a22oi_2 _31191_ (.A1(_09155_),
    .A2(_09156_),
    .B1(_09006_),
    .B2(_09002_),
    .Y(_09162_));
 sky130_fd_sc_hd__o2111a_2 _31192_ (.A1(_09005_),
    .A2(_09151_),
    .B1(_09155_),
    .C1(_09156_),
    .D1(_09006_),
    .X(_09163_));
 sky130_fd_sc_hd__nor3_2 _31193_ (.A(_09161_),
    .B(_09162_),
    .C(_09163_),
    .Y(_09164_));
 sky130_fd_sc_hd__o22ai_2 _31194_ (.A1(_08900_),
    .A2(_08901_),
    .B1(_09160_),
    .B2(_09164_),
    .Y(_09165_));
 sky130_fd_sc_hd__o21ai_2 _31195_ (.A1(_09162_),
    .A2(_09163_),
    .B1(_09161_),
    .Y(_09166_));
 sky130_fd_sc_hd__nand3_2 _31196_ (.A(_09159_),
    .B(_09150_),
    .C(_09157_),
    .Y(_09167_));
 sky130_fd_sc_hd__nor2_2 _31197_ (.A(_08901_),
    .B(_08900_),
    .Y(_09168_));
 sky130_fd_sc_hd__nand3_2 _31198_ (.A(_09166_),
    .B(_09167_),
    .C(_09168_),
    .Y(_09169_));
 sky130_fd_sc_hd__nand2_2 _31199_ (.A(_08863_),
    .B(_08867_),
    .Y(_09170_));
 sky130_fd_sc_hd__nand2_2 _31200_ (.A(_09170_),
    .B(_08857_),
    .Y(_09171_));
 sky130_fd_sc_hd__nand3_2 _31201_ (.A(_09165_),
    .B(_09169_),
    .C(_09171_),
    .Y(_09172_));
 sky130_fd_sc_hd__o21ai_2 _31202_ (.A1(_09160_),
    .A2(_09164_),
    .B1(_09168_),
    .Y(_09173_));
 sky130_fd_sc_hd__a21boi_2 _31203_ (.A1(_08863_),
    .A2(_08867_),
    .B1_N(_08857_),
    .Y(_09174_));
 sky130_fd_sc_hd__or2b_2 _31204_ (.A(_08901_),
    .B_N(_08899_),
    .X(_09175_));
 sky130_fd_sc_hd__nand3_2 _31205_ (.A(_09166_),
    .B(_09167_),
    .C(_09175_),
    .Y(_09176_));
 sky130_fd_sc_hd__nand3_2 _31206_ (.A(_09173_),
    .B(_09174_),
    .C(_09176_),
    .Y(_09177_));
 sky130_fd_sc_hd__nor2_2 _31207_ (.A(_08539_),
    .B(_08537_),
    .Y(_09178_));
 sky130_fd_sc_hd__o2bb2ai_2 _31208_ (.A1_N(_09172_),
    .A2_N(_09177_),
    .B1(_09178_),
    .B2(_08864_),
    .Y(_09179_));
 sky130_fd_sc_hd__nand3_2 _31209_ (.A(_09177_),
    .B(_09172_),
    .C(_08865_),
    .Y(_09180_));
 sky130_fd_sc_hd__nand2_2 _31210_ (.A(_08874_),
    .B(_08883_),
    .Y(_09181_));
 sky130_fd_sc_hd__nand2_2 _31211_ (.A(_09181_),
    .B(_08880_),
    .Y(_09182_));
 sky130_fd_sc_hd__a21oi_2 _31212_ (.A1(_09179_),
    .A2(_09180_),
    .B1(_09182_),
    .Y(_09183_));
 sky130_fd_sc_hd__and3_2 _31213_ (.A(_09165_),
    .B(_09169_),
    .C(_09171_),
    .X(_09184_));
 sky130_fd_sc_hd__nand2_2 _31214_ (.A(_09177_),
    .B(_08865_),
    .Y(_09185_));
 sky130_fd_sc_hd__o211a_2 _31215_ (.A1(_09184_),
    .A2(_09185_),
    .B1(_09182_),
    .C1(_09179_),
    .X(_09186_));
 sky130_fd_sc_hd__nor2_2 _31216_ (.A(_09183_),
    .B(_09186_),
    .Y(_09187_));
 sky130_fd_sc_hd__a21oi_2 _31217_ (.A1(_08874_),
    .A2(_08880_),
    .B1(_08883_),
    .Y(_09188_));
 sky130_fd_sc_hd__a31oi_2 _31218_ (.A1(_08564_),
    .A2(_08565_),
    .A3(_08566_),
    .B1(_08279_),
    .Y(_09189_));
 sky130_fd_sc_hd__o21ai_2 _31219_ (.A1(_08592_),
    .A2(_09189_),
    .B1(_08886_),
    .Y(_09190_));
 sky130_fd_sc_hd__o2111a_2 _31220_ (.A1(_09188_),
    .A2(_09190_),
    .B1(_08895_),
    .C1(_08579_),
    .D1(_08571_),
    .X(_09191_));
 sky130_fd_sc_hd__a21oi_2 _31221_ (.A1(_08885_),
    .A2(_08886_),
    .B1(_08593_),
    .Y(_09192_));
 sky130_fd_sc_hd__a21oi_2 _31222_ (.A1(_08887_),
    .A2(_08579_),
    .B1(_09192_),
    .Y(_09193_));
 sky130_fd_sc_hd__a21o_2 _31223_ (.A1(_08589_),
    .A2(_09191_),
    .B1(_09193_),
    .X(_09194_));
 sky130_fd_sc_hd__xor2_2 _31224_ (.A(_09187_),
    .B(_09194_),
    .X(_02645_));
 sky130_fd_sc_hd__a31o_2 _31225_ (.A1(_09006_),
    .A2(_09155_),
    .A3(_09002_),
    .B1(_09149_),
    .X(_09195_));
 sky130_fd_sc_hd__inv_2 _31226_ (.A(_08919_),
    .Y(_09196_));
 sky130_fd_sc_hd__o21a_2 _31227_ (.A1(_08929_),
    .A2(_08928_),
    .B1(_08914_),
    .X(_09197_));
 sky130_fd_sc_hd__nand2_2 _31228_ (.A(_05402_),
    .B(_08103_),
    .Y(_09198_));
 sky130_fd_sc_hd__buf_1 _31229_ (.A(_08085_),
    .X(_09199_));
 sky130_fd_sc_hd__nand2_2 _31230_ (.A(_05721_),
    .B(_09199_),
    .Y(_09200_));
 sky130_fd_sc_hd__nor2_2 _31231_ (.A(_09198_),
    .B(_09200_),
    .Y(_09201_));
 sky130_fd_sc_hd__and2_2 _31232_ (.A(_09198_),
    .B(_09200_),
    .X(_09202_));
 sky130_fd_sc_hd__buf_1 _31233_ (.A(\pcpi_mul.rs1[27] ),
    .X(_09203_));
 sky130_fd_sc_hd__nand2_2 _31234_ (.A(_06057_),
    .B(_09203_),
    .Y(_09204_));
 sky130_fd_sc_hd__inv_2 _31235_ (.A(_09204_),
    .Y(_09205_));
 sky130_fd_sc_hd__o21ai_2 _31236_ (.A1(_09201_),
    .A2(_09202_),
    .B1(_09205_),
    .Y(_09206_));
 sky130_fd_sc_hd__or2_2 _31237_ (.A(_09198_),
    .B(_09200_),
    .X(_09207_));
 sky130_fd_sc_hd__nand2_2 _31238_ (.A(_09198_),
    .B(_09200_),
    .Y(_09208_));
 sky130_fd_sc_hd__nand3_2 _31239_ (.A(_09207_),
    .B(_09204_),
    .C(_09208_),
    .Y(_09209_));
 sky130_fd_sc_hd__a21oi_2 _31240_ (.A1(_08907_),
    .A2(_08908_),
    .B1(_08904_),
    .Y(_09210_));
 sky130_fd_sc_hd__nand3_2 _31241_ (.A(_09206_),
    .B(_09209_),
    .C(_09210_),
    .Y(_09211_));
 sky130_fd_sc_hd__o21ai_2 _31242_ (.A1(_09201_),
    .A2(_09202_),
    .B1(_09204_),
    .Y(_09212_));
 sky130_fd_sc_hd__nand3_2 _31243_ (.A(_09207_),
    .B(_09205_),
    .C(_09208_),
    .Y(_09213_));
 sky130_fd_sc_hd__nand2_2 _31244_ (.A(_08915_),
    .B(_08909_),
    .Y(_09214_));
 sky130_fd_sc_hd__nand3_2 _31245_ (.A(_09212_),
    .B(_09213_),
    .C(_09214_),
    .Y(_09215_));
 sky130_fd_sc_hd__buf_1 _31246_ (.A(_08905_),
    .X(_09216_));
 sky130_fd_sc_hd__nand2_2 _31247_ (.A(_06219_),
    .B(_19565_),
    .Y(_09217_));
 sky130_fd_sc_hd__a21o_2 _31248_ (.A1(_05144_),
    .A2(_09216_),
    .B1(_09217_),
    .X(_09218_));
 sky130_fd_sc_hd__buf_1 _31249_ (.A(_08920_),
    .X(_09219_));
 sky130_fd_sc_hd__buf_1 _31250_ (.A(_19561_),
    .X(_09220_));
 sky130_fd_sc_hd__nand2_2 _31251_ (.A(_19401_),
    .B(_09220_),
    .Y(_09221_));
 sky130_fd_sc_hd__a21o_2 _31252_ (.A1(_05141_),
    .A2(_09219_),
    .B1(_09221_),
    .X(_09222_));
 sky130_fd_sc_hd__buf_1 _31253_ (.A(_08662_),
    .X(_09223_));
 sky130_fd_sc_hd__nand2_2 _31254_ (.A(_05116_),
    .B(_09223_),
    .Y(_09224_));
 sky130_fd_sc_hd__a21oi_2 _31255_ (.A1(_09218_),
    .A2(_09222_),
    .B1(_09224_),
    .Y(_09225_));
 sky130_fd_sc_hd__buf_1 _31256_ (.A(_08487_),
    .X(_09226_));
 sky130_fd_sc_hd__o211a_2 _31257_ (.A1(_05151_),
    .A2(_09226_),
    .B1(_09222_),
    .C1(_09218_),
    .X(_09227_));
 sky130_fd_sc_hd__nor2_2 _31258_ (.A(_09225_),
    .B(_09227_),
    .Y(_09228_));
 sky130_fd_sc_hd__a21oi_2 _31259_ (.A1(_09211_),
    .A2(_09215_),
    .B1(_09228_),
    .Y(_09229_));
 sky130_fd_sc_hd__o21a_2 _31260_ (.A1(_09201_),
    .A2(_09202_),
    .B1(_09204_),
    .X(_09230_));
 sky130_fd_sc_hd__nand2_2 _31261_ (.A(_09213_),
    .B(_09214_),
    .Y(_09231_));
 sky130_fd_sc_hd__o211a_2 _31262_ (.A1(_09230_),
    .A2(_09231_),
    .B1(_09211_),
    .C1(_09228_),
    .X(_09232_));
 sky130_fd_sc_hd__o22ai_2 _31263_ (.A1(_09196_),
    .A2(_09197_),
    .B1(_09229_),
    .B2(_09232_),
    .Y(_09233_));
 sky130_fd_sc_hd__nand2_2 _31264_ (.A(_08931_),
    .B(_08919_),
    .Y(_09234_));
 sky130_fd_sc_hd__nand2_2 _31265_ (.A(_09234_),
    .B(_08914_),
    .Y(_09235_));
 sky130_fd_sc_hd__nand3_2 _31266_ (.A(_09228_),
    .B(_09215_),
    .C(_09211_),
    .Y(_09236_));
 sky130_fd_sc_hd__a21o_2 _31267_ (.A1(_09211_),
    .A2(_09215_),
    .B1(_09228_),
    .X(_09237_));
 sky130_fd_sc_hd__nand3_2 _31268_ (.A(_09235_),
    .B(_09236_),
    .C(_09237_),
    .Y(_09238_));
 sky130_fd_sc_hd__nor2_2 _31269_ (.A(_08923_),
    .B(_08925_),
    .Y(_09239_));
 sky130_fd_sc_hd__or2_2 _31270_ (.A(_09239_),
    .B(_08929_),
    .X(_09240_));
 sky130_fd_sc_hd__a21oi_2 _31271_ (.A1(_09233_),
    .A2(_09238_),
    .B1(_09240_),
    .Y(_09241_));
 sky130_fd_sc_hd__o211a_2 _31272_ (.A1(_09239_),
    .A2(_08929_),
    .B1(_09238_),
    .C1(_09233_),
    .X(_09242_));
 sky130_fd_sc_hd__nor2_2 _31273_ (.A(_09241_),
    .B(_09242_),
    .Y(_09243_));
 sky130_fd_sc_hd__and2_2 _31274_ (.A(_08966_),
    .B(_08969_),
    .X(_09244_));
 sky130_fd_sc_hd__inv_2 _31275_ (.A(\pcpi_mul.rs1[20] ),
    .Y(_09245_));
 sky130_fd_sc_hd__buf_1 _31276_ (.A(_09245_),
    .X(_09246_));
 sky130_fd_sc_hd__buf_1 _31277_ (.A(_06334_),
    .X(_09247_));
 sky130_fd_sc_hd__buf_1 _31278_ (.A(\pcpi_mul.rs1[19] ),
    .X(_09248_));
 sky130_fd_sc_hd__nand3_2 _31279_ (.A(_19380_),
    .B(_09247_),
    .C(_09248_),
    .Y(_09249_));
 sky130_fd_sc_hd__buf_1 _31280_ (.A(_07605_),
    .X(_09250_));
 sky130_fd_sc_hd__nand2_2 _31281_ (.A(_05764_),
    .B(_09250_),
    .Y(_09251_));
 sky130_fd_sc_hd__a22o_2 _31282_ (.A1(_07797_),
    .A2(_19582_),
    .B1(_08949_),
    .B2(_19580_),
    .X(_09252_));
 sky130_fd_sc_hd__o211ai_2 _31283_ (.A1(_09246_),
    .A2(_09249_),
    .B1(_09251_),
    .C1(_09252_),
    .Y(_09253_));
 sky130_fd_sc_hd__buf_1 _31284_ (.A(_05760_),
    .X(_09254_));
 sky130_fd_sc_hd__a22oi_2 _31285_ (.A1(_08948_),
    .A2(_08490_),
    .B1(_09254_),
    .B2(_08108_),
    .Y(_09255_));
 sky130_fd_sc_hd__buf_1 _31286_ (.A(_09245_),
    .X(_09256_));
 sky130_fd_sc_hd__nor2_2 _31287_ (.A(_09256_),
    .B(_09249_),
    .Y(_09257_));
 sky130_fd_sc_hd__inv_2 _31288_ (.A(_09251_),
    .Y(_09258_));
 sky130_fd_sc_hd__o21ai_2 _31289_ (.A1(_09255_),
    .A2(_09257_),
    .B1(_09258_),
    .Y(_09259_));
 sky130_fd_sc_hd__o2111ai_2 _31290_ (.A1(_09053_),
    .A2(_09050_),
    .B1(_09057_),
    .C1(_09253_),
    .D1(_09259_),
    .Y(_09260_));
 sky130_fd_sc_hd__o21ai_2 _31291_ (.A1(_09255_),
    .A2(_09257_),
    .B1(_09251_),
    .Y(_09261_));
 sky130_fd_sc_hd__o21ai_2 _31292_ (.A1(_09053_),
    .A2(_09050_),
    .B1(_09057_),
    .Y(_09262_));
 sky130_fd_sc_hd__buf_1 _31293_ (.A(_09256_),
    .X(_09263_));
 sky130_fd_sc_hd__o211ai_2 _31294_ (.A1(_09263_),
    .A2(_09249_),
    .B1(_09258_),
    .C1(_09252_),
    .Y(_09264_));
 sky130_fd_sc_hd__nand3_2 _31295_ (.A(_09261_),
    .B(_09262_),
    .C(_09264_),
    .Y(_09265_));
 sky130_fd_sc_hd__a21o_2 _31296_ (.A1(_08960_),
    .A2(_08958_),
    .B1(_08952_),
    .X(_09266_));
 sky130_fd_sc_hd__a21o_2 _31297_ (.A1(_09260_),
    .A2(_09265_),
    .B1(_09266_),
    .X(_09267_));
 sky130_fd_sc_hd__nand3_2 _31298_ (.A(_09260_),
    .B(_09266_),
    .C(_09265_),
    .Y(_09268_));
 sky130_fd_sc_hd__a21oi_2 _31299_ (.A1(_09043_),
    .A2(_09044_),
    .B1(_09040_),
    .Y(_09269_));
 sky130_fd_sc_hd__a32o_2 _31300_ (.A1(_09043_),
    .A2(_09040_),
    .A3(_09044_),
    .B1(_08742_),
    .B2(_08749_),
    .X(_09270_));
 sky130_fd_sc_hd__o2bb2ai_2 _31301_ (.A1_N(_09062_),
    .A2_N(_09049_),
    .B1(_09269_),
    .B2(_09270_),
    .Y(_09271_));
 sky130_fd_sc_hd__a21oi_2 _31302_ (.A1(_09267_),
    .A2(_09268_),
    .B1(_09271_),
    .Y(_09272_));
 sky130_fd_sc_hd__inv_2 _31303_ (.A(_09265_),
    .Y(_09273_));
 sky130_fd_sc_hd__nand2_2 _31304_ (.A(_09260_),
    .B(_09266_),
    .Y(_09274_));
 sky130_fd_sc_hd__o211a_2 _31305_ (.A1(_09273_),
    .A2(_09274_),
    .B1(_09271_),
    .C1(_09267_),
    .X(_09275_));
 sky130_fd_sc_hd__o22ai_2 _31306_ (.A1(_08975_),
    .A2(_09244_),
    .B1(_09272_),
    .B2(_09275_),
    .Y(_09276_));
 sky130_fd_sc_hd__a21oi_2 _31307_ (.A1(_08980_),
    .A2(_08977_),
    .B1(_08976_),
    .Y(_09277_));
 sky130_fd_sc_hd__a21o_2 _31308_ (.A1(_09267_),
    .A2(_09268_),
    .B1(_09271_),
    .X(_09278_));
 sky130_fd_sc_hd__nand2_2 _31309_ (.A(_08974_),
    .B(_08962_),
    .Y(_09279_));
 sky130_fd_sc_hd__inv_2 _31310_ (.A(_09279_),
    .Y(_09280_));
 sky130_fd_sc_hd__nand3_2 _31311_ (.A(_09267_),
    .B(_09271_),
    .C(_09268_),
    .Y(_09281_));
 sky130_fd_sc_hd__nand3_2 _31312_ (.A(_09278_),
    .B(_09280_),
    .C(_09281_),
    .Y(_09282_));
 sky130_fd_sc_hd__nand3_2 _31313_ (.A(_09276_),
    .B(_09277_),
    .C(_09282_),
    .Y(_09283_));
 sky130_fd_sc_hd__o21ai_2 _31314_ (.A1(_09272_),
    .A2(_09275_),
    .B1(_09280_),
    .Y(_09284_));
 sky130_fd_sc_hd__o21ai_2 _31315_ (.A1(_08978_),
    .A2(_08973_),
    .B1(_08981_),
    .Y(_09285_));
 sky130_fd_sc_hd__nand3_2 _31316_ (.A(_09278_),
    .B(_09279_),
    .C(_09281_),
    .Y(_09286_));
 sky130_fd_sc_hd__nand3_2 _31317_ (.A(_09284_),
    .B(_09285_),
    .C(_09286_),
    .Y(_09287_));
 sky130_fd_sc_hd__nand3_2 _31318_ (.A(_09243_),
    .B(_09283_),
    .C(_09287_),
    .Y(_09288_));
 sky130_fd_sc_hd__o2bb2ai_2 _31319_ (.A1_N(_09283_),
    .A2_N(_09287_),
    .B1(_09242_),
    .B2(_09241_),
    .Y(_09289_));
 sky130_fd_sc_hd__a21oi_2 _31320_ (.A1(_08770_),
    .A2(_08768_),
    .B1(_08731_),
    .Y(_09290_));
 sky130_fd_sc_hd__nand2_2 _31321_ (.A(_09078_),
    .B(_09290_),
    .Y(_09291_));
 sky130_fd_sc_hd__inv_2 _31322_ (.A(_09291_),
    .Y(_09292_));
 sky130_fd_sc_hd__and3_2 _31323_ (.A(_09066_),
    .B(_09074_),
    .C(_08826_),
    .X(_09293_));
 sky130_fd_sc_hd__o2bb2ai_2 _31324_ (.A1_N(_09288_),
    .A2_N(_09289_),
    .B1(_09292_),
    .B2(_09293_),
    .Y(_09294_));
 sky130_fd_sc_hd__and3_2 _31325_ (.A(_09076_),
    .B(_09077_),
    .C(_08830_),
    .X(_09295_));
 sky130_fd_sc_hd__a31oi_2 _31326_ (.A1(_09066_),
    .A2(_09074_),
    .A3(_08826_),
    .B1(_09290_),
    .Y(_09296_));
 sky130_fd_sc_hd__o211ai_2 _31327_ (.A1(_09295_),
    .A2(_09296_),
    .B1(_09288_),
    .C1(_09289_),
    .Y(_09297_));
 sky130_fd_sc_hd__nand2_2 _31328_ (.A(_08944_),
    .B(_08989_),
    .Y(_09298_));
 sky130_fd_sc_hd__nand2_2 _31329_ (.A(_09298_),
    .B(_08984_),
    .Y(_09299_));
 sky130_fd_sc_hd__a21oi_2 _31330_ (.A1(_09294_),
    .A2(_09297_),
    .B1(_09299_),
    .Y(_09300_));
 sky130_fd_sc_hd__inv_2 _31331_ (.A(_09299_),
    .Y(_09301_));
 sky130_fd_sc_hd__a22oi_2 _31332_ (.A1(_09075_),
    .A2(_09291_),
    .B1(_09289_),
    .B2(_09288_),
    .Y(_09302_));
 sky130_fd_sc_hd__o211a_2 _31333_ (.A1(_09295_),
    .A2(_09296_),
    .B1(_09288_),
    .C1(_09289_),
    .X(_09303_));
 sky130_fd_sc_hd__nor3_2 _31334_ (.A(_09301_),
    .B(_09302_),
    .C(_09303_),
    .Y(_09304_));
 sky130_fd_sc_hd__inv_2 _31335_ (.A(_09112_),
    .Y(_09305_));
 sky130_fd_sc_hd__nand2_2 _31336_ (.A(_09119_),
    .B(_09133_),
    .Y(_09306_));
 sky130_fd_sc_hd__a22oi_2 _31337_ (.A1(_08385_),
    .A2(_06629_),
    .B1(_08383_),
    .B2(_06502_),
    .Y(_09307_));
 sky130_fd_sc_hd__nand3_2 _31338_ (.A(_19336_),
    .B(\pcpi_mul.rs2[22] ),
    .C(_05206_),
    .Y(_09308_));
 sky130_fd_sc_hd__nor2_2 _31339_ (.A(_05856_),
    .B(_09308_),
    .Y(_09309_));
 sky130_fd_sc_hd__nand2_2 _31340_ (.A(\pcpi_mul.rs2[21] ),
    .B(_06609_),
    .Y(_09310_));
 sky130_fd_sc_hd__inv_2 _31341_ (.A(_09310_),
    .Y(_09311_));
 sky130_fd_sc_hd__o21ai_2 _31342_ (.A1(_09307_),
    .A2(_09309_),
    .B1(_09311_),
    .Y(_09312_));
 sky130_fd_sc_hd__a21oi_2 _31343_ (.A1(_09085_),
    .A2(_09087_),
    .B1(_09084_),
    .Y(_09313_));
 sky130_fd_sc_hd__a22o_2 _31344_ (.A1(_08385_),
    .A2(_05338_),
    .B1(_07974_),
    .B2(_05765_),
    .X(_09314_));
 sky130_fd_sc_hd__o211ai_2 _31345_ (.A1(_05865_),
    .A2(_09308_),
    .B1(_09310_),
    .C1(_09314_),
    .Y(_09315_));
 sky130_fd_sc_hd__nand3_2 _31346_ (.A(_09312_),
    .B(_09313_),
    .C(_09315_),
    .Y(_09316_));
 sky130_fd_sc_hd__o21ai_2 _31347_ (.A1(_09307_),
    .A2(_09309_),
    .B1(_09310_),
    .Y(_09317_));
 sky130_fd_sc_hd__o21ai_2 _31348_ (.A1(_09086_),
    .A2(_09090_),
    .B1(_09096_),
    .Y(_09318_));
 sky130_fd_sc_hd__o211ai_2 _31349_ (.A1(_05865_),
    .A2(_09308_),
    .B1(_09311_),
    .C1(_09314_),
    .Y(_09319_));
 sky130_fd_sc_hd__nand3_2 _31350_ (.A(_09317_),
    .B(_09318_),
    .C(_09319_),
    .Y(_09320_));
 sky130_fd_sc_hd__a22oi_2 _31351_ (.A1(_09101_),
    .A2(_06617_),
    .B1(_19350_),
    .B2(_06052_),
    .Y(_09321_));
 sky130_fd_sc_hd__nand3_2 _31352_ (.A(_07903_),
    .B(_07723_),
    .C(_05426_),
    .Y(_09322_));
 sky130_fd_sc_hd__nor2_2 _31353_ (.A(_05731_),
    .B(_09322_),
    .Y(_09323_));
 sky130_fd_sc_hd__nand2_2 _31354_ (.A(_07475_),
    .B(_06327_),
    .Y(_09324_));
 sky130_fd_sc_hd__inv_2 _31355_ (.A(_09324_),
    .Y(_09325_));
 sky130_fd_sc_hd__o21ai_2 _31356_ (.A1(_09321_),
    .A2(_09323_),
    .B1(_09325_),
    .Y(_09326_));
 sky130_fd_sc_hd__a22o_2 _31357_ (.A1(_19347_),
    .A2(_06617_),
    .B1(_19350_),
    .B2(_06052_),
    .X(_09327_));
 sky130_fd_sc_hd__o211ai_2 _31358_ (.A1(_05732_),
    .A2(_09322_),
    .B1(_09324_),
    .C1(_09327_),
    .Y(_09328_));
 sky130_fd_sc_hd__nand2_2 _31359_ (.A(_09326_),
    .B(_09328_),
    .Y(_09329_));
 sky130_fd_sc_hd__a21oi_2 _31360_ (.A1(_09316_),
    .A2(_09320_),
    .B1(_09329_),
    .Y(_09330_));
 sky130_fd_sc_hd__and3_2 _31361_ (.A(_09316_),
    .B(_09320_),
    .C(_09329_),
    .X(_09331_));
 sky130_fd_sc_hd__nand2_2 _31362_ (.A(_09130_),
    .B(_08787_),
    .Y(_09332_));
 sky130_fd_sc_hd__o21ai_2 _31363_ (.A1(_09330_),
    .A2(_09331_),
    .B1(_09332_),
    .Y(_09333_));
 sky130_fd_sc_hd__a21o_2 _31364_ (.A1(_09316_),
    .A2(_09320_),
    .B1(_09329_),
    .X(_09334_));
 sky130_fd_sc_hd__nand3_2 _31365_ (.A(_09316_),
    .B(_09320_),
    .C(_09329_),
    .Y(_09335_));
 sky130_fd_sc_hd__nand3_2 _31366_ (.A(_09334_),
    .B(_09129_),
    .C(_09335_),
    .Y(_09336_));
 sky130_fd_sc_hd__nand2_2 _31367_ (.A(_09111_),
    .B(_09092_),
    .Y(_09337_));
 sky130_fd_sc_hd__a21oi_2 _31368_ (.A1(_09333_),
    .A2(_09336_),
    .B1(_09337_),
    .Y(_09338_));
 sky130_fd_sc_hd__buf_1 _31369_ (.A(\pcpi_mul.rs2[26] ),
    .X(_09339_));
 sky130_fd_sc_hd__nand2_2 _31370_ (.A(_09339_),
    .B(_05105_),
    .Y(_09340_));
 sky130_fd_sc_hd__nand2_2 _31371_ (.A(_19330_),
    .B(_05323_),
    .Y(_09341_));
 sky130_fd_sc_hd__nor2_2 _31372_ (.A(_09340_),
    .B(_09341_),
    .Y(_09342_));
 sky130_fd_sc_hd__nand2_2 _31373_ (.A(\pcpi_mul.rs2[24] ),
    .B(_05271_),
    .Y(_09343_));
 sky130_fd_sc_hd__inv_2 _31374_ (.A(_09343_),
    .Y(_09344_));
 sky130_fd_sc_hd__nand2_2 _31375_ (.A(_09340_),
    .B(_09341_),
    .Y(_09345_));
 sky130_fd_sc_hd__nand2_2 _31376_ (.A(_09344_),
    .B(_09345_),
    .Y(_09346_));
 sky130_fd_sc_hd__a31o_2 _31377_ (.A1(_09127_),
    .A2(_19334_),
    .A3(_19634_),
    .B1(_09123_),
    .X(_09347_));
 sky130_fd_sc_hd__and2_2 _31378_ (.A(_09340_),
    .B(_09341_),
    .X(_09348_));
 sky130_fd_sc_hd__o21ai_2 _31379_ (.A1(_09342_),
    .A2(_09348_),
    .B1(_09343_),
    .Y(_09349_));
 sky130_fd_sc_hd__o211ai_2 _31380_ (.A1(_09342_),
    .A2(_09346_),
    .B1(_09347_),
    .C1(_09349_),
    .Y(_09350_));
 sky130_fd_sc_hd__o21ai_2 _31381_ (.A1(_09342_),
    .A2(_09348_),
    .B1(_09344_),
    .Y(_09351_));
 sky130_fd_sc_hd__nand3b_2 _31382_ (.A_N(_09342_),
    .B(_09345_),
    .C(_09343_),
    .Y(_09352_));
 sky130_fd_sc_hd__a21oi_2 _31383_ (.A1(_09125_),
    .A2(_09127_),
    .B1(_09123_),
    .Y(_09353_));
 sky130_fd_sc_hd__nand3_2 _31384_ (.A(_09351_),
    .B(_09352_),
    .C(_09353_),
    .Y(_09354_));
 sky130_fd_sc_hd__nand2_2 _31385_ (.A(_09350_),
    .B(_09354_),
    .Y(_09355_));
 sky130_fd_sc_hd__inv_2 _31386_ (.A(\pcpi_mul.rs2[27] ),
    .Y(_09356_));
 sky130_fd_sc_hd__buf_1 _31387_ (.A(_09356_),
    .X(_09357_));
 sky130_fd_sc_hd__buf_1 _31388_ (.A(_09357_),
    .X(_09358_));
 sky130_fd_sc_hd__nor2_2 _31389_ (.A(_09358_),
    .B(_04839_),
    .Y(_09359_));
 sky130_fd_sc_hd__and2_2 _31390_ (.A(_09355_),
    .B(_09359_),
    .X(_09360_));
 sky130_fd_sc_hd__nor2_2 _31391_ (.A(_09359_),
    .B(_09355_),
    .Y(_09361_));
 sky130_fd_sc_hd__a21oi_2 _31392_ (.A1(_09334_),
    .A2(_09335_),
    .B1(_09129_),
    .Y(_09362_));
 sky130_fd_sc_hd__nand2_2 _31393_ (.A(_09336_),
    .B(_09337_),
    .Y(_09363_));
 sky130_fd_sc_hd__o22ai_2 _31394_ (.A1(_09360_),
    .A2(_09361_),
    .B1(_09362_),
    .B2(_09363_),
    .Y(_09364_));
 sky130_fd_sc_hd__nor2_2 _31395_ (.A(_09338_),
    .B(_09364_),
    .Y(_09365_));
 sky130_fd_sc_hd__nand3_2 _31396_ (.A(_09350_),
    .B(_09354_),
    .C(_09359_),
    .Y(_09366_));
 sky130_fd_sc_hd__inv_2 _31397_ (.A(_09359_),
    .Y(_09367_));
 sky130_fd_sc_hd__nand2_2 _31398_ (.A(_09355_),
    .B(_09367_),
    .Y(_09368_));
 sky130_fd_sc_hd__nor3_2 _31399_ (.A(_09330_),
    .B(_09332_),
    .C(_09331_),
    .Y(_09369_));
 sky130_fd_sc_hd__a21boi_2 _31400_ (.A1(_09107_),
    .A2(_09098_),
    .B1_N(_09092_),
    .Y(_09370_));
 sky130_fd_sc_hd__o21ai_2 _31401_ (.A1(_09362_),
    .A2(_09369_),
    .B1(_09370_),
    .Y(_09371_));
 sky130_fd_sc_hd__nand3_2 _31402_ (.A(_09333_),
    .B(_09336_),
    .C(_09337_),
    .Y(_09372_));
 sky130_fd_sc_hd__a22oi_2 _31403_ (.A1(_09366_),
    .A2(_09368_),
    .B1(_09371_),
    .B2(_09372_),
    .Y(_09373_));
 sky130_fd_sc_hd__o22ai_2 _31404_ (.A1(_09305_),
    .A2(_09306_),
    .B1(_09365_),
    .B2(_09373_),
    .Y(_09374_));
 sky130_fd_sc_hd__nor2_2 _31405_ (.A(_09362_),
    .B(_09363_),
    .Y(_09375_));
 sky130_fd_sc_hd__nand2_2 _31406_ (.A(_09368_),
    .B(_09366_),
    .Y(_09376_));
 sky130_fd_sc_hd__o21ai_2 _31407_ (.A1(_09338_),
    .A2(_09375_),
    .B1(_09376_),
    .Y(_09377_));
 sky130_fd_sc_hd__nand3b_2 _31408_ (.A_N(_09376_),
    .B(_09371_),
    .C(_09372_),
    .Y(_09378_));
 sky130_fd_sc_hd__nand3_2 _31409_ (.A(_09377_),
    .B(_09378_),
    .C(_09139_),
    .Y(_09379_));
 sky130_fd_sc_hd__nand2_2 _31410_ (.A(_09374_),
    .B(_09379_),
    .Y(_09380_));
 sky130_fd_sc_hd__a22oi_2 _31411_ (.A1(_07481_),
    .A2(_19623_),
    .B1(_07907_),
    .B2(_19620_),
    .Y(_09381_));
 sky130_fd_sc_hd__o21a_2 _31412_ (.A1(_09381_),
    .A2(_09103_),
    .B1(_09100_),
    .X(_09382_));
 sky130_fd_sc_hd__a22oi_2 _31413_ (.A1(_19355_),
    .A2(_09010_),
    .B1(_19358_),
    .B2(_06074_),
    .Y(_09383_));
 sky130_fd_sc_hd__nand3_2 _31414_ (.A(_06822_),
    .B(_06824_),
    .C(_19609_),
    .Y(_09384_));
 sky130_fd_sc_hd__nor2_2 _31415_ (.A(_06688_),
    .B(_09384_),
    .Y(_09385_));
 sky130_fd_sc_hd__buf_1 _31416_ (.A(_07890_),
    .X(_09386_));
 sky130_fd_sc_hd__nand2_2 _31417_ (.A(_09386_),
    .B(_06538_),
    .Y(_09387_));
 sky130_fd_sc_hd__inv_2 _31418_ (.A(_09387_),
    .Y(_09388_));
 sky130_fd_sc_hd__o21ai_2 _31419_ (.A1(_09383_),
    .A2(_09385_),
    .B1(_09388_),
    .Y(_09389_));
 sky130_fd_sc_hd__a22o_2 _31420_ (.A1(_19355_),
    .A2(_09010_),
    .B1(_09009_),
    .B2(_05911_),
    .X(_09390_));
 sky130_fd_sc_hd__o211ai_2 _31421_ (.A1(_06225_),
    .A2(_09384_),
    .B1(_09387_),
    .C1(_09390_),
    .Y(_09391_));
 sky130_fd_sc_hd__nand3_2 _31422_ (.A(_09382_),
    .B(_09389_),
    .C(_09391_),
    .Y(_09392_));
 sky130_fd_sc_hd__o21ai_2 _31423_ (.A1(_09383_),
    .A2(_09385_),
    .B1(_09387_),
    .Y(_09393_));
 sky130_fd_sc_hd__o211ai_2 _31424_ (.A1(_06225_),
    .A2(_09384_),
    .B1(_09388_),
    .C1(_09390_),
    .Y(_09394_));
 sky130_fd_sc_hd__o21ai_2 _31425_ (.A1(_09103_),
    .A2(_09381_),
    .B1(_09100_),
    .Y(_09395_));
 sky130_fd_sc_hd__nand3_2 _31426_ (.A(_09393_),
    .B(_09394_),
    .C(_09395_),
    .Y(_09396_));
 sky130_fd_sc_hd__nand2_2 _31427_ (.A(_09392_),
    .B(_09396_),
    .Y(_09397_));
 sky130_fd_sc_hd__a21oi_2 _31428_ (.A1(_09020_),
    .A2(_09017_),
    .B1(_09014_),
    .Y(_09398_));
 sky130_fd_sc_hd__nand2_2 _31429_ (.A(_09397_),
    .B(_09398_),
    .Y(_09399_));
 sky130_fd_sc_hd__inv_2 _31430_ (.A(_09398_),
    .Y(_09400_));
 sky130_fd_sc_hd__nand3_2 _31431_ (.A(_09392_),
    .B(_09396_),
    .C(_09400_),
    .Y(_09401_));
 sky130_fd_sc_hd__nand2_2 _31432_ (.A(_09028_),
    .B(_09031_),
    .Y(_09402_));
 sky130_fd_sc_hd__nand2_2 _31433_ (.A(_09402_),
    .B(_09023_),
    .Y(_09403_));
 sky130_fd_sc_hd__a21oi_2 _31434_ (.A1(_09399_),
    .A2(_09401_),
    .B1(_09403_),
    .Y(_09404_));
 sky130_fd_sc_hd__inv_2 _31435_ (.A(_09396_),
    .Y(_09405_));
 sky130_fd_sc_hd__nand2_2 _31436_ (.A(_09392_),
    .B(_09400_),
    .Y(_09406_));
 sky130_fd_sc_hd__o211a_2 _31437_ (.A1(_09405_),
    .A2(_09406_),
    .B1(_09403_),
    .C1(_09399_),
    .X(_09407_));
 sky130_fd_sc_hd__o21ai_2 _31438_ (.A1(_09039_),
    .A2(_09037_),
    .B1(_09043_),
    .Y(_09408_));
 sky130_fd_sc_hd__nand2_2 _31439_ (.A(_07012_),
    .B(_07311_),
    .Y(_09409_));
 sky130_fd_sc_hd__nand2_2 _31440_ (.A(_19365_),
    .B(_08761_),
    .Y(_09410_));
 sky130_fd_sc_hd__nor2_2 _31441_ (.A(_09409_),
    .B(_09410_),
    .Y(_09411_));
 sky130_fd_sc_hd__and2_2 _31442_ (.A(_09409_),
    .B(_09410_),
    .X(_09412_));
 sky130_fd_sc_hd__nand2_2 _31443_ (.A(_06628_),
    .B(_19594_),
    .Y(_09413_));
 sky130_fd_sc_hd__inv_2 _31444_ (.A(_09413_),
    .Y(_09414_));
 sky130_fd_sc_hd__o21ai_2 _31445_ (.A1(_09411_),
    .A2(_09412_),
    .B1(_09414_),
    .Y(_09415_));
 sky130_fd_sc_hd__or2_2 _31446_ (.A(_09409_),
    .B(_09410_),
    .X(_09416_));
 sky130_fd_sc_hd__nand2_2 _31447_ (.A(_09409_),
    .B(_09410_),
    .Y(_09417_));
 sky130_fd_sc_hd__nand3_2 _31448_ (.A(_09416_),
    .B(_09417_),
    .C(_09413_),
    .Y(_09418_));
 sky130_fd_sc_hd__nand3b_2 _31449_ (.A_N(_09408_),
    .B(_09415_),
    .C(_09418_),
    .Y(_09419_));
 sky130_fd_sc_hd__nand2_2 _31450_ (.A(_09414_),
    .B(_09417_),
    .Y(_09420_));
 sky130_fd_sc_hd__o21ai_2 _31451_ (.A1(_09411_),
    .A2(_09412_),
    .B1(_09413_),
    .Y(_09421_));
 sky130_fd_sc_hd__o211ai_2 _31452_ (.A1(_09411_),
    .A2(_09420_),
    .B1(_09408_),
    .C1(_09421_),
    .Y(_09422_));
 sky130_fd_sc_hd__nand2_2 _31453_ (.A(_09419_),
    .B(_09422_),
    .Y(_09423_));
 sky130_fd_sc_hd__nand2_2 _31454_ (.A(_06500_),
    .B(_19590_),
    .Y(_09424_));
 sky130_fd_sc_hd__nand2_2 _31455_ (.A(_05670_),
    .B(_06728_),
    .Y(_09425_));
 sky130_fd_sc_hd__or2_2 _31456_ (.A(_09424_),
    .B(_09425_),
    .X(_09426_));
 sky130_fd_sc_hd__nand2_2 _31457_ (.A(_06616_),
    .B(_08596_),
    .Y(_09427_));
 sky130_fd_sc_hd__nand2_2 _31458_ (.A(_09424_),
    .B(_09425_),
    .Y(_09428_));
 sky130_fd_sc_hd__nand3_2 _31459_ (.A(_09426_),
    .B(_09427_),
    .C(_09428_),
    .Y(_09429_));
 sky130_fd_sc_hd__a22oi_2 _31460_ (.A1(_19371_),
    .A2(_06750_),
    .B1(_19374_),
    .B2(_07380_),
    .Y(_09430_));
 sky130_fd_sc_hd__nor2_2 _31461_ (.A(_09424_),
    .B(_09425_),
    .Y(_09431_));
 sky130_fd_sc_hd__inv_2 _31462_ (.A(_09427_),
    .Y(_09432_));
 sky130_fd_sc_hd__o21ai_2 _31463_ (.A1(_09430_),
    .A2(_09431_),
    .B1(_09432_),
    .Y(_09433_));
 sky130_fd_sc_hd__nand2_2 _31464_ (.A(_09429_),
    .B(_09433_),
    .Y(_09434_));
 sky130_fd_sc_hd__nand2_2 _31465_ (.A(_09423_),
    .B(_09434_),
    .Y(_09435_));
 sky130_fd_sc_hd__inv_2 _31466_ (.A(_09434_),
    .Y(_09436_));
 sky130_fd_sc_hd__nand3_2 _31467_ (.A(_09436_),
    .B(_09419_),
    .C(_09422_),
    .Y(_09437_));
 sky130_fd_sc_hd__nand2_2 _31468_ (.A(_09435_),
    .B(_09437_),
    .Y(_09438_));
 sky130_fd_sc_hd__o21ai_2 _31469_ (.A1(_09404_),
    .A2(_09407_),
    .B1(_09438_),
    .Y(_09439_));
 sky130_fd_sc_hd__a21o_2 _31470_ (.A1(_09399_),
    .A2(_09401_),
    .B1(_09403_),
    .X(_09440_));
 sky130_fd_sc_hd__nand3_2 _31471_ (.A(_09399_),
    .B(_09403_),
    .C(_09401_),
    .Y(_09441_));
 sky130_fd_sc_hd__nand3b_2 _31472_ (.A_N(_09438_),
    .B(_09440_),
    .C(_09441_),
    .Y(_09442_));
 sky130_fd_sc_hd__nand3_2 _31473_ (.A(_09439_),
    .B(_09112_),
    .C(_09442_),
    .Y(_09443_));
 sky130_fd_sc_hd__nand3_2 _31474_ (.A(_09419_),
    .B(_09422_),
    .C(_09434_),
    .Y(_09444_));
 sky130_fd_sc_hd__inv_2 _31475_ (.A(_09444_),
    .Y(_09445_));
 sky130_fd_sc_hd__and2_2 _31476_ (.A(_09423_),
    .B(_09436_),
    .X(_09446_));
 sky130_fd_sc_hd__o22ai_2 _31477_ (.A1(_09445_),
    .A2(_09446_),
    .B1(_09404_),
    .B2(_09407_),
    .Y(_09447_));
 sky130_fd_sc_hd__nand3_2 _31478_ (.A(_09440_),
    .B(_09438_),
    .C(_09441_),
    .Y(_09448_));
 sky130_fd_sc_hd__nand3_2 _31479_ (.A(_09447_),
    .B(_09305_),
    .C(_09448_),
    .Y(_09449_));
 sky130_fd_sc_hd__nor2_2 _31480_ (.A(_09036_),
    .B(_09065_),
    .Y(_09450_));
 sky130_fd_sc_hd__nor2_2 _31481_ (.A(_09033_),
    .B(_09450_),
    .Y(_09451_));
 sky130_fd_sc_hd__nand3_2 _31482_ (.A(_09443_),
    .B(_09449_),
    .C(_09451_),
    .Y(_09452_));
 sky130_fd_sc_hd__o2bb2ai_2 _31483_ (.A1_N(_09449_),
    .A2_N(_09443_),
    .B1(_09033_),
    .B2(_09450_),
    .Y(_09453_));
 sky130_fd_sc_hd__nand3_2 _31484_ (.A(_09380_),
    .B(_09452_),
    .C(_09453_),
    .Y(_09454_));
 sky130_fd_sc_hd__nand2_2 _31485_ (.A(_09453_),
    .B(_09452_),
    .Y(_09455_));
 sky130_fd_sc_hd__nand3_2 _31486_ (.A(_09455_),
    .B(_09374_),
    .C(_09379_),
    .Y(_09456_));
 sky130_fd_sc_hd__a31oi_2 _31487_ (.A1(_09082_),
    .A2(_09142_),
    .A3(_09081_),
    .B1(_09137_),
    .Y(_09457_));
 sky130_fd_sc_hd__nand3_2 _31488_ (.A(_09454_),
    .B(_09456_),
    .C(_09457_),
    .Y(_09458_));
 sky130_fd_sc_hd__nand2_2 _31489_ (.A(_09143_),
    .B(_09136_),
    .Y(_09459_));
 sky130_fd_sc_hd__a21oi_2 _31490_ (.A1(_09443_),
    .A2(_09449_),
    .B1(_09451_),
    .Y(_09460_));
 sky130_fd_sc_hd__and3_2 _31491_ (.A(_09443_),
    .B(_09449_),
    .C(_09451_),
    .X(_09461_));
 sky130_fd_sc_hd__o2bb2ai_2 _31492_ (.A1_N(_09379_),
    .A2_N(_09374_),
    .B1(_09460_),
    .B2(_09461_),
    .Y(_09462_));
 sky130_fd_sc_hd__and3_2 _31493_ (.A(_09447_),
    .B(_09305_),
    .C(_09448_),
    .X(_09463_));
 sky130_fd_sc_hd__nand2_2 _31494_ (.A(_09443_),
    .B(_09451_),
    .Y(_09464_));
 sky130_fd_sc_hd__o2111ai_2 _31495_ (.A1(_09463_),
    .A2(_09464_),
    .B1(_09379_),
    .C1(_09453_),
    .D1(_09374_),
    .Y(_09465_));
 sky130_fd_sc_hd__nand3_2 _31496_ (.A(_09459_),
    .B(_09462_),
    .C(_09465_),
    .Y(_09466_));
 sky130_fd_sc_hd__nand2_2 _31497_ (.A(_09458_),
    .B(_09466_),
    .Y(_09467_));
 sky130_fd_sc_hd__o21ai_2 _31498_ (.A1(_09300_),
    .A2(_09304_),
    .B1(_09467_),
    .Y(_09468_));
 sky130_fd_sc_hd__nand2_2 _31499_ (.A(_09294_),
    .B(_09299_),
    .Y(_09469_));
 sky130_fd_sc_hd__o21ai_2 _31500_ (.A1(_09302_),
    .A2(_09303_),
    .B1(_09301_),
    .Y(_09470_));
 sky130_fd_sc_hd__o2111ai_2 _31501_ (.A1(_09303_),
    .A2(_09469_),
    .B1(_09466_),
    .C1(_09458_),
    .D1(_09470_),
    .Y(_09471_));
 sky130_fd_sc_hd__nand3_2 _31502_ (.A(_09195_),
    .B(_09468_),
    .C(_09471_),
    .Y(_09472_));
 sky130_fd_sc_hd__nand3_2 _31503_ (.A(_09294_),
    .B(_09297_),
    .C(_09299_),
    .Y(_09473_));
 sky130_fd_sc_hd__nand2_2 _31504_ (.A(_09470_),
    .B(_09473_),
    .Y(_09474_));
 sky130_fd_sc_hd__nand3_2 _31505_ (.A(_09474_),
    .B(_09458_),
    .C(_09466_),
    .Y(_09475_));
 sky130_fd_sc_hd__nand3_2 _31506_ (.A(_09467_),
    .B(_09473_),
    .C(_09470_),
    .Y(_09476_));
 sky130_fd_sc_hd__a31oi_2 _31507_ (.A1(_09006_),
    .A2(_09155_),
    .A3(_09002_),
    .B1(_09149_),
    .Y(_09477_));
 sky130_fd_sc_hd__nand3_2 _31508_ (.A(_09475_),
    .B(_09476_),
    .C(_09477_),
    .Y(_09478_));
 sky130_fd_sc_hd__nand2_2 _31509_ (.A(_08941_),
    .B(_08939_),
    .Y(_09479_));
 sky130_fd_sc_hd__nand2_2 _31510_ (.A(_09479_),
    .B(_08942_),
    .Y(_09480_));
 sky130_fd_sc_hd__inv_2 _31511_ (.A(_09480_),
    .Y(_09481_));
 sky130_fd_sc_hd__a21o_2 _31512_ (.A1(_09151_),
    .A2(_09000_),
    .B1(_09481_),
    .X(_09482_));
 sky130_fd_sc_hd__inv_2 _31513_ (.A(_09482_),
    .Y(_09483_));
 sky130_fd_sc_hd__and3_2 _31514_ (.A(_09151_),
    .B(_09000_),
    .C(_09481_),
    .X(_09484_));
 sky130_fd_sc_hd__o2bb2ai_2 _31515_ (.A1_N(_09472_),
    .A2_N(_09478_),
    .B1(_09483_),
    .B2(_09484_),
    .Y(_09485_));
 sky130_fd_sc_hd__nand2_2 _31516_ (.A(_09159_),
    .B(_09157_),
    .Y(_09486_));
 sky130_fd_sc_hd__o22ai_2 _31517_ (.A1(_09162_),
    .A2(_09486_),
    .B1(_09175_),
    .B2(_09160_),
    .Y(_09487_));
 sky130_fd_sc_hd__nor2_2 _31518_ (.A(_09484_),
    .B(_09483_),
    .Y(_09488_));
 sky130_fd_sc_hd__nand3_2 _31519_ (.A(_09488_),
    .B(_09478_),
    .C(_09472_),
    .Y(_09489_));
 sky130_fd_sc_hd__nand3_2 _31520_ (.A(_09485_),
    .B(_09487_),
    .C(_09489_),
    .Y(_09490_));
 sky130_fd_sc_hd__a21oi_2 _31521_ (.A1(_09166_),
    .A2(_09168_),
    .B1(_09164_),
    .Y(_09491_));
 sky130_fd_sc_hd__and2_2 _31522_ (.A(_09151_),
    .B(_09000_),
    .X(_09492_));
 sky130_fd_sc_hd__nor2_2 _31523_ (.A(_09480_),
    .B(_09492_),
    .Y(_09493_));
 sky130_fd_sc_hd__and3_2 _31524_ (.A(_09151_),
    .B(_09000_),
    .C(_09480_),
    .X(_09494_));
 sky130_fd_sc_hd__o2bb2ai_2 _31525_ (.A1_N(_09472_),
    .A2_N(_09478_),
    .B1(_09493_),
    .B2(_09494_),
    .Y(_09495_));
 sky130_fd_sc_hd__o211ai_2 _31526_ (.A1(_09483_),
    .A2(_09484_),
    .B1(_09472_),
    .C1(_09478_),
    .Y(_09496_));
 sky130_fd_sc_hd__nand3_2 _31527_ (.A(_09491_),
    .B(_09495_),
    .C(_09496_),
    .Y(_09497_));
 sky130_fd_sc_hd__nor2_2 _31528_ (.A(_08852_),
    .B(_08711_),
    .Y(_09498_));
 sky130_fd_sc_hd__o2bb2ai_2 _31529_ (.A1_N(_09490_),
    .A2_N(_09497_),
    .B1(_09498_),
    .B2(_08898_),
    .Y(_09499_));
 sky130_fd_sc_hd__nand3_2 _31530_ (.A(_09497_),
    .B(_09490_),
    .C(_08900_),
    .Y(_09500_));
 sky130_fd_sc_hd__nand2_2 _31531_ (.A(_09185_),
    .B(_09172_),
    .Y(_09501_));
 sky130_fd_sc_hd__a21oi_2 _31532_ (.A1(_09499_),
    .A2(_09500_),
    .B1(_09501_),
    .Y(_09502_));
 sky130_fd_sc_hd__inv_2 _31533_ (.A(_08865_),
    .Y(_09503_));
 sky130_fd_sc_hd__a31oi_2 _31534_ (.A1(_09173_),
    .A2(_09174_),
    .A3(_09176_),
    .B1(_09503_),
    .Y(_09504_));
 sky130_fd_sc_hd__o211a_2 _31535_ (.A1(_09184_),
    .A2(_09504_),
    .B1(_09500_),
    .C1(_09499_),
    .X(_09505_));
 sky130_fd_sc_hd__nor2_2 _31536_ (.A(_09502_),
    .B(_09505_),
    .Y(_09506_));
 sky130_fd_sc_hd__and2_2 _31537_ (.A(_09179_),
    .B(_09180_),
    .X(_09507_));
 sky130_fd_sc_hd__o21ai_2 _31538_ (.A1(_09182_),
    .A2(_09507_),
    .B1(_09194_),
    .Y(_09508_));
 sky130_fd_sc_hd__inv_2 _31539_ (.A(_09186_),
    .Y(_09509_));
 sky130_fd_sc_hd__nand2_2 _31540_ (.A(_09508_),
    .B(_09509_),
    .Y(_09510_));
 sky130_fd_sc_hd__xor2_2 _31541_ (.A(_09506_),
    .B(_09510_),
    .X(_02646_));
 sky130_fd_sc_hd__nand2_2 _31542_ (.A(_09469_),
    .B(_09297_),
    .Y(_09511_));
 sky130_fd_sc_hd__inv_2 _31543_ (.A(_09240_),
    .Y(_09512_));
 sky130_fd_sc_hd__inv_2 _31544_ (.A(_09233_),
    .Y(_09513_));
 sky130_fd_sc_hd__o21a_2 _31545_ (.A1(_09512_),
    .A2(_09513_),
    .B1(_09238_),
    .X(_09514_));
 sky130_fd_sc_hd__inv_2 _31546_ (.A(_09514_),
    .Y(_09515_));
 sky130_fd_sc_hd__nand2_2 _31547_ (.A(_09511_),
    .B(_09515_),
    .Y(_09516_));
 sky130_fd_sc_hd__inv_2 _31548_ (.A(_09516_),
    .Y(_09517_));
 sky130_fd_sc_hd__nor2_2 _31549_ (.A(_09515_),
    .B(_09511_),
    .Y(_09518_));
 sky130_fd_sc_hd__nor2_2 _31550_ (.A(_09324_),
    .B(_09321_),
    .Y(_09519_));
 sky130_fd_sc_hd__nand3_2 _31551_ (.A(_19354_),
    .B(_07652_),
    .C(_05910_),
    .Y(_09520_));
 sky130_fd_sc_hd__nand2_2 _31552_ (.A(_07890_),
    .B(_08218_),
    .Y(_09521_));
 sky130_fd_sc_hd__inv_2 _31553_ (.A(_09521_),
    .Y(_09522_));
 sky130_fd_sc_hd__a22o_2 _31554_ (.A1(_07886_),
    .A2(_06540_),
    .B1(_06824_),
    .B2(_06538_),
    .X(_09523_));
 sky130_fd_sc_hd__o211ai_2 _31555_ (.A1(_06391_),
    .A2(_09520_),
    .B1(_09522_),
    .C1(_09523_),
    .Y(_09524_));
 sky130_fd_sc_hd__a22oi_2 _31556_ (.A1(_09018_),
    .A2(_06540_),
    .B1(_09019_),
    .B2(_06726_),
    .Y(_09525_));
 sky130_fd_sc_hd__nor2_2 _31557_ (.A(_06391_),
    .B(_09520_),
    .Y(_09526_));
 sky130_fd_sc_hd__o21ai_2 _31558_ (.A1(_09525_),
    .A2(_09526_),
    .B1(_09521_),
    .Y(_09527_));
 sky130_fd_sc_hd__o211ai_2 _31559_ (.A1(_09323_),
    .A2(_09519_),
    .B1(_09524_),
    .C1(_09527_),
    .Y(_09528_));
 sky130_fd_sc_hd__o21ai_2 _31560_ (.A1(_09525_),
    .A2(_09526_),
    .B1(_09522_),
    .Y(_09529_));
 sky130_fd_sc_hd__a21oi_2 _31561_ (.A1(_09327_),
    .A2(_09325_),
    .B1(_09323_),
    .Y(_09530_));
 sky130_fd_sc_hd__o211ai_2 _31562_ (.A1(_06391_),
    .A2(_09520_),
    .B1(_09521_),
    .C1(_09523_),
    .Y(_09531_));
 sky130_fd_sc_hd__nand3_2 _31563_ (.A(_09529_),
    .B(_09530_),
    .C(_09531_),
    .Y(_09532_));
 sky130_fd_sc_hd__nand2_2 _31564_ (.A(_09528_),
    .B(_09532_),
    .Y(_09533_));
 sky130_fd_sc_hd__a21oi_2 _31565_ (.A1(_09390_),
    .A2(_09388_),
    .B1(_09385_),
    .Y(_09534_));
 sky130_fd_sc_hd__nand2_2 _31566_ (.A(_09533_),
    .B(_09534_),
    .Y(_09535_));
 sky130_fd_sc_hd__nand3b_2 _31567_ (.A_N(_09534_),
    .B(_09528_),
    .C(_09532_),
    .Y(_09536_));
 sky130_fd_sc_hd__nand2_2 _31568_ (.A(_09406_),
    .B(_09396_),
    .Y(_09537_));
 sky130_fd_sc_hd__a21oi_2 _31569_ (.A1(_09535_),
    .A2(_09536_),
    .B1(_09537_),
    .Y(_09538_));
 sky130_fd_sc_hd__a31oi_2 _31570_ (.A1(_09382_),
    .A2(_09389_),
    .A3(_09391_),
    .B1(_09398_),
    .Y(_09539_));
 sky130_fd_sc_hd__o211a_2 _31571_ (.A1(_09405_),
    .A2(_09539_),
    .B1(_09536_),
    .C1(_09535_),
    .X(_09540_));
 sky130_fd_sc_hd__nand2_2 _31572_ (.A(_06278_),
    .B(_07143_),
    .Y(_09541_));
 sky130_fd_sc_hd__nand2_2 _31573_ (.A(_07450_),
    .B(_06560_),
    .Y(_09542_));
 sky130_fd_sc_hd__nor2_2 _31574_ (.A(_09541_),
    .B(_09542_),
    .Y(_09543_));
 sky130_fd_sc_hd__and2_2 _31575_ (.A(_09541_),
    .B(_09542_),
    .X(_09544_));
 sky130_fd_sc_hd__nand2_2 _31576_ (.A(_06446_),
    .B(_06946_),
    .Y(_09545_));
 sky130_fd_sc_hd__inv_2 _31577_ (.A(_09545_),
    .Y(_09546_));
 sky130_fd_sc_hd__o21ai_2 _31578_ (.A1(_09543_),
    .A2(_09544_),
    .B1(_09546_),
    .Y(_09547_));
 sky130_fd_sc_hd__or2_2 _31579_ (.A(_09541_),
    .B(_09542_),
    .X(_09548_));
 sky130_fd_sc_hd__nand2_2 _31580_ (.A(_09541_),
    .B(_09542_),
    .Y(_09549_));
 sky130_fd_sc_hd__nand3_2 _31581_ (.A(_09548_),
    .B(_09549_),
    .C(_09545_),
    .Y(_09550_));
 sky130_fd_sc_hd__a21oi_2 _31582_ (.A1(_09414_),
    .A2(_09417_),
    .B1(_09411_),
    .Y(_09551_));
 sky130_fd_sc_hd__a21o_2 _31583_ (.A1(_09547_),
    .A2(_09550_),
    .B1(_09551_),
    .X(_09552_));
 sky130_fd_sc_hd__nand3_2 _31584_ (.A(_09547_),
    .B(_09550_),
    .C(_09551_),
    .Y(_09553_));
 sky130_fd_sc_hd__nand2_2 _31585_ (.A(_09552_),
    .B(_09553_),
    .Y(_09554_));
 sky130_fd_sc_hd__nand2_2 _31586_ (.A(_05956_),
    .B(_06944_),
    .Y(_09555_));
 sky130_fd_sc_hd__nand2_2 _31587_ (.A(_07034_),
    .B(_08089_),
    .Y(_09556_));
 sky130_fd_sc_hd__nor2_2 _31588_ (.A(_09555_),
    .B(_09556_),
    .Y(_09557_));
 sky130_fd_sc_hd__nand2_2 _31589_ (.A(_09555_),
    .B(_09556_),
    .Y(_09558_));
 sky130_fd_sc_hd__inv_2 _31590_ (.A(_09558_),
    .Y(_09559_));
 sky130_fd_sc_hd__nand2_2 _31591_ (.A(_05673_),
    .B(_07593_),
    .Y(_09560_));
 sky130_fd_sc_hd__inv_2 _31592_ (.A(_09560_),
    .Y(_09561_));
 sky130_fd_sc_hd__o21ai_2 _31593_ (.A1(_09557_),
    .A2(_09559_),
    .B1(_09561_),
    .Y(_09562_));
 sky130_fd_sc_hd__nand3b_2 _31594_ (.A_N(_09557_),
    .B(_09558_),
    .C(_09560_),
    .Y(_09563_));
 sky130_fd_sc_hd__nand2_2 _31595_ (.A(_09562_),
    .B(_09563_),
    .Y(_09564_));
 sky130_fd_sc_hd__inv_2 _31596_ (.A(_09564_),
    .Y(_09565_));
 sky130_fd_sc_hd__nand2_2 _31597_ (.A(_09554_),
    .B(_09565_),
    .Y(_09566_));
 sky130_fd_sc_hd__nand3_2 _31598_ (.A(_09552_),
    .B(_09553_),
    .C(_09564_),
    .Y(_09567_));
 sky130_fd_sc_hd__nand2_2 _31599_ (.A(_09566_),
    .B(_09567_),
    .Y(_09568_));
 sky130_fd_sc_hd__o21ai_2 _31600_ (.A1(_09538_),
    .A2(_09540_),
    .B1(_09568_),
    .Y(_09569_));
 sky130_fd_sc_hd__nand2_2 _31601_ (.A(_09554_),
    .B(_09564_),
    .Y(_09570_));
 sky130_fd_sc_hd__nand3_2 _31602_ (.A(_09565_),
    .B(_09553_),
    .C(_09552_),
    .Y(_09571_));
 sky130_fd_sc_hd__nand2_2 _31603_ (.A(_09570_),
    .B(_09571_),
    .Y(_09572_));
 sky130_fd_sc_hd__a21o_2 _31604_ (.A1(_09535_),
    .A2(_09536_),
    .B1(_09537_),
    .X(_09573_));
 sky130_fd_sc_hd__nand3_2 _31605_ (.A(_09537_),
    .B(_09535_),
    .C(_09536_),
    .Y(_09574_));
 sky130_fd_sc_hd__nand3_2 _31606_ (.A(_09572_),
    .B(_09573_),
    .C(_09574_),
    .Y(_09575_));
 sky130_fd_sc_hd__o21ai_2 _31607_ (.A1(_09370_),
    .A2(_09362_),
    .B1(_09336_),
    .Y(_09576_));
 sky130_fd_sc_hd__nand3_2 _31608_ (.A(_09569_),
    .B(_09575_),
    .C(_09576_),
    .Y(_09577_));
 sky130_fd_sc_hd__o21ai_2 _31609_ (.A1(_09538_),
    .A2(_09540_),
    .B1(_09572_),
    .Y(_09578_));
 sky130_fd_sc_hd__a21oi_2 _31610_ (.A1(_09333_),
    .A2(_09337_),
    .B1(_09369_),
    .Y(_09579_));
 sky130_fd_sc_hd__nand3_2 _31611_ (.A(_09568_),
    .B(_09573_),
    .C(_09574_),
    .Y(_09580_));
 sky130_fd_sc_hd__nand3_2 _31612_ (.A(_09578_),
    .B(_09579_),
    .C(_09580_),
    .Y(_09581_));
 sky130_fd_sc_hd__nor2_2 _31613_ (.A(_09438_),
    .B(_09407_),
    .Y(_09582_));
 sky130_fd_sc_hd__nor2_2 _31614_ (.A(_09404_),
    .B(_09582_),
    .Y(_09583_));
 sky130_fd_sc_hd__a21oi_2 _31615_ (.A1(_09577_),
    .A2(_09581_),
    .B1(_09583_),
    .Y(_09584_));
 sky130_fd_sc_hd__and3_2 _31616_ (.A(_09577_),
    .B(_09581_),
    .C(_09583_),
    .X(_09585_));
 sky130_fd_sc_hd__a21oi_2 _31617_ (.A1(_09344_),
    .A2(_09345_),
    .B1(_09342_),
    .Y(_09586_));
 sky130_fd_sc_hd__nand2_2 _31618_ (.A(_09339_),
    .B(_05323_),
    .Y(_09587_));
 sky130_fd_sc_hd__nand2_2 _31619_ (.A(_19330_),
    .B(_06792_),
    .Y(_09588_));
 sky130_fd_sc_hd__nor2_2 _31620_ (.A(_09587_),
    .B(_09588_),
    .Y(_09589_));
 sky130_fd_sc_hd__and2_2 _31621_ (.A(_09587_),
    .B(_09588_),
    .X(_09590_));
 sky130_fd_sc_hd__nand2_2 _31622_ (.A(_19333_),
    .B(_05212_),
    .Y(_09591_));
 sky130_fd_sc_hd__o21ai_2 _31623_ (.A1(_09589_),
    .A2(_09590_),
    .B1(_09591_),
    .Y(_09592_));
 sky130_fd_sc_hd__or2_2 _31624_ (.A(_09587_),
    .B(_09588_),
    .X(_09593_));
 sky130_fd_sc_hd__nand2_2 _31625_ (.A(_09587_),
    .B(_09588_),
    .Y(_09594_));
 sky130_fd_sc_hd__inv_2 _31626_ (.A(_09591_),
    .Y(_09595_));
 sky130_fd_sc_hd__nand3_2 _31627_ (.A(_09593_),
    .B(_09594_),
    .C(_09595_),
    .Y(_09596_));
 sky130_fd_sc_hd__nand3b_2 _31628_ (.A_N(_09586_),
    .B(_09592_),
    .C(_09596_),
    .Y(_09597_));
 sky130_fd_sc_hd__o21ai_2 _31629_ (.A1(_09589_),
    .A2(_09590_),
    .B1(_09595_),
    .Y(_09598_));
 sky130_fd_sc_hd__nand3_2 _31630_ (.A(_09593_),
    .B(_09594_),
    .C(_09591_),
    .Y(_09599_));
 sky130_fd_sc_hd__nand3_2 _31631_ (.A(_09598_),
    .B(_09599_),
    .C(_09586_),
    .Y(_09600_));
 sky130_fd_sc_hd__nand2_2 _31632_ (.A(_09597_),
    .B(_09600_),
    .Y(_09601_));
 sky130_fd_sc_hd__buf_1 _31633_ (.A(\pcpi_mul.rs2[28] ),
    .X(_09602_));
 sky130_fd_sc_hd__nand2_2 _31634_ (.A(_09602_),
    .B(_05188_),
    .Y(_09603_));
 sky130_fd_sc_hd__nand2_2 _31635_ (.A(_19322_),
    .B(_05190_),
    .Y(_09604_));
 sky130_fd_sc_hd__nor2_2 _31636_ (.A(_09603_),
    .B(_09604_),
    .Y(_09605_));
 sky130_fd_sc_hd__and2_2 _31637_ (.A(_09603_),
    .B(_09604_),
    .X(_09606_));
 sky130_fd_sc_hd__or2_2 _31638_ (.A(_09605_),
    .B(_09606_),
    .X(_09607_));
 sky130_fd_sc_hd__nand2_2 _31639_ (.A(_09601_),
    .B(_09607_),
    .Y(_09608_));
 sky130_fd_sc_hd__inv_2 _31640_ (.A(_09607_),
    .Y(_09609_));
 sky130_fd_sc_hd__nand3_2 _31641_ (.A(_09609_),
    .B(_09600_),
    .C(_09597_),
    .Y(_09610_));
 sky130_fd_sc_hd__nor2_2 _31642_ (.A(_09367_),
    .B(_09355_),
    .Y(_09611_));
 sky130_fd_sc_hd__a21oi_2 _31643_ (.A1(_09608_),
    .A2(_09610_),
    .B1(_09611_),
    .Y(_09612_));
 sky130_fd_sc_hd__and3_2 _31644_ (.A(_09611_),
    .B(_09608_),
    .C(_09610_),
    .X(_09613_));
 sky130_fd_sc_hd__buf_1 _31645_ (.A(\pcpi_mul.rs2[22] ),
    .X(_09614_));
 sky130_fd_sc_hd__nand3_2 _31646_ (.A(_09094_),
    .B(_09614_),
    .C(_19625_),
    .Y(_09615_));
 sky130_fd_sc_hd__nor2_2 _31647_ (.A(_05261_),
    .B(_09615_),
    .Y(_09616_));
 sky130_fd_sc_hd__buf_1 _31648_ (.A(_19339_),
    .X(_09617_));
 sky130_fd_sc_hd__a22o_2 _31649_ (.A1(_08382_),
    .A2(_06502_),
    .B1(_09617_),
    .B2(_05425_),
    .X(_09618_));
 sky130_fd_sc_hd__nand2_2 _31650_ (.A(_08388_),
    .B(_06808_),
    .Y(_09619_));
 sky130_fd_sc_hd__inv_2 _31651_ (.A(_09619_),
    .Y(_09620_));
 sky130_fd_sc_hd__nand2_2 _31652_ (.A(_09618_),
    .B(_09620_),
    .Y(_09621_));
 sky130_fd_sc_hd__a22oi_2 _31653_ (.A1(_08382_),
    .A2(_05341_),
    .B1(_08791_),
    .B2(_05425_),
    .Y(_09622_));
 sky130_fd_sc_hd__o21ai_2 _31654_ (.A1(_09622_),
    .A2(_09616_),
    .B1(_09619_),
    .Y(_09623_));
 sky130_fd_sc_hd__o21bai_2 _31655_ (.A1(_09310_),
    .A2(_09307_),
    .B1_N(_09309_),
    .Y(_09624_));
 sky130_fd_sc_hd__o211ai_2 _31656_ (.A1(_09616_),
    .A2(_09621_),
    .B1(_09623_),
    .C1(_09624_),
    .Y(_09625_));
 sky130_fd_sc_hd__o21ai_2 _31657_ (.A1(_09622_),
    .A2(_09616_),
    .B1(_09620_),
    .Y(_09626_));
 sky130_fd_sc_hd__a21oi_2 _31658_ (.A1(_09314_),
    .A2(_09311_),
    .B1(_09309_),
    .Y(_09627_));
 sky130_fd_sc_hd__o211ai_2 _31659_ (.A1(_05501_),
    .A2(_09615_),
    .B1(_09619_),
    .C1(_09618_),
    .Y(_09628_));
 sky130_fd_sc_hd__nand3_2 _31660_ (.A(_09626_),
    .B(_09627_),
    .C(_09628_),
    .Y(_09629_));
 sky130_fd_sc_hd__nand2_2 _31661_ (.A(_07483_),
    .B(_05506_),
    .Y(_09630_));
 sky130_fd_sc_hd__nand2_2 _31662_ (.A(_07478_),
    .B(_06327_),
    .Y(_09631_));
 sky130_fd_sc_hd__nor2_2 _31663_ (.A(_09630_),
    .B(_09631_),
    .Y(_09632_));
 sky130_fd_sc_hd__and2_2 _31664_ (.A(_09630_),
    .B(_09631_),
    .X(_09633_));
 sky130_fd_sc_hd__nand2_2 _31665_ (.A(_07475_),
    .B(_06889_),
    .Y(_09634_));
 sky130_fd_sc_hd__inv_2 _31666_ (.A(_09634_),
    .Y(_09635_));
 sky130_fd_sc_hd__o21ai_2 _31667_ (.A1(_09632_),
    .A2(_09633_),
    .B1(_09635_),
    .Y(_09636_));
 sky130_fd_sc_hd__nand2_2 _31668_ (.A(_09630_),
    .B(_09631_),
    .Y(_09637_));
 sky130_fd_sc_hd__nand3b_2 _31669_ (.A_N(_09632_),
    .B(_09634_),
    .C(_09637_),
    .Y(_09638_));
 sky130_fd_sc_hd__nand2_2 _31670_ (.A(_09636_),
    .B(_09638_),
    .Y(_09639_));
 sky130_fd_sc_hd__a21oi_2 _31671_ (.A1(_09625_),
    .A2(_09629_),
    .B1(_09639_),
    .Y(_09640_));
 sky130_fd_sc_hd__and3_2 _31672_ (.A(_09625_),
    .B(_09639_),
    .C(_09629_),
    .X(_09641_));
 sky130_fd_sc_hd__o21ai_2 _31673_ (.A1(_09640_),
    .A2(_09641_),
    .B1(_09350_),
    .Y(_09642_));
 sky130_fd_sc_hd__a21o_2 _31674_ (.A1(_09625_),
    .A2(_09629_),
    .B1(_09639_),
    .X(_09643_));
 sky130_fd_sc_hd__inv_2 _31675_ (.A(_09350_),
    .Y(_09644_));
 sky130_fd_sc_hd__nand3_2 _31676_ (.A(_09625_),
    .B(_09639_),
    .C(_09629_),
    .Y(_09645_));
 sky130_fd_sc_hd__nand3_2 _31677_ (.A(_09643_),
    .B(_09644_),
    .C(_09645_),
    .Y(_09646_));
 sky130_fd_sc_hd__nand2_2 _31678_ (.A(_09335_),
    .B(_09320_),
    .Y(_09647_));
 sky130_fd_sc_hd__inv_2 _31679_ (.A(_09647_),
    .Y(_09648_));
 sky130_fd_sc_hd__nand3_2 _31680_ (.A(_09642_),
    .B(_09646_),
    .C(_09648_),
    .Y(_09649_));
 sky130_fd_sc_hd__a21oi_2 _31681_ (.A1(_09643_),
    .A2(_09645_),
    .B1(_09644_),
    .Y(_09650_));
 sky130_fd_sc_hd__nor3_2 _31682_ (.A(_09350_),
    .B(_09640_),
    .C(_09641_),
    .Y(_09651_));
 sky130_fd_sc_hd__o21ai_2 _31683_ (.A1(_09650_),
    .A2(_09651_),
    .B1(_09647_),
    .Y(_09652_));
 sky130_fd_sc_hd__o211ai_2 _31684_ (.A1(_09612_),
    .A2(_09613_),
    .B1(_09649_),
    .C1(_09652_),
    .Y(_09653_));
 sky130_fd_sc_hd__o21ai_2 _31685_ (.A1(_09650_),
    .A2(_09651_),
    .B1(_09648_),
    .Y(_09654_));
 sky130_fd_sc_hd__nand3_2 _31686_ (.A(_09642_),
    .B(_09646_),
    .C(_09647_),
    .Y(_09655_));
 sky130_fd_sc_hd__a21oi_2 _31687_ (.A1(_09601_),
    .A2(_09607_),
    .B1(_09366_),
    .Y(_09656_));
 sky130_fd_sc_hd__a21oi_2 _31688_ (.A1(_09656_),
    .A2(_09610_),
    .B1(_09612_),
    .Y(_09657_));
 sky130_fd_sc_hd__nand3_2 _31689_ (.A(_09654_),
    .B(_09655_),
    .C(_09657_),
    .Y(_09658_));
 sky130_fd_sc_hd__nand3_2 _31690_ (.A(_09653_),
    .B(_09365_),
    .C(_09658_),
    .Y(_09659_));
 sky130_fd_sc_hd__o2bb2ai_2 _31691_ (.A1_N(_09658_),
    .A2_N(_09653_),
    .B1(_09338_),
    .B2(_09364_),
    .Y(_09660_));
 sky130_fd_sc_hd__o211ai_2 _31692_ (.A1(_09584_),
    .A2(_09585_),
    .B1(_09659_),
    .C1(_09660_),
    .Y(_09661_));
 sky130_fd_sc_hd__and3_2 _31693_ (.A(_09377_),
    .B(_09139_),
    .C(_09378_),
    .X(_09662_));
 sky130_fd_sc_hd__a31oi_2 _31694_ (.A1(_09374_),
    .A2(_09452_),
    .A3(_09453_),
    .B1(_09662_),
    .Y(_09663_));
 sky130_fd_sc_hd__nand2_2 _31695_ (.A(_09660_),
    .B(_09659_),
    .Y(_09664_));
 sky130_fd_sc_hd__nand3_2 _31696_ (.A(_09577_),
    .B(_09581_),
    .C(_09583_),
    .Y(_09665_));
 sky130_fd_sc_hd__o2bb2ai_2 _31697_ (.A1_N(_09577_),
    .A2_N(_09581_),
    .B1(_09404_),
    .B2(_09582_),
    .Y(_09666_));
 sky130_fd_sc_hd__nand3_2 _31698_ (.A(_09664_),
    .B(_09665_),
    .C(_09666_),
    .Y(_09667_));
 sky130_fd_sc_hd__nand3_2 _31699_ (.A(_09661_),
    .B(_09663_),
    .C(_09667_),
    .Y(_09668_));
 sky130_fd_sc_hd__nand3_2 _31700_ (.A(_09374_),
    .B(_09453_),
    .C(_09452_),
    .Y(_09669_));
 sky130_fd_sc_hd__nand2_2 _31701_ (.A(_09669_),
    .B(_09379_),
    .Y(_09670_));
 sky130_fd_sc_hd__o2bb2ai_2 _31702_ (.A1_N(_09659_),
    .A2_N(_09660_),
    .B1(_09584_),
    .B2(_09585_),
    .Y(_09671_));
 sky130_fd_sc_hd__and3_2 _31703_ (.A(_09569_),
    .B(_09575_),
    .C(_09576_),
    .X(_09672_));
 sky130_fd_sc_hd__nand2_2 _31704_ (.A(_09581_),
    .B(_09583_),
    .Y(_09673_));
 sky130_fd_sc_hd__o2111ai_2 _31705_ (.A1(_09672_),
    .A2(_09673_),
    .B1(_09659_),
    .C1(_09666_),
    .D1(_09660_),
    .Y(_09674_));
 sky130_fd_sc_hd__nand3_2 _31706_ (.A(_09670_),
    .B(_09671_),
    .C(_09674_),
    .Y(_09675_));
 sky130_fd_sc_hd__nand2_2 _31707_ (.A(_09668_),
    .B(_09675_),
    .Y(_09676_));
 sky130_fd_sc_hd__inv_2 _31708_ (.A(\pcpi_mul.rs1[21] ),
    .Y(_09677_));
 sky130_fd_sc_hd__buf_1 _31709_ (.A(_09677_),
    .X(_09678_));
 sky130_fd_sc_hd__buf_1 _31710_ (.A(_09678_),
    .X(_09679_));
 sky130_fd_sc_hd__nand3_2 _31711_ (.A(_05448_),
    .B(_05445_),
    .C(_07594_),
    .Y(_09680_));
 sky130_fd_sc_hd__nand2_2 _31712_ (.A(_08953_),
    .B(_19574_),
    .Y(_09681_));
 sky130_fd_sc_hd__a22oi_2 _31713_ (.A1(_07797_),
    .A2(_08650_),
    .B1(_08949_),
    .B2(_07849_),
    .Y(_09682_));
 sky130_fd_sc_hd__nor2_2 _31714_ (.A(_09681_),
    .B(_09682_),
    .Y(_09683_));
 sky130_fd_sc_hd__o21ai_2 _31715_ (.A1(_09679_),
    .A2(_09680_),
    .B1(_09683_),
    .Y(_09684_));
 sky130_fd_sc_hd__a21o_2 _31716_ (.A1(_09432_),
    .A2(_09428_),
    .B1(_09431_),
    .X(_09685_));
 sky130_fd_sc_hd__nor2_2 _31717_ (.A(_09678_),
    .B(_09680_),
    .Y(_09686_));
 sky130_fd_sc_hd__o21ai_2 _31718_ (.A1(_09682_),
    .A2(_09686_),
    .B1(_09681_),
    .Y(_09687_));
 sky130_fd_sc_hd__nand3_2 _31719_ (.A(_09684_),
    .B(_09685_),
    .C(_09687_),
    .Y(_09688_));
 sky130_fd_sc_hd__a22o_2 _31720_ (.A1(_08948_),
    .A2(_08108_),
    .B1(_09254_),
    .B2(_19578_),
    .X(_09689_));
 sky130_fd_sc_hd__nand3b_2 _31721_ (.A_N(_09686_),
    .B(_09681_),
    .C(_09689_),
    .Y(_09690_));
 sky130_fd_sc_hd__a21oi_2 _31722_ (.A1(_09432_),
    .A2(_09428_),
    .B1(_09431_),
    .Y(_09691_));
 sky130_fd_sc_hd__o21bai_2 _31723_ (.A1(_09682_),
    .A2(_09686_),
    .B1_N(_09681_),
    .Y(_09692_));
 sky130_fd_sc_hd__nand3_2 _31724_ (.A(_09690_),
    .B(_09691_),
    .C(_09692_),
    .Y(_09693_));
 sky130_fd_sc_hd__a21o_2 _31725_ (.A1(_09252_),
    .A2(_09258_),
    .B1(_09257_),
    .X(_09694_));
 sky130_fd_sc_hd__a21o_2 _31726_ (.A1(_09688_),
    .A2(_09693_),
    .B1(_09694_),
    .X(_09695_));
 sky130_fd_sc_hd__nand3_2 _31727_ (.A(_09688_),
    .B(_09693_),
    .C(_09694_),
    .Y(_09696_));
 sky130_fd_sc_hd__nand2_2 _31728_ (.A(_09419_),
    .B(_09434_),
    .Y(_09697_));
 sky130_fd_sc_hd__nand2_2 _31729_ (.A(_09697_),
    .B(_09422_),
    .Y(_09698_));
 sky130_fd_sc_hd__a21oi_2 _31730_ (.A1(_09695_),
    .A2(_09696_),
    .B1(_09698_),
    .Y(_09699_));
 sky130_fd_sc_hd__inv_2 _31731_ (.A(_09688_),
    .Y(_09700_));
 sky130_fd_sc_hd__nand2_2 _31732_ (.A(_09693_),
    .B(_09694_),
    .Y(_09701_));
 sky130_fd_sc_hd__o211a_2 _31733_ (.A1(_09700_),
    .A2(_09701_),
    .B1(_09695_),
    .C1(_09698_),
    .X(_09702_));
 sky130_fd_sc_hd__nand2_2 _31734_ (.A(_09274_),
    .B(_09265_),
    .Y(_09703_));
 sky130_fd_sc_hd__o21ai_2 _31735_ (.A1(_09699_),
    .A2(_09702_),
    .B1(_09703_),
    .Y(_09704_));
 sky130_fd_sc_hd__a21oi_2 _31736_ (.A1(_09278_),
    .A2(_09279_),
    .B1(_09275_),
    .Y(_09705_));
 sky130_fd_sc_hd__a21o_2 _31737_ (.A1(_09695_),
    .A2(_09696_),
    .B1(_09698_),
    .X(_09706_));
 sky130_fd_sc_hd__inv_2 _31738_ (.A(_09703_),
    .Y(_09707_));
 sky130_fd_sc_hd__nand3_2 _31739_ (.A(_09698_),
    .B(_09695_),
    .C(_09696_),
    .Y(_09708_));
 sky130_fd_sc_hd__nand3_2 _31740_ (.A(_09706_),
    .B(_09707_),
    .C(_09708_),
    .Y(_09709_));
 sky130_fd_sc_hd__nand3_2 _31741_ (.A(_09704_),
    .B(_09705_),
    .C(_09709_),
    .Y(_09710_));
 sky130_fd_sc_hd__o21ai_2 _31742_ (.A1(_09699_),
    .A2(_09702_),
    .B1(_09707_),
    .Y(_09711_));
 sky130_fd_sc_hd__nand3_2 _31743_ (.A(_09706_),
    .B(_09703_),
    .C(_09708_),
    .Y(_09712_));
 sky130_fd_sc_hd__o21ai_2 _31744_ (.A1(_09280_),
    .A2(_09272_),
    .B1(_09281_),
    .Y(_09713_));
 sky130_fd_sc_hd__nand3_2 _31745_ (.A(_09711_),
    .B(_09712_),
    .C(_09713_),
    .Y(_09714_));
 sky130_fd_sc_hd__nand2_2 _31746_ (.A(_09710_),
    .B(_09714_),
    .Y(_09715_));
 sky130_fd_sc_hd__o21ai_2 _31747_ (.A1(_09225_),
    .A2(_09227_),
    .B1(_09215_),
    .Y(_09716_));
 sky130_fd_sc_hd__a21oi_2 _31748_ (.A1(_09205_),
    .A2(_09208_),
    .B1(_09201_),
    .Y(_09717_));
 sky130_fd_sc_hd__nand2_2 _31749_ (.A(_05402_),
    .B(_09199_),
    .Y(_09718_));
 sky130_fd_sc_hd__nand2_2 _31750_ (.A(_06054_),
    .B(_19567_),
    .Y(_09719_));
 sky130_fd_sc_hd__nor2_2 _31751_ (.A(_09718_),
    .B(_09719_),
    .Y(_09720_));
 sky130_fd_sc_hd__and2_2 _31752_ (.A(_09718_),
    .B(_09719_),
    .X(_09721_));
 sky130_fd_sc_hd__buf_1 _31753_ (.A(_19552_),
    .X(_09722_));
 sky130_fd_sc_hd__nand2_2 _31754_ (.A(_06057_),
    .B(_09722_),
    .Y(_09723_));
 sky130_fd_sc_hd__o21ai_2 _31755_ (.A1(_09720_),
    .A2(_09721_),
    .B1(_09723_),
    .Y(_09724_));
 sky130_fd_sc_hd__or2_2 _31756_ (.A(_09718_),
    .B(_09719_),
    .X(_09725_));
 sky130_fd_sc_hd__inv_2 _31757_ (.A(_09723_),
    .Y(_09726_));
 sky130_fd_sc_hd__nand2_2 _31758_ (.A(_09718_),
    .B(_09719_),
    .Y(_09727_));
 sky130_fd_sc_hd__nand3_2 _31759_ (.A(_09725_),
    .B(_09726_),
    .C(_09727_),
    .Y(_09728_));
 sky130_fd_sc_hd__nand3b_2 _31760_ (.A_N(_09717_),
    .B(_09724_),
    .C(_09728_),
    .Y(_09729_));
 sky130_fd_sc_hd__o21ai_2 _31761_ (.A1(_09720_),
    .A2(_09721_),
    .B1(_09726_),
    .Y(_09730_));
 sky130_fd_sc_hd__nand3_2 _31762_ (.A(_09725_),
    .B(_09723_),
    .C(_09727_),
    .Y(_09731_));
 sky130_fd_sc_hd__nand3_2 _31763_ (.A(_09730_),
    .B(_09731_),
    .C(_09717_),
    .Y(_09732_));
 sky130_fd_sc_hd__buf_1 _31764_ (.A(_09203_),
    .X(_09733_));
 sky130_fd_sc_hd__nand2_2 _31765_ (.A(_05123_),
    .B(_08905_),
    .Y(_09734_));
 sky130_fd_sc_hd__a21o_2 _31766_ (.A1(_06220_),
    .A2(_09733_),
    .B1(_09734_),
    .X(_09735_));
 sky130_fd_sc_hd__buf_1 _31767_ (.A(_19557_),
    .X(_09736_));
 sky130_fd_sc_hd__nand2_2 _31768_ (.A(_05118_),
    .B(_09736_),
    .Y(_09737_));
 sky130_fd_sc_hd__a21o_2 _31769_ (.A1(_06219_),
    .A2(_19562_),
    .B1(_09737_),
    .X(_09738_));
 sky130_fd_sc_hd__nand2_2 _31770_ (.A(_19394_),
    .B(_09219_),
    .Y(_09739_));
 sky130_fd_sc_hd__a21oi_2 _31771_ (.A1(_09735_),
    .A2(_09738_),
    .B1(_09739_),
    .Y(_09740_));
 sky130_fd_sc_hd__and3_2 _31772_ (.A(_09735_),
    .B(_09738_),
    .C(_09739_),
    .X(_09741_));
 sky130_fd_sc_hd__nor2_2 _31773_ (.A(_09740_),
    .B(_09741_),
    .Y(_09742_));
 sky130_fd_sc_hd__a21oi_2 _31774_ (.A1(_09729_),
    .A2(_09732_),
    .B1(_09742_),
    .Y(_09743_));
 sky130_fd_sc_hd__and3_2 _31775_ (.A(_09742_),
    .B(_09729_),
    .C(_09732_),
    .X(_09744_));
 sky130_fd_sc_hd__o2bb2ai_2 _31776_ (.A1_N(_09211_),
    .A2_N(_09716_),
    .B1(_09743_),
    .B2(_09744_),
    .Y(_09745_));
 sky130_fd_sc_hd__a21bo_2 _31777_ (.A1(_09211_),
    .A2(_09228_),
    .B1_N(_09215_),
    .X(_09746_));
 sky130_fd_sc_hd__nand3_2 _31778_ (.A(_09742_),
    .B(_09729_),
    .C(_09732_),
    .Y(_09747_));
 sky130_fd_sc_hd__nand3b_2 _31779_ (.A_N(_09743_),
    .B(_09746_),
    .C(_09747_),
    .Y(_09748_));
 sky130_fd_sc_hd__inv_2 _31780_ (.A(_09225_),
    .Y(_09749_));
 sky130_fd_sc_hd__nor2_2 _31781_ (.A(_09217_),
    .B(_09221_),
    .Y(_09750_));
 sky130_fd_sc_hd__inv_2 _31782_ (.A(_09750_),
    .Y(_09751_));
 sky130_fd_sc_hd__nand2_2 _31783_ (.A(_09749_),
    .B(_09751_),
    .Y(_09752_));
 sky130_fd_sc_hd__a21oi_2 _31784_ (.A1(_09745_),
    .A2(_09748_),
    .B1(_09752_),
    .Y(_09753_));
 sky130_fd_sc_hd__and3_2 _31785_ (.A(_09745_),
    .B(_09748_),
    .C(_09752_),
    .X(_09754_));
 sky130_fd_sc_hd__nor2_2 _31786_ (.A(_09753_),
    .B(_09754_),
    .Y(_09755_));
 sky130_fd_sc_hd__nand2_2 _31787_ (.A(_09715_),
    .B(_09755_),
    .Y(_09756_));
 sky130_fd_sc_hd__a21oi_2 _31788_ (.A1(_09443_),
    .A2(_09451_),
    .B1(_09463_),
    .Y(_09757_));
 sky130_fd_sc_hd__a21o_2 _31789_ (.A1(_09745_),
    .A2(_09748_),
    .B1(_09752_),
    .X(_09758_));
 sky130_fd_sc_hd__nand3_2 _31790_ (.A(_09745_),
    .B(_09752_),
    .C(_09748_),
    .Y(_09759_));
 sky130_fd_sc_hd__nand2_2 _31791_ (.A(_09758_),
    .B(_09759_),
    .Y(_09760_));
 sky130_fd_sc_hd__nand3_2 _31792_ (.A(_09760_),
    .B(_09714_),
    .C(_09710_),
    .Y(_09761_));
 sky130_fd_sc_hd__nand3_2 _31793_ (.A(_09756_),
    .B(_09757_),
    .C(_09761_),
    .Y(_09762_));
 sky130_fd_sc_hd__nand2_2 _31794_ (.A(_09715_),
    .B(_09760_),
    .Y(_09763_));
 sky130_fd_sc_hd__nand3_2 _31795_ (.A(_09755_),
    .B(_09714_),
    .C(_09710_),
    .Y(_09764_));
 sky130_fd_sc_hd__nand2_2 _31796_ (.A(_09464_),
    .B(_09449_),
    .Y(_09765_));
 sky130_fd_sc_hd__nand3_2 _31797_ (.A(_09763_),
    .B(_09764_),
    .C(_09765_),
    .Y(_09766_));
 sky130_fd_sc_hd__inv_2 _31798_ (.A(_09283_),
    .Y(_09767_));
 sky130_fd_sc_hd__inv_2 _31799_ (.A(_09287_),
    .Y(_09768_));
 sky130_fd_sc_hd__nor2_2 _31800_ (.A(_09243_),
    .B(_09768_),
    .Y(_09769_));
 sky130_fd_sc_hd__o2bb2ai_2 _31801_ (.A1_N(_09762_),
    .A2_N(_09766_),
    .B1(_09767_),
    .B2(_09769_),
    .Y(_09770_));
 sky130_fd_sc_hd__nor2_2 _31802_ (.A(_09767_),
    .B(_09769_),
    .Y(_09771_));
 sky130_fd_sc_hd__nand3_2 _31803_ (.A(_09771_),
    .B(_09762_),
    .C(_09766_),
    .Y(_09772_));
 sky130_fd_sc_hd__nand2_2 _31804_ (.A(_09770_),
    .B(_09772_),
    .Y(_09773_));
 sky130_fd_sc_hd__nand2_2 _31805_ (.A(_09676_),
    .B(_09773_),
    .Y(_09774_));
 sky130_fd_sc_hd__and3_2 _31806_ (.A(_09763_),
    .B(_09764_),
    .C(_09765_),
    .X(_09775_));
 sky130_fd_sc_hd__nand2_2 _31807_ (.A(_09771_),
    .B(_09762_),
    .Y(_09776_));
 sky130_fd_sc_hd__o2111ai_2 _31808_ (.A1(_09775_),
    .A2(_09776_),
    .B1(_09675_),
    .C1(_09770_),
    .D1(_09668_),
    .Y(_09777_));
 sky130_fd_sc_hd__nand3_2 _31809_ (.A(_09470_),
    .B(_09458_),
    .C(_09473_),
    .Y(_09778_));
 sky130_fd_sc_hd__nand2_2 _31810_ (.A(_09778_),
    .B(_09466_),
    .Y(_09779_));
 sky130_fd_sc_hd__a21oi_2 _31811_ (.A1(_09774_),
    .A2(_09777_),
    .B1(_09779_),
    .Y(_09780_));
 sky130_fd_sc_hd__nand2_2 _31812_ (.A(_09668_),
    .B(_09770_),
    .Y(_09781_));
 sky130_fd_sc_hd__nand2_2 _31813_ (.A(_09675_),
    .B(_09772_),
    .Y(_09782_));
 sky130_fd_sc_hd__o211a_2 _31814_ (.A1(_09781_),
    .A2(_09782_),
    .B1(_09774_),
    .C1(_09779_),
    .X(_09783_));
 sky130_fd_sc_hd__o22ai_2 _31815_ (.A1(_09517_),
    .A2(_09518_),
    .B1(_09780_),
    .B2(_09783_),
    .Y(_09784_));
 sky130_fd_sc_hd__nand2_2 _31816_ (.A(_09488_),
    .B(_09478_),
    .Y(_09785_));
 sky130_fd_sc_hd__nand2_2 _31817_ (.A(_09785_),
    .B(_09472_),
    .Y(_09786_));
 sky130_fd_sc_hd__nand2_2 _31818_ (.A(_09774_),
    .B(_09777_),
    .Y(_09787_));
 sky130_fd_sc_hd__and2_2 _31819_ (.A(_09778_),
    .B(_09466_),
    .X(_09788_));
 sky130_fd_sc_hd__nand2_2 _31820_ (.A(_09787_),
    .B(_09788_),
    .Y(_09789_));
 sky130_fd_sc_hd__nand3_2 _31821_ (.A(_09779_),
    .B(_09774_),
    .C(_09777_),
    .Y(_09790_));
 sky130_fd_sc_hd__inv_2 _31822_ (.A(_09511_),
    .Y(_09791_));
 sky130_fd_sc_hd__nand2_2 _31823_ (.A(_09791_),
    .B(_09515_),
    .Y(_09792_));
 sky130_fd_sc_hd__nand2_2 _31824_ (.A(_09511_),
    .B(_09514_),
    .Y(_09793_));
 sky130_fd_sc_hd__nand2_2 _31825_ (.A(_09792_),
    .B(_09793_),
    .Y(_09794_));
 sky130_fd_sc_hd__nand3_2 _31826_ (.A(_09789_),
    .B(_09790_),
    .C(_09794_),
    .Y(_09795_));
 sky130_fd_sc_hd__nand3_2 _31827_ (.A(_09784_),
    .B(_09786_),
    .C(_09795_),
    .Y(_09796_));
 sky130_fd_sc_hd__o21ai_2 _31828_ (.A1(_09780_),
    .A2(_09783_),
    .B1(_09794_),
    .Y(_09797_));
 sky130_fd_sc_hd__a21boi_2 _31829_ (.A1(_09488_),
    .A2(_09478_),
    .B1_N(_09472_),
    .Y(_09798_));
 sky130_fd_sc_hd__or2b_2 _31830_ (.A(_09518_),
    .B_N(_09516_),
    .X(_09799_));
 sky130_fd_sc_hd__nand3_2 _31831_ (.A(_09789_),
    .B(_09790_),
    .C(_09799_),
    .Y(_09800_));
 sky130_fd_sc_hd__nand3_2 _31832_ (.A(_09797_),
    .B(_09798_),
    .C(_09800_),
    .Y(_09801_));
 sky130_fd_sc_hd__o2bb2ai_2 _31833_ (.A1_N(_09796_),
    .A2_N(_09801_),
    .B1(_09492_),
    .B2(_09481_),
    .Y(_09802_));
 sky130_fd_sc_hd__nand3_2 _31834_ (.A(_09801_),
    .B(_09796_),
    .C(_09483_),
    .Y(_09803_));
 sky130_fd_sc_hd__a21bo_2 _31835_ (.A1(_08900_),
    .A2(_09497_),
    .B1_N(_09490_),
    .X(_09804_));
 sky130_fd_sc_hd__a21o_2 _31836_ (.A1(_09802_),
    .A2(_09803_),
    .B1(_09804_),
    .X(_09805_));
 sky130_fd_sc_hd__nand3_2 _31837_ (.A(_09804_),
    .B(_09802_),
    .C(_09803_),
    .Y(_09806_));
 sky130_fd_sc_hd__nand2_2 _31838_ (.A(_09805_),
    .B(_09806_),
    .Y(_09807_));
 sky130_fd_sc_hd__inv_2 _31839_ (.A(_09505_),
    .Y(_09808_));
 sky130_fd_sc_hd__nand3_2 _31840_ (.A(_09187_),
    .B(_09506_),
    .C(_09193_),
    .Y(_09809_));
 sky130_fd_sc_hd__o211ai_2 _31841_ (.A1(_09509_),
    .A2(_09502_),
    .B1(_09808_),
    .C1(_09809_),
    .Y(_09810_));
 sky130_fd_sc_hd__nand3_2 _31842_ (.A(_09191_),
    .B(_09187_),
    .C(_09506_),
    .Y(_09811_));
 sky130_fd_sc_hd__a21oi_2 _31843_ (.A1(_08583_),
    .A2(_08588_),
    .B1(_09811_),
    .Y(_09812_));
 sky130_fd_sc_hd__nor2_2 _31844_ (.A(_09810_),
    .B(_09812_),
    .Y(_09813_));
 sky130_fd_sc_hd__xor2_2 _31845_ (.A(_09807_),
    .B(_09813_),
    .X(_02647_));
 sky130_fd_sc_hd__nand3_2 _31846_ (.A(_09668_),
    .B(_09770_),
    .C(_09772_),
    .Y(_09814_));
 sky130_fd_sc_hd__nand2_2 _31847_ (.A(_09814_),
    .B(_09675_),
    .Y(_09815_));
 sky130_fd_sc_hd__and3_2 _31848_ (.A(_09653_),
    .B(_09365_),
    .C(_09658_),
    .X(_09816_));
 sky130_fd_sc_hd__a31o_2 _31849_ (.A1(_09660_),
    .A2(_09666_),
    .A3(_09665_),
    .B1(_09816_),
    .X(_09817_));
 sky130_fd_sc_hd__a31oi_2 _31850_ (.A1(_09654_),
    .A2(_09657_),
    .A3(_09655_),
    .B1(_09613_),
    .Y(_09818_));
 sky130_fd_sc_hd__buf_1 _31851_ (.A(\pcpi_mul.rs2[26] ),
    .X(_09819_));
 sky130_fd_sc_hd__a22oi_2 _31852_ (.A1(_09819_),
    .A2(_05330_),
    .B1(_19331_),
    .B2(_06501_),
    .Y(_09820_));
 sky130_fd_sc_hd__nand3_2 _31853_ (.A(_09339_),
    .B(_19330_),
    .C(_06792_),
    .Y(_09821_));
 sky130_fd_sc_hd__nor2_2 _31854_ (.A(_06105_),
    .B(_09821_),
    .Y(_09822_));
 sky130_fd_sc_hd__nand2_2 _31855_ (.A(\pcpi_mul.rs2[24] ),
    .B(_05184_),
    .Y(_09823_));
 sky130_fd_sc_hd__inv_2 _31856_ (.A(_09823_),
    .Y(_09824_));
 sky130_fd_sc_hd__o21ai_2 _31857_ (.A1(_09820_),
    .A2(_09822_),
    .B1(_09824_),
    .Y(_09825_));
 sky130_fd_sc_hd__buf_1 _31858_ (.A(\pcpi_mul.rs2[26] ),
    .X(_09826_));
 sky130_fd_sc_hd__buf_1 _31859_ (.A(\pcpi_mul.rs2[25] ),
    .X(_09827_));
 sky130_fd_sc_hd__a22o_2 _31860_ (.A1(_09826_),
    .A2(_19630_),
    .B1(_09827_),
    .B2(_06629_),
    .X(_09828_));
 sky130_fd_sc_hd__o211ai_2 _31861_ (.A1(_05850_),
    .A2(_09821_),
    .B1(_09823_),
    .C1(_09828_),
    .Y(_09829_));
 sky130_fd_sc_hd__nand3b_2 _31862_ (.A_N(_09605_),
    .B(_09825_),
    .C(_09829_),
    .Y(_09830_));
 sky130_fd_sc_hd__o21ai_2 _31863_ (.A1(_09820_),
    .A2(_09822_),
    .B1(_09823_),
    .Y(_09831_));
 sky130_fd_sc_hd__o211ai_2 _31864_ (.A1(_05850_),
    .A2(_09821_),
    .B1(_09824_),
    .C1(_09828_),
    .Y(_09832_));
 sky130_fd_sc_hd__nand3_2 _31865_ (.A(_09831_),
    .B(_09605_),
    .C(_09832_),
    .Y(_09833_));
 sky130_fd_sc_hd__a21o_2 _31866_ (.A1(_09595_),
    .A2(_09594_),
    .B1(_09589_),
    .X(_09834_));
 sky130_fd_sc_hd__a21o_2 _31867_ (.A1(_09830_),
    .A2(_09833_),
    .B1(_09834_),
    .X(_09835_));
 sky130_fd_sc_hd__nand3_2 _31868_ (.A(_09830_),
    .B(_09833_),
    .C(_09834_),
    .Y(_09836_));
 sky130_fd_sc_hd__nand2_2 _31869_ (.A(_19323_),
    .B(_08393_),
    .Y(_09837_));
 sky130_fd_sc_hd__buf_1 _31870_ (.A(_19319_),
    .X(_09838_));
 sky130_fd_sc_hd__a22oi_2 _31871_ (.A1(_19316_),
    .A2(_05805_),
    .B1(_09838_),
    .B2(_05804_),
    .Y(_09839_));
 sky130_fd_sc_hd__nand2_2 _31872_ (.A(_09602_),
    .B(_05543_),
    .Y(_09840_));
 sky130_fd_sc_hd__buf_2 _31873_ (.A(\pcpi_mul.rs2[29] ),
    .X(_09841_));
 sky130_fd_sc_hd__buf_1 _31874_ (.A(_09841_),
    .X(_09842_));
 sky130_fd_sc_hd__nand2_2 _31875_ (.A(_09842_),
    .B(_19640_),
    .Y(_09843_));
 sky130_fd_sc_hd__nor2_2 _31876_ (.A(_09840_),
    .B(_09843_),
    .Y(_09844_));
 sky130_fd_sc_hd__nor2_2 _31877_ (.A(_09839_),
    .B(_09844_),
    .Y(_09845_));
 sky130_fd_sc_hd__xnor2_2 _31878_ (.A(_09837_),
    .B(_09845_),
    .Y(_09846_));
 sky130_fd_sc_hd__a21oi_2 _31879_ (.A1(_09835_),
    .A2(_09836_),
    .B1(_09846_),
    .Y(_09847_));
 sky130_fd_sc_hd__and3_2 _31880_ (.A(_09835_),
    .B(_09846_),
    .C(_09836_),
    .X(_09848_));
 sky130_fd_sc_hd__o22ai_2 _31881_ (.A1(_09601_),
    .A2(_09607_),
    .B1(_09847_),
    .B2(_09848_),
    .Y(_09849_));
 sky130_fd_sc_hd__nand2_2 _31882_ (.A(_09835_),
    .B(_09836_),
    .Y(_09850_));
 sky130_fd_sc_hd__xor2_2 _31883_ (.A(_09837_),
    .B(_09845_),
    .X(_09851_));
 sky130_fd_sc_hd__nand2_2 _31884_ (.A(_09850_),
    .B(_09851_),
    .Y(_09852_));
 sky130_fd_sc_hd__a21oi_2 _31885_ (.A1(_09830_),
    .A2(_09833_),
    .B1(_09834_),
    .Y(_09853_));
 sky130_fd_sc_hd__nor2_2 _31886_ (.A(_09851_),
    .B(_09853_),
    .Y(_09854_));
 sky130_fd_sc_hd__nand2_2 _31887_ (.A(_09854_),
    .B(_09836_),
    .Y(_09855_));
 sky130_fd_sc_hd__inv_2 _31888_ (.A(_09610_),
    .Y(_09856_));
 sky130_fd_sc_hd__nand3_2 _31889_ (.A(_09852_),
    .B(_09855_),
    .C(_09856_),
    .Y(_09857_));
 sky130_fd_sc_hd__nand2_2 _31890_ (.A(_09849_),
    .B(_09857_),
    .Y(_09858_));
 sky130_fd_sc_hd__a22oi_2 _31891_ (.A1(_08790_),
    .A2(_05343_),
    .B1(_08791_),
    .B2(_06617_),
    .Y(_09859_));
 sky130_fd_sc_hd__nand3_2 _31892_ (.A(_09094_),
    .B(_09614_),
    .C(_19622_),
    .Y(_09860_));
 sky130_fd_sc_hd__nor2_2 _31893_ (.A(_06332_),
    .B(_09860_),
    .Y(_09861_));
 sky130_fd_sc_hd__nand2_2 _31894_ (.A(_19342_),
    .B(_05506_),
    .Y(_09862_));
 sky130_fd_sc_hd__inv_2 _31895_ (.A(_09862_),
    .Y(_09863_));
 sky130_fd_sc_hd__o21ai_2 _31896_ (.A1(_09859_),
    .A2(_09861_),
    .B1(_09863_),
    .Y(_09864_));
 sky130_fd_sc_hd__a21oi_2 _31897_ (.A1(_09618_),
    .A2(_09620_),
    .B1(_09616_),
    .Y(_09865_));
 sky130_fd_sc_hd__a22o_2 _31898_ (.A1(_08790_),
    .A2(_05425_),
    .B1(_08791_),
    .B2(_06617_),
    .X(_09866_));
 sky130_fd_sc_hd__o211ai_2 _31899_ (.A1(_06333_),
    .A2(_09860_),
    .B1(_09862_),
    .C1(_09866_),
    .Y(_09867_));
 sky130_fd_sc_hd__nand3_2 _31900_ (.A(_09864_),
    .B(_09865_),
    .C(_09867_),
    .Y(_09868_));
 sky130_fd_sc_hd__nand2_2 _31901_ (.A(_09866_),
    .B(_09863_),
    .Y(_09869_));
 sky130_fd_sc_hd__o22ai_2 _31902_ (.A1(_05501_),
    .A2(_09615_),
    .B1(_09619_),
    .B2(_09622_),
    .Y(_09870_));
 sky130_fd_sc_hd__o21ai_2 _31903_ (.A1(_09859_),
    .A2(_09861_),
    .B1(_09862_),
    .Y(_09871_));
 sky130_fd_sc_hd__o211ai_2 _31904_ (.A1(_09861_),
    .A2(_09869_),
    .B1(_09870_),
    .C1(_09871_),
    .Y(_09872_));
 sky130_fd_sc_hd__nand2_2 _31905_ (.A(_08407_),
    .B(_05717_),
    .Y(_09873_));
 sky130_fd_sc_hd__a22oi_2 _31906_ (.A1(_09101_),
    .A2(_05737_),
    .B1(_08809_),
    .B2(_09010_),
    .Y(_09874_));
 sky130_fd_sc_hd__nand3_2 _31907_ (.A(_07722_),
    .B(_07478_),
    .C(_06327_),
    .Y(_09875_));
 sky130_fd_sc_hd__nor2_2 _31908_ (.A(_06694_),
    .B(_09875_),
    .Y(_09876_));
 sky130_fd_sc_hd__nor3_2 _31909_ (.A(_09873_),
    .B(_09874_),
    .C(_09876_),
    .Y(_09877_));
 sky130_fd_sc_hd__o21a_2 _31910_ (.A1(_09874_),
    .A2(_09876_),
    .B1(_09873_),
    .X(_09878_));
 sky130_fd_sc_hd__o2bb2ai_2 _31911_ (.A1_N(_09868_),
    .A2_N(_09872_),
    .B1(_09877_),
    .B2(_09878_),
    .Y(_09879_));
 sky130_fd_sc_hd__a22o_2 _31912_ (.A1(_08808_),
    .A2(_05737_),
    .B1(_08809_),
    .B2(_09010_),
    .X(_09880_));
 sky130_fd_sc_hd__nand3b_2 _31913_ (.A_N(_09876_),
    .B(_09880_),
    .C(_09873_),
    .Y(_09881_));
 sky130_fd_sc_hd__inv_2 _31914_ (.A(_09873_),
    .Y(_09882_));
 sky130_fd_sc_hd__o21ai_2 _31915_ (.A1(_09874_),
    .A2(_09876_),
    .B1(_09882_),
    .Y(_09883_));
 sky130_fd_sc_hd__nand2_2 _31916_ (.A(_09881_),
    .B(_09883_),
    .Y(_09884_));
 sky130_fd_sc_hd__nand3_2 _31917_ (.A(_09872_),
    .B(_09868_),
    .C(_09884_),
    .Y(_09885_));
 sky130_fd_sc_hd__inv_2 _31918_ (.A(_09597_),
    .Y(_09886_));
 sky130_fd_sc_hd__a21o_2 _31919_ (.A1(_09879_),
    .A2(_09885_),
    .B1(_09886_),
    .X(_09887_));
 sky130_fd_sc_hd__nand3_2 _31920_ (.A(_09879_),
    .B(_09886_),
    .C(_09885_),
    .Y(_09888_));
 sky130_fd_sc_hd__nand2_2 _31921_ (.A(_09639_),
    .B(_09629_),
    .Y(_09889_));
 sky130_fd_sc_hd__nand2_2 _31922_ (.A(_09889_),
    .B(_09625_),
    .Y(_09890_));
 sky130_fd_sc_hd__nand3_2 _31923_ (.A(_09887_),
    .B(_09888_),
    .C(_09890_),
    .Y(_09891_));
 sky130_fd_sc_hd__inv_2 _31924_ (.A(_09629_),
    .Y(_09892_));
 sky130_fd_sc_hd__and3_2 _31925_ (.A(_09625_),
    .B(_09636_),
    .C(_09638_),
    .X(_09893_));
 sky130_fd_sc_hd__a21oi_2 _31926_ (.A1(_09879_),
    .A2(_09885_),
    .B1(_09886_),
    .Y(_09894_));
 sky130_fd_sc_hd__and3_2 _31927_ (.A(_09879_),
    .B(_09886_),
    .C(_09885_),
    .X(_09895_));
 sky130_fd_sc_hd__o22ai_2 _31928_ (.A1(_09892_),
    .A2(_09893_),
    .B1(_09894_),
    .B2(_09895_),
    .Y(_09896_));
 sky130_fd_sc_hd__nand3_2 _31929_ (.A(_09858_),
    .B(_09891_),
    .C(_09896_),
    .Y(_09897_));
 sky130_fd_sc_hd__nand2_2 _31930_ (.A(_09896_),
    .B(_09891_),
    .Y(_09898_));
 sky130_fd_sc_hd__nand3_2 _31931_ (.A(_09898_),
    .B(_09849_),
    .C(_09857_),
    .Y(_09899_));
 sky130_fd_sc_hd__nand3_2 _31932_ (.A(_09818_),
    .B(_09897_),
    .C(_09899_),
    .Y(_09900_));
 sky130_fd_sc_hd__inv_2 _31933_ (.A(_09613_),
    .Y(_09901_));
 sky130_fd_sc_hd__nand2_2 _31934_ (.A(_09658_),
    .B(_09901_),
    .Y(_09902_));
 sky130_fd_sc_hd__nand2_2 _31935_ (.A(_09858_),
    .B(_09898_),
    .Y(_09903_));
 sky130_fd_sc_hd__nand2_2 _31936_ (.A(_09852_),
    .B(_09856_),
    .Y(_09904_));
 sky130_fd_sc_hd__o2111ai_2 _31937_ (.A1(_09848_),
    .A2(_09904_),
    .B1(_09849_),
    .C1(_09891_),
    .D1(_09896_),
    .Y(_09905_));
 sky130_fd_sc_hd__nand3_2 _31938_ (.A(_09902_),
    .B(_09903_),
    .C(_09905_),
    .Y(_09906_));
 sky130_fd_sc_hd__nand2_2 _31939_ (.A(_09900_),
    .B(_09906_),
    .Y(_09907_));
 sky130_fd_sc_hd__a21oi_2 _31940_ (.A1(_09635_),
    .A2(_09637_),
    .B1(_09632_),
    .Y(_09908_));
 sky130_fd_sc_hd__nand2_2 _31941_ (.A(_07236_),
    .B(_05896_),
    .Y(_09909_));
 sky130_fd_sc_hd__nand2_2 _31942_ (.A(_06827_),
    .B(_19599_),
    .Y(_09910_));
 sky130_fd_sc_hd__nor2_2 _31943_ (.A(_09909_),
    .B(_09910_),
    .Y(_09911_));
 sky130_fd_sc_hd__buf_1 _31944_ (.A(_09911_),
    .X(_09912_));
 sky130_fd_sc_hd__and2_2 _31945_ (.A(_09909_),
    .B(_09910_),
    .X(_09913_));
 sky130_fd_sc_hd__nand2_2 _31946_ (.A(_19359_),
    .B(_08761_),
    .Y(_09914_));
 sky130_fd_sc_hd__o21ai_2 _31947_ (.A1(_09912_),
    .A2(_09913_),
    .B1(_09914_),
    .Y(_09915_));
 sky130_fd_sc_hd__inv_2 _31948_ (.A(_09914_),
    .Y(_09916_));
 sky130_fd_sc_hd__nand2_2 _31949_ (.A(_09909_),
    .B(_09910_),
    .Y(_09917_));
 sky130_fd_sc_hd__nand3b_2 _31950_ (.A_N(_09912_),
    .B(_09916_),
    .C(_09917_),
    .Y(_09918_));
 sky130_fd_sc_hd__nand3b_2 _31951_ (.A_N(_09908_),
    .B(_09915_),
    .C(_09918_),
    .Y(_09919_));
 sky130_fd_sc_hd__o21ai_2 _31952_ (.A1(_09912_),
    .A2(_09913_),
    .B1(_09916_),
    .Y(_09920_));
 sky130_fd_sc_hd__nand3b_2 _31953_ (.A_N(_09911_),
    .B(_09914_),
    .C(_09917_),
    .Y(_09921_));
 sky130_fd_sc_hd__nand3_2 _31954_ (.A(_09920_),
    .B(_09921_),
    .C(_09908_),
    .Y(_09922_));
 sky130_fd_sc_hd__a21oi_2 _31955_ (.A1(_09523_),
    .A2(_09522_),
    .B1(_09526_),
    .Y(_09923_));
 sky130_fd_sc_hd__inv_2 _31956_ (.A(_09923_),
    .Y(_09924_));
 sky130_fd_sc_hd__a21oi_2 _31957_ (.A1(_09919_),
    .A2(_09922_),
    .B1(_09924_),
    .Y(_09925_));
 sky130_fd_sc_hd__nand3_2 _31958_ (.A(_09919_),
    .B(_09922_),
    .C(_09924_),
    .Y(_09926_));
 sky130_fd_sc_hd__nand2_2 _31959_ (.A(_09528_),
    .B(_09534_),
    .Y(_09927_));
 sky130_fd_sc_hd__nand3_2 _31960_ (.A(_09926_),
    .B(_09532_),
    .C(_09927_),
    .Y(_09928_));
 sky130_fd_sc_hd__nor2_2 _31961_ (.A(_09925_),
    .B(_09928_),
    .Y(_09929_));
 sky130_fd_sc_hd__a21o_2 _31962_ (.A1(_09919_),
    .A2(_09922_),
    .B1(_09924_),
    .X(_09930_));
 sky130_fd_sc_hd__nand2_2 _31963_ (.A(_09536_),
    .B(_09528_),
    .Y(_09931_));
 sky130_fd_sc_hd__a21oi_2 _31964_ (.A1(_09930_),
    .A2(_09926_),
    .B1(_09931_),
    .Y(_09932_));
 sky130_fd_sc_hd__buf_1 _31965_ (.A(_07138_),
    .X(_09933_));
 sky130_fd_sc_hd__a22oi_2 _31966_ (.A1(_05807_),
    .A2(_08950_),
    .B1(_05808_),
    .B2(_09933_),
    .Y(_09934_));
 sky130_fd_sc_hd__nand2_2 _31967_ (.A(_09051_),
    .B(_19585_),
    .Y(_09935_));
 sky130_fd_sc_hd__nand2_2 _31968_ (.A(_06433_),
    .B(_09248_),
    .Y(_09936_));
 sky130_fd_sc_hd__nor2_2 _31969_ (.A(_09935_),
    .B(_09936_),
    .Y(_09937_));
 sky130_fd_sc_hd__nand2_2 _31970_ (.A(_19376_),
    .B(_08650_),
    .Y(_09938_));
 sky130_fd_sc_hd__inv_2 _31971_ (.A(_09938_),
    .Y(_09939_));
 sky130_fd_sc_hd__o21ai_2 _31972_ (.A1(_09934_),
    .A2(_09937_),
    .B1(_09939_),
    .Y(_09940_));
 sky130_fd_sc_hd__nor2_2 _31973_ (.A(_09934_),
    .B(_09937_),
    .Y(_09941_));
 sky130_fd_sc_hd__nand2_2 _31974_ (.A(_09941_),
    .B(_09938_),
    .Y(_09942_));
 sky130_fd_sc_hd__a21oi_2 _31975_ (.A1(_09546_),
    .A2(_09549_),
    .B1(_09543_),
    .Y(_09943_));
 sky130_fd_sc_hd__nand2_2 _31976_ (.A(_19363_),
    .B(_06560_),
    .Y(_09944_));
 sky130_fd_sc_hd__nand2_2 _31977_ (.A(_07450_),
    .B(_06946_),
    .Y(_09945_));
 sky130_fd_sc_hd__nor2_2 _31978_ (.A(_09944_),
    .B(_09945_),
    .Y(_09946_));
 sky130_fd_sc_hd__and2_2 _31979_ (.A(_09944_),
    .B(_09945_),
    .X(_09947_));
 sky130_fd_sc_hd__nand2_2 _31980_ (.A(_06446_),
    .B(_06728_),
    .Y(_09948_));
 sky130_fd_sc_hd__o21ai_2 _31981_ (.A1(_09946_),
    .A2(_09947_),
    .B1(_09948_),
    .Y(_09949_));
 sky130_fd_sc_hd__or2_2 _31982_ (.A(_09944_),
    .B(_09945_),
    .X(_09950_));
 sky130_fd_sc_hd__nand2_2 _31983_ (.A(_09944_),
    .B(_09945_),
    .Y(_09951_));
 sky130_fd_sc_hd__inv_2 _31984_ (.A(_09948_),
    .Y(_09952_));
 sky130_fd_sc_hd__nand3_2 _31985_ (.A(_09950_),
    .B(_09951_),
    .C(_09952_),
    .Y(_09953_));
 sky130_fd_sc_hd__nand3b_2 _31986_ (.A_N(_09943_),
    .B(_09949_),
    .C(_09953_),
    .Y(_09954_));
 sky130_fd_sc_hd__o21ai_2 _31987_ (.A1(_09946_),
    .A2(_09947_),
    .B1(_09952_),
    .Y(_09955_));
 sky130_fd_sc_hd__nand3_2 _31988_ (.A(_09950_),
    .B(_09951_),
    .C(_09948_),
    .Y(_09956_));
 sky130_fd_sc_hd__nand3_2 _31989_ (.A(_09955_),
    .B(_09956_),
    .C(_09943_),
    .Y(_09957_));
 sky130_fd_sc_hd__a22o_2 _31990_ (.A1(_09940_),
    .A2(_09942_),
    .B1(_09954_),
    .B2(_09957_),
    .X(_09958_));
 sky130_fd_sc_hd__nand2_2 _31991_ (.A(_09942_),
    .B(_09940_),
    .Y(_09959_));
 sky130_fd_sc_hd__nand3b_2 _31992_ (.A_N(_09959_),
    .B(_09957_),
    .C(_09954_),
    .Y(_09960_));
 sky130_fd_sc_hd__and2_2 _31993_ (.A(_09958_),
    .B(_09960_),
    .X(_09961_));
 sky130_fd_sc_hd__o21ai_2 _31994_ (.A1(_09929_),
    .A2(_09932_),
    .B1(_09961_),
    .Y(_09962_));
 sky130_fd_sc_hd__a21o_2 _31995_ (.A1(_09930_),
    .A2(_09926_),
    .B1(_09931_),
    .X(_09963_));
 sky130_fd_sc_hd__nand3_2 _31996_ (.A(_09930_),
    .B(_09931_),
    .C(_09926_),
    .Y(_09964_));
 sky130_fd_sc_hd__nand2_2 _31997_ (.A(_09958_),
    .B(_09960_),
    .Y(_09965_));
 sky130_fd_sc_hd__nand3_2 _31998_ (.A(_09963_),
    .B(_09964_),
    .C(_09965_),
    .Y(_09966_));
 sky130_fd_sc_hd__o21ai_2 _31999_ (.A1(_09648_),
    .A2(_09650_),
    .B1(_09646_),
    .Y(_09967_));
 sky130_fd_sc_hd__nand3_2 _32000_ (.A(_09962_),
    .B(_09966_),
    .C(_09967_),
    .Y(_09968_));
 sky130_fd_sc_hd__o21ai_2 _32001_ (.A1(_09929_),
    .A2(_09932_),
    .B1(_09965_),
    .Y(_09969_));
 sky130_fd_sc_hd__nand3_2 _32002_ (.A(_09963_),
    .B(_09961_),
    .C(_09964_),
    .Y(_09970_));
 sky130_fd_sc_hd__a21oi_2 _32003_ (.A1(_09642_),
    .A2(_09647_),
    .B1(_09651_),
    .Y(_09971_));
 sky130_fd_sc_hd__nand3_2 _32004_ (.A(_09969_),
    .B(_09970_),
    .C(_09971_),
    .Y(_09972_));
 sky130_fd_sc_hd__nor2_2 _32005_ (.A(_09540_),
    .B(_09572_),
    .Y(_09973_));
 sky130_fd_sc_hd__o2bb2ai_2 _32006_ (.A1_N(_09968_),
    .A2_N(_09972_),
    .B1(_09538_),
    .B2(_09973_),
    .Y(_09974_));
 sky130_fd_sc_hd__nor2_2 _32007_ (.A(_09538_),
    .B(_09973_),
    .Y(_09975_));
 sky130_fd_sc_hd__nand3_2 _32008_ (.A(_09972_),
    .B(_09968_),
    .C(_09975_),
    .Y(_09976_));
 sky130_fd_sc_hd__nand2_2 _32009_ (.A(_09974_),
    .B(_09976_),
    .Y(_09977_));
 sky130_fd_sc_hd__nand2_2 _32010_ (.A(_09907_),
    .B(_09977_),
    .Y(_09978_));
 sky130_fd_sc_hd__and3_2 _32011_ (.A(_09962_),
    .B(_09966_),
    .C(_09967_),
    .X(_09979_));
 sky130_fd_sc_hd__nand2_2 _32012_ (.A(_09972_),
    .B(_09975_),
    .Y(_09980_));
 sky130_fd_sc_hd__o2111ai_2 _32013_ (.A1(_09979_),
    .A2(_09980_),
    .B1(_09974_),
    .C1(_09906_),
    .D1(_09900_),
    .Y(_09981_));
 sky130_fd_sc_hd__nand3_2 _32014_ (.A(_09817_),
    .B(_09978_),
    .C(_09981_),
    .Y(_09982_));
 sky130_fd_sc_hd__a21oi_2 _32015_ (.A1(_09572_),
    .A2(_09573_),
    .B1(_09540_),
    .Y(_09983_));
 sky130_fd_sc_hd__a31oi_2 _32016_ (.A1(_09969_),
    .A2(_09970_),
    .A3(_09971_),
    .B1(_09983_),
    .Y(_09984_));
 sky130_fd_sc_hd__a2bb2oi_2 _32017_ (.A1_N(_09538_),
    .A2_N(_09973_),
    .B1(_09968_),
    .B2(_09972_),
    .Y(_09985_));
 sky130_fd_sc_hd__a21oi_2 _32018_ (.A1(_09968_),
    .A2(_09984_),
    .B1(_09985_),
    .Y(_09986_));
 sky130_fd_sc_hd__nand2_2 _32019_ (.A(_09986_),
    .B(_09907_),
    .Y(_09987_));
 sky130_fd_sc_hd__a31oi_2 _32020_ (.A1(_09660_),
    .A2(_09666_),
    .A3(_09665_),
    .B1(_09816_),
    .Y(_09988_));
 sky130_fd_sc_hd__nand3_2 _32021_ (.A(_09977_),
    .B(_09900_),
    .C(_09906_),
    .Y(_09989_));
 sky130_fd_sc_hd__nand3_2 _32022_ (.A(_09987_),
    .B(_09988_),
    .C(_09989_),
    .Y(_09990_));
 sky130_fd_sc_hd__and4_2 _32023_ (.A(_19380_),
    .B(_09247_),
    .C(_08497_),
    .D(_09250_),
    .X(_09991_));
 sky130_fd_sc_hd__nand2_2 _32024_ (.A(_05764_),
    .B(_09199_),
    .Y(_09992_));
 sky130_fd_sc_hd__inv_2 _32025_ (.A(_09992_),
    .Y(_09993_));
 sky130_fd_sc_hd__buf_1 _32026_ (.A(_19573_),
    .X(_09994_));
 sky130_fd_sc_hd__a22o_2 _32027_ (.A1(_08948_),
    .A2(_19578_),
    .B1(_09254_),
    .B2(_09994_),
    .X(_09995_));
 sky130_fd_sc_hd__nand3b_2 _32028_ (.A_N(_09991_),
    .B(_09993_),
    .C(_09995_),
    .Y(_09996_));
 sky130_fd_sc_hd__a21o_2 _32029_ (.A1(_09561_),
    .A2(_09558_),
    .B1(_09557_),
    .X(_09997_));
 sky130_fd_sc_hd__a22oi_2 _32030_ (.A1(_07797_),
    .A2(_08651_),
    .B1(_08949_),
    .B2(_19574_),
    .Y(_09998_));
 sky130_fd_sc_hd__o21ai_2 _32031_ (.A1(_09998_),
    .A2(_09991_),
    .B1(_09992_),
    .Y(_09999_));
 sky130_fd_sc_hd__nand3_2 _32032_ (.A(_09996_),
    .B(_09997_),
    .C(_09999_),
    .Y(_10000_));
 sky130_fd_sc_hd__nand3b_2 _32033_ (.A_N(_09991_),
    .B(_09992_),
    .C(_09995_),
    .Y(_10001_));
 sky130_fd_sc_hd__a21oi_2 _32034_ (.A1(_09561_),
    .A2(_09558_),
    .B1(_09557_),
    .Y(_10002_));
 sky130_fd_sc_hd__o21ai_2 _32035_ (.A1(_09998_),
    .A2(_09991_),
    .B1(_09993_),
    .Y(_10003_));
 sky130_fd_sc_hd__nand3_2 _32036_ (.A(_10001_),
    .B(_10002_),
    .C(_10003_),
    .Y(_10004_));
 sky130_fd_sc_hd__nand2_2 _32037_ (.A(_10000_),
    .B(_10004_),
    .Y(_10005_));
 sky130_fd_sc_hd__nor2_2 _32038_ (.A(_09686_),
    .B(_09683_),
    .Y(_10006_));
 sky130_fd_sc_hd__nand2_2 _32039_ (.A(_10005_),
    .B(_10006_),
    .Y(_10007_));
 sky130_fd_sc_hd__inv_2 _32040_ (.A(_10006_),
    .Y(_10008_));
 sky130_fd_sc_hd__nand3_2 _32041_ (.A(_10008_),
    .B(_10004_),
    .C(_10000_),
    .Y(_10009_));
 sky130_fd_sc_hd__o21a_2 _32042_ (.A1(_09543_),
    .A2(_09544_),
    .B1(_09545_),
    .X(_10010_));
 sky130_fd_sc_hd__a31o_2 _32043_ (.A1(_09549_),
    .A2(_09546_),
    .A3(_09548_),
    .B1(_09551_),
    .X(_10011_));
 sky130_fd_sc_hd__o2bb2ai_2 _32044_ (.A1_N(_09553_),
    .A2_N(_09564_),
    .B1(_10010_),
    .B2(_10011_),
    .Y(_10012_));
 sky130_fd_sc_hd__a21oi_2 _32045_ (.A1(_10007_),
    .A2(_10009_),
    .B1(_10012_),
    .Y(_10013_));
 sky130_fd_sc_hd__inv_2 _32046_ (.A(_10000_),
    .Y(_10014_));
 sky130_fd_sc_hd__nand2_2 _32047_ (.A(_10008_),
    .B(_10004_),
    .Y(_10015_));
 sky130_fd_sc_hd__o211a_2 _32048_ (.A1(_10014_),
    .A2(_10015_),
    .B1(_10007_),
    .C1(_10012_),
    .X(_10016_));
 sky130_fd_sc_hd__and2_2 _32049_ (.A(_09693_),
    .B(_09694_),
    .X(_10017_));
 sky130_fd_sc_hd__nor2_2 _32050_ (.A(_09700_),
    .B(_10017_),
    .Y(_10018_));
 sky130_fd_sc_hd__o21ai_2 _32051_ (.A1(_10013_),
    .A2(_10016_),
    .B1(_10018_),
    .Y(_10019_));
 sky130_fd_sc_hd__a21o_2 _32052_ (.A1(_10007_),
    .A2(_10009_),
    .B1(_10012_),
    .X(_10020_));
 sky130_fd_sc_hd__nand3_2 _32053_ (.A(_10012_),
    .B(_10007_),
    .C(_10009_),
    .Y(_10021_));
 sky130_fd_sc_hd__nand3b_2 _32054_ (.A_N(_10018_),
    .B(_10020_),
    .C(_10021_),
    .Y(_10022_));
 sky130_fd_sc_hd__o21ai_2 _32055_ (.A1(_09707_),
    .A2(_09699_),
    .B1(_09708_),
    .Y(_10023_));
 sky130_fd_sc_hd__nand3_2 _32056_ (.A(_10019_),
    .B(_10022_),
    .C(_10023_),
    .Y(_10024_));
 sky130_fd_sc_hd__o22ai_2 _32057_ (.A1(_09700_),
    .A2(_10017_),
    .B1(_10013_),
    .B2(_10016_),
    .Y(_10025_));
 sky130_fd_sc_hd__nand2_2 _32058_ (.A(_09708_),
    .B(_09707_),
    .Y(_10026_));
 sky130_fd_sc_hd__nand2_2 _32059_ (.A(_10026_),
    .B(_09706_),
    .Y(_10027_));
 sky130_fd_sc_hd__nand3_2 _32060_ (.A(_10020_),
    .B(_10021_),
    .C(_10018_),
    .Y(_10028_));
 sky130_fd_sc_hd__nand3_2 _32061_ (.A(_10025_),
    .B(_10027_),
    .C(_10028_),
    .Y(_10029_));
 sky130_fd_sc_hd__nand2_2 _32062_ (.A(_10024_),
    .B(_10029_),
    .Y(_10030_));
 sky130_fd_sc_hd__nand2_2 _32063_ (.A(_09742_),
    .B(_09732_),
    .Y(_10031_));
 sky130_fd_sc_hd__nand2_2 _32064_ (.A(_10031_),
    .B(_09729_),
    .Y(_10032_));
 sky130_fd_sc_hd__nand2_2 _32065_ (.A(_06051_),
    .B(_08664_),
    .Y(_10033_));
 sky130_fd_sc_hd__nand2_2 _32066_ (.A(_06054_),
    .B(_08920_),
    .Y(_10034_));
 sky130_fd_sc_hd__nor2_2 _32067_ (.A(_10033_),
    .B(_10034_),
    .Y(_10035_));
 sky130_fd_sc_hd__and2_2 _32068_ (.A(_10033_),
    .B(_10034_),
    .X(_10036_));
 sky130_fd_sc_hd__nand2_2 _32069_ (.A(_19404_),
    .B(_19549_),
    .Y(_10037_));
 sky130_fd_sc_hd__o21ai_2 _32070_ (.A1(_10035_),
    .A2(_10036_),
    .B1(_10037_),
    .Y(_10038_));
 sky130_fd_sc_hd__or2_2 _32071_ (.A(_10033_),
    .B(_10034_),
    .X(_10039_));
 sky130_fd_sc_hd__inv_2 _32072_ (.A(_10037_),
    .Y(_10040_));
 sky130_fd_sc_hd__nand2_2 _32073_ (.A(_10033_),
    .B(_10034_),
    .Y(_10041_));
 sky130_fd_sc_hd__nand3_2 _32074_ (.A(_10039_),
    .B(_10040_),
    .C(_10041_),
    .Y(_10042_));
 sky130_fd_sc_hd__a21o_2 _32075_ (.A1(_09726_),
    .A2(_09727_),
    .B1(_09720_),
    .X(_10043_));
 sky130_fd_sc_hd__nand3_2 _32076_ (.A(_10038_),
    .B(_10042_),
    .C(_10043_),
    .Y(_10044_));
 sky130_fd_sc_hd__o21ai_2 _32077_ (.A1(_10035_),
    .A2(_10036_),
    .B1(_10040_),
    .Y(_10045_));
 sky130_fd_sc_hd__nand3_2 _32078_ (.A(_10039_),
    .B(_10037_),
    .C(_10041_),
    .Y(_10046_));
 sky130_fd_sc_hd__a21oi_2 _32079_ (.A1(_09726_),
    .A2(_09727_),
    .B1(_09720_),
    .Y(_10047_));
 sky130_fd_sc_hd__nand3_2 _32080_ (.A(_10045_),
    .B(_10046_),
    .C(_10047_),
    .Y(_10048_));
 sky130_fd_sc_hd__nand2_2 _32081_ (.A(_10044_),
    .B(_10048_),
    .Y(_10049_));
 sky130_fd_sc_hd__buf_1 _32082_ (.A(_19552_),
    .X(_10050_));
 sky130_fd_sc_hd__nand2_2 _32083_ (.A(_06072_),
    .B(_19558_),
    .Y(_10051_));
 sky130_fd_sc_hd__a21o_2 _32084_ (.A1(_05144_),
    .A2(_10050_),
    .B1(_10051_),
    .X(_10052_));
 sky130_fd_sc_hd__nand2_2 _32085_ (.A(_06220_),
    .B(_19553_),
    .Y(_10053_));
 sky130_fd_sc_hd__a21o_2 _32086_ (.A1(_05141_),
    .A2(_09733_),
    .B1(_10053_),
    .X(_10054_));
 sky130_fd_sc_hd__buf_1 _32087_ (.A(_09220_),
    .X(_10055_));
 sky130_fd_sc_hd__nand2_2 _32088_ (.A(_05116_),
    .B(_10055_),
    .Y(_10056_));
 sky130_fd_sc_hd__a21o_2 _32089_ (.A1(_10052_),
    .A2(_10054_),
    .B1(_10056_),
    .X(_10057_));
 sky130_fd_sc_hd__nand3_2 _32090_ (.A(_10052_),
    .B(_10054_),
    .C(_10056_),
    .Y(_10058_));
 sky130_fd_sc_hd__nand2_2 _32091_ (.A(_10057_),
    .B(_10058_),
    .Y(_10059_));
 sky130_fd_sc_hd__nand2_2 _32092_ (.A(_10049_),
    .B(_10059_),
    .Y(_10060_));
 sky130_fd_sc_hd__and2_2 _32093_ (.A(_10057_),
    .B(_10058_),
    .X(_10061_));
 sky130_fd_sc_hd__nand3_2 _32094_ (.A(_10061_),
    .B(_10044_),
    .C(_10048_),
    .Y(_10062_));
 sky130_fd_sc_hd__nand3_2 _32095_ (.A(_10032_),
    .B(_10060_),
    .C(_10062_),
    .Y(_10063_));
 sky130_fd_sc_hd__inv_2 _32096_ (.A(_09740_),
    .Y(_10064_));
 sky130_fd_sc_hd__or2_2 _32097_ (.A(_09734_),
    .B(_09737_),
    .X(_10065_));
 sky130_fd_sc_hd__nand2_2 _32098_ (.A(_10064_),
    .B(_10065_),
    .Y(_10066_));
 sky130_fd_sc_hd__nand2_2 _32099_ (.A(_10063_),
    .B(_10066_),
    .Y(_10067_));
 sky130_fd_sc_hd__inv_2 _32100_ (.A(_09732_),
    .Y(_10068_));
 sky130_fd_sc_hd__o21a_2 _32101_ (.A1(_09740_),
    .A2(_09741_),
    .B1(_09729_),
    .X(_10069_));
 sky130_fd_sc_hd__o2bb2ai_2 _32102_ (.A1_N(_10062_),
    .A2_N(_10060_),
    .B1(_10068_),
    .B2(_10069_),
    .Y(_10070_));
 sky130_fd_sc_hd__inv_2 _32103_ (.A(_10070_),
    .Y(_10071_));
 sky130_fd_sc_hd__a21o_2 _32104_ (.A1(_10070_),
    .A2(_10063_),
    .B1(_10066_),
    .X(_10072_));
 sky130_fd_sc_hd__o21ai_2 _32105_ (.A1(_10067_),
    .A2(_10071_),
    .B1(_10072_),
    .Y(_10073_));
 sky130_fd_sc_hd__nand2_2 _32106_ (.A(_10030_),
    .B(_10073_),
    .Y(_10074_));
 sky130_fd_sc_hd__a21oi_2 _32107_ (.A1(_10070_),
    .A2(_10063_),
    .B1(_10066_),
    .Y(_10075_));
 sky130_fd_sc_hd__and3_2 _32108_ (.A(_10070_),
    .B(_10066_),
    .C(_10063_),
    .X(_10076_));
 sky130_fd_sc_hd__nor2_2 _32109_ (.A(_10075_),
    .B(_10076_),
    .Y(_10077_));
 sky130_fd_sc_hd__nand3_2 _32110_ (.A(_10077_),
    .B(_10024_),
    .C(_10029_),
    .Y(_10078_));
 sky130_fd_sc_hd__nand2_2 _32111_ (.A(_09673_),
    .B(_09577_),
    .Y(_10079_));
 sky130_fd_sc_hd__nand3_2 _32112_ (.A(_10074_),
    .B(_10078_),
    .C(_10079_),
    .Y(_10080_));
 sky130_fd_sc_hd__nand2_2 _32113_ (.A(_10030_),
    .B(_10077_),
    .Y(_10081_));
 sky130_fd_sc_hd__a21boi_2 _32114_ (.A1(_09581_),
    .A2(_09583_),
    .B1_N(_09577_),
    .Y(_10082_));
 sky130_fd_sc_hd__nand3_2 _32115_ (.A(_10073_),
    .B(_10024_),
    .C(_10029_),
    .Y(_10083_));
 sky130_fd_sc_hd__nand3_2 _32116_ (.A(_10081_),
    .B(_10082_),
    .C(_10083_),
    .Y(_10084_));
 sky130_fd_sc_hd__and3_2 _32117_ (.A(_09711_),
    .B(_09712_),
    .C(_09713_),
    .X(_10085_));
 sky130_fd_sc_hd__a21o_2 _32118_ (.A1(_09755_),
    .A2(_09710_),
    .B1(_10085_),
    .X(_10086_));
 sky130_fd_sc_hd__a21oi_2 _32119_ (.A1(_10080_),
    .A2(_10084_),
    .B1(_10086_),
    .Y(_10087_));
 sky130_fd_sc_hd__a21oi_2 _32120_ (.A1(_10081_),
    .A2(_10083_),
    .B1(_10082_),
    .Y(_10088_));
 sky130_fd_sc_hd__nand2_2 _32121_ (.A(_10084_),
    .B(_10086_),
    .Y(_10089_));
 sky130_fd_sc_hd__nor2_2 _32122_ (.A(_10088_),
    .B(_10089_),
    .Y(_10090_));
 sky130_fd_sc_hd__o2bb2ai_2 _32123_ (.A1_N(_09982_),
    .A2_N(_09990_),
    .B1(_10087_),
    .B2(_10090_),
    .Y(_10091_));
 sky130_fd_sc_hd__nand2_2 _32124_ (.A(_10080_),
    .B(_10084_),
    .Y(_10092_));
 sky130_fd_sc_hd__a21oi_2 _32125_ (.A1(_09755_),
    .A2(_09710_),
    .B1(_10085_),
    .Y(_10093_));
 sky130_fd_sc_hd__nand2_2 _32126_ (.A(_10092_),
    .B(_10093_),
    .Y(_10094_));
 sky130_fd_sc_hd__o2111ai_2 _32127_ (.A1(_10088_),
    .A2(_10089_),
    .B1(_10094_),
    .C1(_09990_),
    .D1(_09982_),
    .Y(_10095_));
 sky130_fd_sc_hd__nand3_2 _32128_ (.A(_09815_),
    .B(_10091_),
    .C(_10095_),
    .Y(_10096_));
 sky130_fd_sc_hd__and3_2 _32129_ (.A(_09670_),
    .B(_09671_),
    .C(_09674_),
    .X(_10097_));
 sky130_fd_sc_hd__a31oi_2 _32130_ (.A1(_09770_),
    .A2(_09668_),
    .A3(_09772_),
    .B1(_10097_),
    .Y(_10098_));
 sky130_fd_sc_hd__nand2_2 _32131_ (.A(_09982_),
    .B(_09990_),
    .Y(_10099_));
 sky130_fd_sc_hd__a31oi_2 _32132_ (.A1(_10081_),
    .A2(_10082_),
    .A3(_10083_),
    .B1(_10093_),
    .Y(_10100_));
 sky130_fd_sc_hd__a21oi_2 _32133_ (.A1(_10080_),
    .A2(_10100_),
    .B1(_10087_),
    .Y(_10101_));
 sky130_fd_sc_hd__nand2_2 _32134_ (.A(_10099_),
    .B(_10101_),
    .Y(_10102_));
 sky130_fd_sc_hd__o211ai_2 _32135_ (.A1(_10087_),
    .A2(_10090_),
    .B1(_09982_),
    .C1(_09990_),
    .Y(_10103_));
 sky130_fd_sc_hd__nand3_2 _32136_ (.A(_10098_),
    .B(_10102_),
    .C(_10103_),
    .Y(_10104_));
 sky130_fd_sc_hd__nand2_2 _32137_ (.A(_09745_),
    .B(_09752_),
    .Y(_10105_));
 sky130_fd_sc_hd__and2_2 _32138_ (.A(_10105_),
    .B(_09748_),
    .X(_10106_));
 sky130_fd_sc_hd__a21o_2 _32139_ (.A1(_09776_),
    .A2(_09766_),
    .B1(_10106_),
    .X(_10107_));
 sky130_fd_sc_hd__inv_2 _32140_ (.A(_10107_),
    .Y(_10108_));
 sky130_fd_sc_hd__nand3_2 _32141_ (.A(_09776_),
    .B(_09766_),
    .C(_10106_),
    .Y(_10109_));
 sky130_fd_sc_hd__inv_2 _32142_ (.A(_10109_),
    .Y(_10110_));
 sky130_fd_sc_hd__o2bb2ai_2 _32143_ (.A1_N(_10096_),
    .A2_N(_10104_),
    .B1(_10108_),
    .B2(_10110_),
    .Y(_10111_));
 sky130_fd_sc_hd__and2_2 _32144_ (.A(_10107_),
    .B(_10109_),
    .X(_10112_));
 sky130_fd_sc_hd__nand3_2 _32145_ (.A(_10104_),
    .B(_10096_),
    .C(_10112_),
    .Y(_10113_));
 sky130_fd_sc_hd__o21ai_2 _32146_ (.A1(_09799_),
    .A2(_09780_),
    .B1(_09790_),
    .Y(_10114_));
 sky130_fd_sc_hd__a21oi_2 _32147_ (.A1(_10111_),
    .A2(_10113_),
    .B1(_10114_),
    .Y(_10115_));
 sky130_fd_sc_hd__and3_2 _32148_ (.A(_09815_),
    .B(_10091_),
    .C(_10095_),
    .X(_10116_));
 sky130_fd_sc_hd__nand2_2 _32149_ (.A(_10104_),
    .B(_10112_),
    .Y(_10117_));
 sky130_fd_sc_hd__o211a_2 _32150_ (.A1(_10116_),
    .A2(_10117_),
    .B1(_10111_),
    .C1(_10114_),
    .X(_10118_));
 sky130_fd_sc_hd__o21ai_2 _32151_ (.A1(_10115_),
    .A2(_10118_),
    .B1(_09517_),
    .Y(_10119_));
 sky130_fd_sc_hd__a21boi_2 _32152_ (.A1(_09801_),
    .A2(_09483_),
    .B1_N(_09796_),
    .Y(_10120_));
 sky130_fd_sc_hd__a21o_2 _32153_ (.A1(_10111_),
    .A2(_10113_),
    .B1(_10114_),
    .X(_10121_));
 sky130_fd_sc_hd__nand3_2 _32154_ (.A(_10114_),
    .B(_10111_),
    .C(_10113_),
    .Y(_10122_));
 sky130_fd_sc_hd__nand3_2 _32155_ (.A(_10121_),
    .B(_09516_),
    .C(_10122_),
    .Y(_10123_));
 sky130_fd_sc_hd__nand3_2 _32156_ (.A(_10119_),
    .B(_10120_),
    .C(_10123_),
    .Y(_10124_));
 sky130_fd_sc_hd__o21ai_2 _32157_ (.A1(_10115_),
    .A2(_10118_),
    .B1(_09516_),
    .Y(_10125_));
 sky130_fd_sc_hd__nand2_2 _32158_ (.A(_09786_),
    .B(_09795_),
    .Y(_10126_));
 sky130_fd_sc_hd__inv_2 _32159_ (.A(_09784_),
    .Y(_10127_));
 sky130_fd_sc_hd__o2bb2ai_2 _32160_ (.A1_N(_09483_),
    .A2_N(_09801_),
    .B1(_10126_),
    .B2(_10127_),
    .Y(_10128_));
 sky130_fd_sc_hd__nand3_2 _32161_ (.A(_10121_),
    .B(_09517_),
    .C(_10122_),
    .Y(_10129_));
 sky130_fd_sc_hd__nand3_2 _32162_ (.A(_10125_),
    .B(_10128_),
    .C(_10129_),
    .Y(_10130_));
 sky130_fd_sc_hd__nand2_2 _32163_ (.A(_10124_),
    .B(_10130_),
    .Y(_10131_));
 sky130_fd_sc_hd__nand2_2 _32164_ (.A(_09813_),
    .B(_09806_),
    .Y(_10132_));
 sky130_fd_sc_hd__nand2_2 _32165_ (.A(_10132_),
    .B(_09805_),
    .Y(_10133_));
 sky130_fd_sc_hd__xor2_2 _32166_ (.A(_10131_),
    .B(_10133_),
    .X(_02648_));
 sky130_fd_sc_hd__nand3_2 _32167_ (.A(_09849_),
    .B(_09896_),
    .C(_09891_),
    .Y(_10134_));
 sky130_fd_sc_hd__nand2_2 _32168_ (.A(_10134_),
    .B(_09857_),
    .Y(_10135_));
 sky130_fd_sc_hd__buf_1 _32169_ (.A(_19319_),
    .X(_10136_));
 sky130_fd_sc_hd__nand2_2 _32170_ (.A(_10136_),
    .B(_08393_),
    .Y(_10137_));
 sky130_fd_sc_hd__buf_1 _32171_ (.A(_09841_),
    .X(_10138_));
 sky130_fd_sc_hd__buf_1 _32172_ (.A(_10138_),
    .X(_10139_));
 sky130_fd_sc_hd__nand3b_2 _32173_ (.A_N(_10137_),
    .B(_10139_),
    .C(_19637_),
    .Y(_10140_));
 sky130_fd_sc_hd__buf_1 _32174_ (.A(\pcpi_mul.rs2[28] ),
    .X(_10141_));
 sky130_fd_sc_hd__a22o_2 _32175_ (.A1(_10138_),
    .A2(_07904_),
    .B1(_10141_),
    .B2(_05215_),
    .X(_10142_));
 sky130_fd_sc_hd__nand2_2 _32176_ (.A(_19322_),
    .B(_06792_),
    .Y(_10143_));
 sky130_fd_sc_hd__inv_2 _32177_ (.A(_10143_),
    .Y(_10144_));
 sky130_fd_sc_hd__nand3_2 _32178_ (.A(_10140_),
    .B(_10142_),
    .C(_10144_),
    .Y(_10145_));
 sky130_fd_sc_hd__buf_1 _32179_ (.A(_09841_),
    .X(_10146_));
 sky130_fd_sc_hd__a22oi_2 _32180_ (.A1(_10146_),
    .A2(_05124_),
    .B1(_19320_),
    .B2(_05120_),
    .Y(_10147_));
 sky130_fd_sc_hd__and4_2 _32181_ (.A(_19315_),
    .B(_09602_),
    .C(_05545_),
    .D(_07904_),
    .X(_10148_));
 sky130_fd_sc_hd__o21ai_2 _32182_ (.A1(_10147_),
    .A2(_10148_),
    .B1(_10143_),
    .Y(_10149_));
 sky130_fd_sc_hd__inv_2 _32183_ (.A(\pcpi_mul.rs2[30] ),
    .Y(_10150_));
 sky130_fd_sc_hd__buf_1 _32184_ (.A(_10150_),
    .X(_10151_));
 sky130_fd_sc_hd__buf_1 _32185_ (.A(_10151_),
    .X(_10152_));
 sky130_fd_sc_hd__o2bb2ai_2 _32186_ (.A1_N(_10145_),
    .A2_N(_10149_),
    .B1(_10152_),
    .B2(_04839_),
    .Y(_10153_));
 sky130_fd_sc_hd__nor2_2 _32187_ (.A(_10151_),
    .B(_04839_),
    .Y(_10154_));
 sky130_fd_sc_hd__nand3_2 _32188_ (.A(_10149_),
    .B(_10145_),
    .C(_10154_),
    .Y(_10155_));
 sky130_fd_sc_hd__buf_1 _32189_ (.A(_09120_),
    .X(_10156_));
 sky130_fd_sc_hd__a22oi_2 _32190_ (.A1(_19328_),
    .A2(_05207_),
    .B1(_10156_),
    .B2(_05341_),
    .Y(_10157_));
 sky130_fd_sc_hd__buf_1 _32191_ (.A(\pcpi_mul.rs2[25] ),
    .X(_10158_));
 sky130_fd_sc_hd__nand3_2 _32192_ (.A(_19327_),
    .B(_10158_),
    .C(_05222_),
    .Y(_10159_));
 sky130_fd_sc_hd__nor2_2 _32193_ (.A(_05856_),
    .B(_10159_),
    .Y(_10160_));
 sky130_fd_sc_hd__nand2_2 _32194_ (.A(_19333_),
    .B(_05347_),
    .Y(_10161_));
 sky130_fd_sc_hd__inv_2 _32195_ (.A(_10161_),
    .Y(_10162_));
 sky130_fd_sc_hd__o21ai_2 _32196_ (.A1(_10157_),
    .A2(_10160_),
    .B1(_10162_),
    .Y(_10163_));
 sky130_fd_sc_hd__nand2_2 _32197_ (.A(_09840_),
    .B(_09843_),
    .Y(_10164_));
 sky130_fd_sc_hd__a31oi_2 _32198_ (.A1(_10164_),
    .A2(_19324_),
    .A3(_19634_),
    .B1(_09844_),
    .Y(_10165_));
 sky130_fd_sc_hd__buf_1 _32199_ (.A(_09339_),
    .X(_10166_));
 sky130_fd_sc_hd__a22o_2 _32200_ (.A1(_10166_),
    .A2(_05207_),
    .B1(_10156_),
    .B2(_05341_),
    .X(_10167_));
 sky130_fd_sc_hd__o211ai_2 _32201_ (.A1(_05865_),
    .A2(_10159_),
    .B1(_10161_),
    .C1(_10167_),
    .Y(_10168_));
 sky130_fd_sc_hd__nand3_2 _32202_ (.A(_10163_),
    .B(_10165_),
    .C(_10168_),
    .Y(_10169_));
 sky130_fd_sc_hd__o21ai_2 _32203_ (.A1(_10157_),
    .A2(_10160_),
    .B1(_10161_),
    .Y(_10170_));
 sky130_fd_sc_hd__nand3b_2 _32204_ (.A_N(_09840_),
    .B(_10146_),
    .C(_06598_),
    .Y(_10171_));
 sky130_fd_sc_hd__o21ai_2 _32205_ (.A1(_09837_),
    .A2(_09839_),
    .B1(_10171_),
    .Y(_10172_));
 sky130_fd_sc_hd__o211ai_2 _32206_ (.A1(_05865_),
    .A2(_10159_),
    .B1(_10162_),
    .C1(_10167_),
    .Y(_10173_));
 sky130_fd_sc_hd__nand3_2 _32207_ (.A(_10170_),
    .B(_10172_),
    .C(_10173_),
    .Y(_10174_));
 sky130_fd_sc_hd__nand2_2 _32208_ (.A(_10169_),
    .B(_10174_),
    .Y(_10175_));
 sky130_fd_sc_hd__a21oi_2 _32209_ (.A1(_09828_),
    .A2(_09824_),
    .B1(_09822_),
    .Y(_10176_));
 sky130_fd_sc_hd__nand2_2 _32210_ (.A(_10175_),
    .B(_10176_),
    .Y(_10177_));
 sky130_fd_sc_hd__a21o_2 _32211_ (.A1(_09828_),
    .A2(_09824_),
    .B1(_09822_),
    .X(_10178_));
 sky130_fd_sc_hd__nand3_2 _32212_ (.A(_10169_),
    .B(_10174_),
    .C(_10178_),
    .Y(_10179_));
 sky130_fd_sc_hd__a22oi_2 _32213_ (.A1(_10153_),
    .A2(_10155_),
    .B1(_10177_),
    .B2(_10179_),
    .Y(_10180_));
 sky130_fd_sc_hd__nand2_2 _32214_ (.A(_10153_),
    .B(_10155_),
    .Y(_10181_));
 sky130_fd_sc_hd__a21oi_2 _32215_ (.A1(_10169_),
    .A2(_10174_),
    .B1(_10178_),
    .Y(_10182_));
 sky130_fd_sc_hd__nor3b_2 _32216_ (.A(_10181_),
    .B(_10182_),
    .C_N(_10179_),
    .Y(_10183_));
 sky130_fd_sc_hd__o22ai_2 _32217_ (.A1(_09851_),
    .A2(_09850_),
    .B1(_10180_),
    .B2(_10183_),
    .Y(_10184_));
 sky130_fd_sc_hd__nand2_2 _32218_ (.A(_10177_),
    .B(_10179_),
    .Y(_10185_));
 sky130_fd_sc_hd__nand2_2 _32219_ (.A(_10185_),
    .B(_10181_),
    .Y(_10186_));
 sky130_fd_sc_hd__nand3b_2 _32220_ (.A_N(_10181_),
    .B(_10177_),
    .C(_10179_),
    .Y(_10187_));
 sky130_fd_sc_hd__nand3_2 _32221_ (.A(_09848_),
    .B(_10186_),
    .C(_10187_),
    .Y(_10188_));
 sky130_fd_sc_hd__nand2_2 _32222_ (.A(_10184_),
    .B(_10188_),
    .Y(_10189_));
 sky130_fd_sc_hd__inv_2 _32223_ (.A(_09868_),
    .Y(_10190_));
 sky130_fd_sc_hd__and3_2 _32224_ (.A(_09872_),
    .B(_09883_),
    .C(_09881_),
    .X(_10191_));
 sky130_fd_sc_hd__a31o_2 _32225_ (.A1(_09831_),
    .A2(_09605_),
    .A3(_09832_),
    .B1(_09834_),
    .X(_10192_));
 sky130_fd_sc_hd__buf_1 _32226_ (.A(_08391_),
    .X(_10193_));
 sky130_fd_sc_hd__a22oi_2 _32227_ (.A1(_10193_),
    .A2(_05713_),
    .B1(_08799_),
    .B2(_05893_),
    .Y(_10194_));
 sky130_fd_sc_hd__nand3_2 _32228_ (.A(_08396_),
    .B(_07974_),
    .C(_05505_),
    .Y(_10195_));
 sky130_fd_sc_hd__nor2_2 _32229_ (.A(_05731_),
    .B(_10195_),
    .Y(_10196_));
 sky130_fd_sc_hd__nand2_2 _32230_ (.A(_07976_),
    .B(_07210_),
    .Y(_10197_));
 sky130_fd_sc_hd__o21ai_2 _32231_ (.A1(_10194_),
    .A2(_10196_),
    .B1(_10197_),
    .Y(_10198_));
 sky130_fd_sc_hd__o22ai_2 _32232_ (.A1(_06333_),
    .A2(_09860_),
    .B1(_09862_),
    .B2(_09859_),
    .Y(_10199_));
 sky130_fd_sc_hd__inv_2 _32233_ (.A(_10197_),
    .Y(_10200_));
 sky130_fd_sc_hd__a22o_2 _32234_ (.A1(_10193_),
    .A2(_05713_),
    .B1(_08799_),
    .B2(_05893_),
    .X(_10201_));
 sky130_fd_sc_hd__o211ai_2 _32235_ (.A1(_05732_),
    .A2(_10195_),
    .B1(_10200_),
    .C1(_10201_),
    .Y(_10202_));
 sky130_fd_sc_hd__nand3_2 _32236_ (.A(_10198_),
    .B(_10199_),
    .C(_10202_),
    .Y(_10203_));
 sky130_fd_sc_hd__o21ai_2 _32237_ (.A1(_10194_),
    .A2(_10196_),
    .B1(_10200_),
    .Y(_10204_));
 sky130_fd_sc_hd__a21oi_2 _32238_ (.A1(_09866_),
    .A2(_09863_),
    .B1(_09861_),
    .Y(_10205_));
 sky130_fd_sc_hd__o211ai_2 _32239_ (.A1(_05732_),
    .A2(_10195_),
    .B1(_10197_),
    .C1(_10201_),
    .Y(_10206_));
 sky130_fd_sc_hd__nand3_2 _32240_ (.A(_10204_),
    .B(_10205_),
    .C(_10206_),
    .Y(_10207_));
 sky130_fd_sc_hd__nand2_2 _32241_ (.A(_08808_),
    .B(_05738_),
    .Y(_10208_));
 sky130_fd_sc_hd__nand3b_2 _32242_ (.A_N(_10208_),
    .B(_08816_),
    .C(_19607_),
    .Y(_10209_));
 sky130_fd_sc_hd__buf_1 _32243_ (.A(_07722_),
    .X(_10210_));
 sky130_fd_sc_hd__a22o_2 _32244_ (.A1(_10210_),
    .A2(_19610_),
    .B1(_08816_),
    .B2(_06074_),
    .X(_10211_));
 sky130_fd_sc_hd__nand2_2 _32245_ (.A(_08407_),
    .B(_06726_),
    .Y(_10212_));
 sky130_fd_sc_hd__inv_2 _32246_ (.A(_10212_),
    .Y(_10213_));
 sky130_fd_sc_hd__and3_2 _32247_ (.A(_10209_),
    .B(_10211_),
    .C(_10213_),
    .X(_10214_));
 sky130_fd_sc_hd__a21oi_2 _32248_ (.A1(_10209_),
    .A2(_10211_),
    .B1(_10213_),
    .Y(_10215_));
 sky130_fd_sc_hd__o2bb2ai_2 _32249_ (.A1_N(_10203_),
    .A2_N(_10207_),
    .B1(_10214_),
    .B2(_10215_),
    .Y(_10216_));
 sky130_fd_sc_hd__a22oi_2 _32250_ (.A1(_10210_),
    .A2(_19610_),
    .B1(_08816_),
    .B2(_19607_),
    .Y(_10217_));
 sky130_fd_sc_hd__and4_2 _32251_ (.A(_10210_),
    .B(_08809_),
    .C(_06074_),
    .D(_09010_),
    .X(_10218_));
 sky130_fd_sc_hd__o21ai_2 _32252_ (.A1(_10217_),
    .A2(_10218_),
    .B1(_10213_),
    .Y(_10219_));
 sky130_fd_sc_hd__nand3_2 _32253_ (.A(_10209_),
    .B(_10211_),
    .C(_10212_),
    .Y(_10220_));
 sky130_fd_sc_hd__nand2_2 _32254_ (.A(_10219_),
    .B(_10220_),
    .Y(_10221_));
 sky130_fd_sc_hd__nand3_2 _32255_ (.A(_10207_),
    .B(_10203_),
    .C(_10221_),
    .Y(_10222_));
 sky130_fd_sc_hd__a22oi_2 _32256_ (.A1(_09830_),
    .A2(_10192_),
    .B1(_10216_),
    .B2(_10222_),
    .Y(_10223_));
 sky130_fd_sc_hd__a21oi_2 _32257_ (.A1(_10207_),
    .A2(_10203_),
    .B1(_10221_),
    .Y(_10224_));
 sky130_fd_sc_hd__nand3_2 _32258_ (.A(_10222_),
    .B(_10192_),
    .C(_09830_),
    .Y(_10225_));
 sky130_fd_sc_hd__nor2_2 _32259_ (.A(_10224_),
    .B(_10225_),
    .Y(_10226_));
 sky130_fd_sc_hd__o22ai_2 _32260_ (.A1(_10190_),
    .A2(_10191_),
    .B1(_10223_),
    .B2(_10226_),
    .Y(_10227_));
 sky130_fd_sc_hd__nand2_2 _32261_ (.A(_09836_),
    .B(_09833_),
    .Y(_10228_));
 sky130_fd_sc_hd__a21o_2 _32262_ (.A1(_10222_),
    .A2(_10216_),
    .B1(_10228_),
    .X(_10229_));
 sky130_fd_sc_hd__nand3_2 _32263_ (.A(_10228_),
    .B(_10222_),
    .C(_10216_),
    .Y(_10230_));
 sky130_fd_sc_hd__nand2_2 _32264_ (.A(_09868_),
    .B(_09884_),
    .Y(_10231_));
 sky130_fd_sc_hd__nand2_2 _32265_ (.A(_10231_),
    .B(_09872_),
    .Y(_10232_));
 sky130_fd_sc_hd__nand3_2 _32266_ (.A(_10229_),
    .B(_10230_),
    .C(_10232_),
    .Y(_10233_));
 sky130_fd_sc_hd__nand2_2 _32267_ (.A(_10227_),
    .B(_10233_),
    .Y(_10234_));
 sky130_fd_sc_hd__nand2_2 _32268_ (.A(_10189_),
    .B(_10234_),
    .Y(_10235_));
 sky130_fd_sc_hd__nand3_2 _32269_ (.A(_10187_),
    .B(_09836_),
    .C(_09854_),
    .Y(_10236_));
 sky130_fd_sc_hd__o2111ai_2 _32270_ (.A1(_10180_),
    .A2(_10236_),
    .B1(_10233_),
    .C1(_10227_),
    .D1(_10184_),
    .Y(_10237_));
 sky130_fd_sc_hd__nand3_2 _32271_ (.A(_10135_),
    .B(_10235_),
    .C(_10237_),
    .Y(_10238_));
 sky130_fd_sc_hd__nand3_2 _32272_ (.A(_10234_),
    .B(_10184_),
    .C(_10188_),
    .Y(_10239_));
 sky130_fd_sc_hd__nand3_2 _32273_ (.A(_10189_),
    .B(_10227_),
    .C(_10233_),
    .Y(_10240_));
 sky130_fd_sc_hd__o2111ai_2 _32274_ (.A1(_09848_),
    .A2(_09904_),
    .B1(_10134_),
    .C1(_10239_),
    .D1(_10240_),
    .Y(_10241_));
 sky130_fd_sc_hd__a22oi_2 _32275_ (.A1(_09008_),
    .A2(_06736_),
    .B1(_09009_),
    .B2(_06935_),
    .Y(_10242_));
 sky130_fd_sc_hd__nand3_2 _32276_ (.A(_07886_),
    .B(_08345_),
    .C(_19600_),
    .Y(_10243_));
 sky130_fd_sc_hd__nor2_2 _32277_ (.A(_06401_),
    .B(_10243_),
    .Y(_10244_));
 sky130_fd_sc_hd__nand2_2 _32278_ (.A(_19359_),
    .B(_06373_),
    .Y(_10245_));
 sky130_fd_sc_hd__inv_2 _32279_ (.A(_10245_),
    .Y(_10246_));
 sky130_fd_sc_hd__o21ai_2 _32280_ (.A1(_10242_),
    .A2(_10244_),
    .B1(_10246_),
    .Y(_10247_));
 sky130_fd_sc_hd__a21oi_2 _32281_ (.A1(_09880_),
    .A2(_09882_),
    .B1(_09876_),
    .Y(_10248_));
 sky130_fd_sc_hd__a22o_2 _32282_ (.A1(_09008_),
    .A2(_06736_),
    .B1(_09009_),
    .B2(_06935_),
    .X(_10249_));
 sky130_fd_sc_hd__o211ai_2 _32283_ (.A1(_06397_),
    .A2(_10243_),
    .B1(_10245_),
    .C1(_10249_),
    .Y(_10250_));
 sky130_fd_sc_hd__nand3_2 _32284_ (.A(_10247_),
    .B(_10248_),
    .C(_10250_),
    .Y(_10251_));
 sky130_fd_sc_hd__o21ai_2 _32285_ (.A1(_10242_),
    .A2(_10244_),
    .B1(_10245_),
    .Y(_10252_));
 sky130_fd_sc_hd__o22ai_2 _32286_ (.A1(_09012_),
    .A2(_09875_),
    .B1(_09873_),
    .B2(_09874_),
    .Y(_10253_));
 sky130_fd_sc_hd__o211ai_2 _32287_ (.A1(_06401_),
    .A2(_10243_),
    .B1(_10246_),
    .C1(_10249_),
    .Y(_10254_));
 sky130_fd_sc_hd__nand3_2 _32288_ (.A(_10252_),
    .B(_10253_),
    .C(_10254_),
    .Y(_10255_));
 sky130_fd_sc_hd__nand2_2 _32289_ (.A(_10251_),
    .B(_10255_),
    .Y(_10256_));
 sky130_fd_sc_hd__nor2_2 _32290_ (.A(_09914_),
    .B(_09913_),
    .Y(_10257_));
 sky130_fd_sc_hd__nor2_2 _32291_ (.A(_09912_),
    .B(_10257_),
    .Y(_10258_));
 sky130_fd_sc_hd__nand2_2 _32292_ (.A(_10256_),
    .B(_10258_),
    .Y(_10259_));
 sky130_fd_sc_hd__o211ai_2 _32293_ (.A1(_09912_),
    .A2(_10257_),
    .B1(_10255_),
    .C1(_10251_),
    .Y(_10260_));
 sky130_fd_sc_hd__nand2_2 _32294_ (.A(_09922_),
    .B(_09924_),
    .Y(_10261_));
 sky130_fd_sc_hd__nand2_2 _32295_ (.A(_10261_),
    .B(_09919_),
    .Y(_10262_));
 sky130_fd_sc_hd__a21oi_2 _32296_ (.A1(_10259_),
    .A2(_10260_),
    .B1(_10262_),
    .Y(_10263_));
 sky130_fd_sc_hd__a21oi_2 _32297_ (.A1(_09920_),
    .A2(_09921_),
    .B1(_09908_),
    .Y(_10264_));
 sky130_fd_sc_hd__a31oi_2 _32298_ (.A1(_09920_),
    .A2(_09921_),
    .A3(_09908_),
    .B1(_09923_),
    .Y(_10265_));
 sky130_fd_sc_hd__o211a_2 _32299_ (.A1(_10264_),
    .A2(_10265_),
    .B1(_10260_),
    .C1(_10259_),
    .X(_10266_));
 sky130_fd_sc_hd__a21oi_2 _32300_ (.A1(_09952_),
    .A2(_09951_),
    .B1(_09946_),
    .Y(_10267_));
 sky130_fd_sc_hd__buf_1 _32301_ (.A(_08045_),
    .X(_10268_));
 sky130_fd_sc_hd__nand3_2 _32302_ (.A(_08315_),
    .B(_07934_),
    .C(_08447_),
    .Y(_10269_));
 sky130_fd_sc_hd__a22o_2 _32303_ (.A1(_06278_),
    .A2(_19590_),
    .B1(_06276_),
    .B2(_06728_),
    .X(_10270_));
 sky130_fd_sc_hd__o21ai_2 _32304_ (.A1(_10268_),
    .A2(_10269_),
    .B1(_10270_),
    .Y(_10271_));
 sky130_fd_sc_hd__nand2_2 _32305_ (.A(_06446_),
    .B(_08596_),
    .Y(_10272_));
 sky130_fd_sc_hd__nand2_2 _32306_ (.A(_10271_),
    .B(_10272_),
    .Y(_10273_));
 sky130_fd_sc_hd__nor2_2 _32307_ (.A(_10268_),
    .B(_10269_),
    .Y(_10274_));
 sky130_fd_sc_hd__inv_2 _32308_ (.A(_10272_),
    .Y(_10275_));
 sky130_fd_sc_hd__nand3b_2 _32309_ (.A_N(_10274_),
    .B(_10275_),
    .C(_10270_),
    .Y(_10276_));
 sky130_fd_sc_hd__nand3b_2 _32310_ (.A_N(_10267_),
    .B(_10273_),
    .C(_10276_),
    .Y(_10277_));
 sky130_fd_sc_hd__nand2_2 _32311_ (.A(_10271_),
    .B(_10275_),
    .Y(_10278_));
 sky130_fd_sc_hd__buf_1 _32312_ (.A(_08045_),
    .X(_10279_));
 sky130_fd_sc_hd__o211ai_2 _32313_ (.A1(_10279_),
    .A2(_10269_),
    .B1(_10272_),
    .C1(_10270_),
    .Y(_10280_));
 sky130_fd_sc_hd__nand3_2 _32314_ (.A(_10278_),
    .B(_10267_),
    .C(_10280_),
    .Y(_10281_));
 sky130_fd_sc_hd__nand3_2 _32315_ (.A(_09051_),
    .B(_06605_),
    .C(_09248_),
    .Y(_10282_));
 sky130_fd_sc_hd__nor2_2 _32316_ (.A(_09256_),
    .B(_10282_),
    .Y(_10283_));
 sky130_fd_sc_hd__a22o_2 _32317_ (.A1(_19371_),
    .A2(_09933_),
    .B1(_19374_),
    .B2(_07848_),
    .X(_10284_));
 sky130_fd_sc_hd__nand2_2 _32318_ (.A(_19376_),
    .B(_07849_),
    .Y(_10285_));
 sky130_fd_sc_hd__nand3b_2 _32319_ (.A_N(_10283_),
    .B(_10284_),
    .C(_10285_),
    .Y(_10286_));
 sky130_fd_sc_hd__a22oi_2 _32320_ (.A1(_19371_),
    .A2(_07852_),
    .B1(_19374_),
    .B2(_07848_),
    .Y(_10287_));
 sky130_fd_sc_hd__inv_2 _32321_ (.A(_10285_),
    .Y(_10288_));
 sky130_fd_sc_hd__o21ai_2 _32322_ (.A1(_10287_),
    .A2(_10283_),
    .B1(_10288_),
    .Y(_10289_));
 sky130_fd_sc_hd__nand2_2 _32323_ (.A(_10286_),
    .B(_10289_),
    .Y(_10290_));
 sky130_fd_sc_hd__a21oi_2 _32324_ (.A1(_10277_),
    .A2(_10281_),
    .B1(_10290_),
    .Y(_10291_));
 sky130_fd_sc_hd__a21oi_2 _32325_ (.A1(_10278_),
    .A2(_10280_),
    .B1(_10267_),
    .Y(_10292_));
 sky130_fd_sc_hd__nand2_2 _32326_ (.A(_10281_),
    .B(_10290_),
    .Y(_10293_));
 sky130_fd_sc_hd__nor2_2 _32327_ (.A(_10292_),
    .B(_10293_),
    .Y(_10294_));
 sky130_fd_sc_hd__nor2_2 _32328_ (.A(_10291_),
    .B(_10294_),
    .Y(_10295_));
 sky130_fd_sc_hd__o21ai_2 _32329_ (.A1(_10263_),
    .A2(_10266_),
    .B1(_10295_),
    .Y(_10296_));
 sky130_fd_sc_hd__inv_2 _32330_ (.A(_09890_),
    .Y(_10297_));
 sky130_fd_sc_hd__nand2_2 _32331_ (.A(_10297_),
    .B(_09888_),
    .Y(_10298_));
 sky130_fd_sc_hd__nand2_2 _32332_ (.A(_10298_),
    .B(_09887_),
    .Y(_10299_));
 sky130_fd_sc_hd__nand3_2 _32333_ (.A(_10262_),
    .B(_10259_),
    .C(_10260_),
    .Y(_10300_));
 sky130_fd_sc_hd__a21o_2 _32334_ (.A1(_10259_),
    .A2(_10260_),
    .B1(_10262_),
    .X(_10301_));
 sky130_fd_sc_hd__o211ai_2 _32335_ (.A1(_10291_),
    .A2(_10294_),
    .B1(_10300_),
    .C1(_10301_),
    .Y(_10302_));
 sky130_fd_sc_hd__nand3_2 _32336_ (.A(_10296_),
    .B(_10299_),
    .C(_10302_),
    .Y(_10303_));
 sky130_fd_sc_hd__o22ai_2 _32337_ (.A1(_10291_),
    .A2(_10294_),
    .B1(_10263_),
    .B2(_10266_),
    .Y(_10304_));
 sky130_fd_sc_hd__nand3_2 _32338_ (.A(_10301_),
    .B(_10295_),
    .C(_10300_),
    .Y(_10305_));
 sky130_fd_sc_hd__o21ai_2 _32339_ (.A1(_10297_),
    .A2(_09894_),
    .B1(_09888_),
    .Y(_10306_));
 sky130_fd_sc_hd__nand3_2 _32340_ (.A(_10304_),
    .B(_10305_),
    .C(_10306_),
    .Y(_10307_));
 sky130_fd_sc_hd__nor2_2 _32341_ (.A(_09965_),
    .B(_09929_),
    .Y(_10308_));
 sky130_fd_sc_hd__nor2_2 _32342_ (.A(_09932_),
    .B(_10308_),
    .Y(_10309_));
 sky130_fd_sc_hd__and3_2 _32343_ (.A(_10303_),
    .B(_10307_),
    .C(_10309_),
    .X(_10310_));
 sky130_fd_sc_hd__buf_1 _32344_ (.A(_10307_),
    .X(_10311_));
 sky130_fd_sc_hd__a21oi_2 _32345_ (.A1(_10303_),
    .A2(_10311_),
    .B1(_10309_),
    .Y(_10312_));
 sky130_fd_sc_hd__o2bb2ai_2 _32346_ (.A1_N(_10238_),
    .A2_N(_10241_),
    .B1(_10310_),
    .B2(_10312_),
    .Y(_10313_));
 sky130_fd_sc_hd__nand2_2 _32347_ (.A(_10303_),
    .B(_10309_),
    .Y(_10314_));
 sky130_fd_sc_hd__inv_2 _32348_ (.A(_10311_),
    .Y(_10315_));
 sky130_fd_sc_hd__o2bb2ai_2 _32349_ (.A1_N(_10311_),
    .A2_N(_10303_),
    .B1(_09932_),
    .B2(_10308_),
    .Y(_10316_));
 sky130_fd_sc_hd__o2111ai_2 _32350_ (.A1(_10314_),
    .A2(_10315_),
    .B1(_10316_),
    .C1(_10238_),
    .D1(_10241_),
    .Y(_10317_));
 sky130_fd_sc_hd__nand3_2 _32351_ (.A(_09900_),
    .B(_09974_),
    .C(_09976_),
    .Y(_10318_));
 sky130_fd_sc_hd__nand2_2 _32352_ (.A(_10318_),
    .B(_09906_),
    .Y(_10319_));
 sky130_fd_sc_hd__a21oi_2 _32353_ (.A1(_10313_),
    .A2(_10317_),
    .B1(_10319_),
    .Y(_10320_));
 sky130_fd_sc_hd__and3_2 _32354_ (.A(_09902_),
    .B(_09903_),
    .C(_09905_),
    .X(_10321_));
 sky130_fd_sc_hd__a31oi_2 _32355_ (.A1(_09900_),
    .A2(_09976_),
    .A3(_09974_),
    .B1(_10321_),
    .Y(_10322_));
 sky130_fd_sc_hd__nand2_2 _32356_ (.A(_10313_),
    .B(_10317_),
    .Y(_10323_));
 sky130_fd_sc_hd__nor2_2 _32357_ (.A(_10322_),
    .B(_10323_),
    .Y(_10324_));
 sky130_fd_sc_hd__inv_2 _32358_ (.A(_10029_),
    .Y(_10325_));
 sky130_fd_sc_hd__inv_2 _32359_ (.A(_10024_),
    .Y(_10326_));
 sky130_fd_sc_hd__nor2_2 _32360_ (.A(_10077_),
    .B(_10326_),
    .Y(_10327_));
 sky130_fd_sc_hd__nand2_2 _32361_ (.A(_09968_),
    .B(_09983_),
    .Y(_10328_));
 sky130_fd_sc_hd__nor2_2 _32362_ (.A(_10006_),
    .B(_10005_),
    .Y(_10329_));
 sky130_fd_sc_hd__nand2_2 _32363_ (.A(_05857_),
    .B(_08497_),
    .Y(_10330_));
 sky130_fd_sc_hd__nand2_2 _32364_ (.A(_06896_),
    .B(_19570_),
    .Y(_10331_));
 sky130_fd_sc_hd__nor2_2 _32365_ (.A(_10330_),
    .B(_10331_),
    .Y(_10332_));
 sky130_fd_sc_hd__and2_2 _32366_ (.A(_10330_),
    .B(_10331_),
    .X(_10333_));
 sky130_fd_sc_hd__nand2_2 _32367_ (.A(_08953_),
    .B(_08662_),
    .Y(_10334_));
 sky130_fd_sc_hd__o21ai_2 _32368_ (.A1(_10332_),
    .A2(_10333_),
    .B1(_10334_),
    .Y(_10335_));
 sky130_fd_sc_hd__inv_2 _32369_ (.A(_10334_),
    .Y(_10336_));
 sky130_fd_sc_hd__nand2_2 _32370_ (.A(_10330_),
    .B(_10331_),
    .Y(_10337_));
 sky130_fd_sc_hd__nand3b_2 _32371_ (.A_N(_10332_),
    .B(_10336_),
    .C(_10337_),
    .Y(_10338_));
 sky130_fd_sc_hd__nand2_2 _32372_ (.A(_09935_),
    .B(_09936_),
    .Y(_10339_));
 sky130_fd_sc_hd__a21o_2 _32373_ (.A1(_09939_),
    .A2(_10339_),
    .B1(_09937_),
    .X(_10340_));
 sky130_fd_sc_hd__nand3_2 _32374_ (.A(_10335_),
    .B(_10338_),
    .C(_10340_),
    .Y(_10341_));
 sky130_fd_sc_hd__o21ai_2 _32375_ (.A1(_10332_),
    .A2(_10333_),
    .B1(_10336_),
    .Y(_10342_));
 sky130_fd_sc_hd__nand3b_2 _32376_ (.A_N(_10332_),
    .B(_10334_),
    .C(_10337_),
    .Y(_10343_));
 sky130_fd_sc_hd__a21oi_2 _32377_ (.A1(_09939_),
    .A2(_10339_),
    .B1(_09937_),
    .Y(_10344_));
 sky130_fd_sc_hd__nand3_2 _32378_ (.A(_10342_),
    .B(_10343_),
    .C(_10344_),
    .Y(_10345_));
 sky130_fd_sc_hd__nor2_2 _32379_ (.A(_09993_),
    .B(_09991_),
    .Y(_10346_));
 sky130_fd_sc_hd__o2bb2ai_2 _32380_ (.A1_N(_10341_),
    .A2_N(_10345_),
    .B1(_09998_),
    .B2(_10346_),
    .Y(_10347_));
 sky130_fd_sc_hd__nor2_2 _32381_ (.A(_09998_),
    .B(_10346_),
    .Y(_10348_));
 sky130_fd_sc_hd__nand3_2 _32382_ (.A(_10341_),
    .B(_10345_),
    .C(_10348_),
    .Y(_10349_));
 sky130_fd_sc_hd__nand2_2 _32383_ (.A(_09957_),
    .B(_09959_),
    .Y(_10350_));
 sky130_fd_sc_hd__nand2_2 _32384_ (.A(_10350_),
    .B(_09954_),
    .Y(_10351_));
 sky130_fd_sc_hd__a21oi_2 _32385_ (.A1(_10347_),
    .A2(_10349_),
    .B1(_10351_),
    .Y(_10352_));
 sky130_fd_sc_hd__inv_2 _32386_ (.A(_10341_),
    .Y(_10353_));
 sky130_fd_sc_hd__nand2_2 _32387_ (.A(_10345_),
    .B(_10348_),
    .Y(_10354_));
 sky130_fd_sc_hd__o211a_2 _32388_ (.A1(_10353_),
    .A2(_10354_),
    .B1(_10347_),
    .C1(_10351_),
    .X(_10355_));
 sky130_fd_sc_hd__o22ai_2 _32389_ (.A1(_10014_),
    .A2(_10329_),
    .B1(_10352_),
    .B2(_10355_),
    .Y(_10356_));
 sky130_fd_sc_hd__nand2_2 _32390_ (.A(_10021_),
    .B(_10018_),
    .Y(_10357_));
 sky130_fd_sc_hd__nand2_2 _32391_ (.A(_10357_),
    .B(_10020_),
    .Y(_10358_));
 sky130_fd_sc_hd__nand2_2 _32392_ (.A(_10347_),
    .B(_10349_),
    .Y(_10359_));
 sky130_fd_sc_hd__a21boi_2 _32393_ (.A1(_09957_),
    .A2(_09959_),
    .B1_N(_09954_),
    .Y(_10360_));
 sky130_fd_sc_hd__nand2_2 _32394_ (.A(_10359_),
    .B(_10360_),
    .Y(_10361_));
 sky130_fd_sc_hd__nand2_2 _32395_ (.A(_10015_),
    .B(_10000_),
    .Y(_10362_));
 sky130_fd_sc_hd__inv_2 _32396_ (.A(_10362_),
    .Y(_10363_));
 sky130_fd_sc_hd__nand3_2 _32397_ (.A(_10351_),
    .B(_10347_),
    .C(_10349_),
    .Y(_10364_));
 sky130_fd_sc_hd__nand3_2 _32398_ (.A(_10361_),
    .B(_10363_),
    .C(_10364_),
    .Y(_10365_));
 sky130_fd_sc_hd__nand3_2 _32399_ (.A(_10356_),
    .B(_10358_),
    .C(_10365_),
    .Y(_10366_));
 sky130_fd_sc_hd__o21ai_2 _32400_ (.A1(_10352_),
    .A2(_10355_),
    .B1(_10363_),
    .Y(_10367_));
 sky130_fd_sc_hd__o21ai_2 _32401_ (.A1(_10018_),
    .A2(_10013_),
    .B1(_10021_),
    .Y(_10368_));
 sky130_fd_sc_hd__nand3_2 _32402_ (.A(_10361_),
    .B(_10362_),
    .C(_10364_),
    .Y(_10369_));
 sky130_fd_sc_hd__nand3_2 _32403_ (.A(_10367_),
    .B(_10368_),
    .C(_10369_),
    .Y(_10370_));
 sky130_fd_sc_hd__buf_1 _32404_ (.A(_19548_),
    .X(_10371_));
 sky130_fd_sc_hd__nand2_2 _32405_ (.A(_06219_),
    .B(_10050_),
    .Y(_10372_));
 sky130_fd_sc_hd__a21o_2 _32406_ (.A1(_05144_),
    .A2(_10371_),
    .B1(_10372_),
    .X(_10373_));
 sky130_fd_sc_hd__nand2_2 _32407_ (.A(_19401_),
    .B(_19549_),
    .Y(_10374_));
 sky130_fd_sc_hd__a21o_2 _32408_ (.A1(_19399_),
    .A2(_10050_),
    .B1(_10374_),
    .X(_10375_));
 sky130_fd_sc_hd__nand2_2 _32409_ (.A(_05116_),
    .B(_19559_),
    .Y(_10376_));
 sky130_fd_sc_hd__a21oi_2 _32410_ (.A1(_10373_),
    .A2(_10375_),
    .B1(_10376_),
    .Y(_10377_));
 sky130_fd_sc_hd__and3_2 _32411_ (.A(_10373_),
    .B(_10375_),
    .C(_10376_),
    .X(_10378_));
 sky130_fd_sc_hd__nor2_2 _32412_ (.A(_10377_),
    .B(_10378_),
    .Y(_10379_));
 sky130_fd_sc_hd__buf_1 _32413_ (.A(_08645_),
    .X(_10380_));
 sky130_fd_sc_hd__nand2_2 _32414_ (.A(_19389_),
    .B(_10380_),
    .Y(_10381_));
 sky130_fd_sc_hd__nand2_2 _32415_ (.A(_19392_),
    .B(_19562_),
    .Y(_10382_));
 sky130_fd_sc_hd__nor2_2 _32416_ (.A(_10381_),
    .B(_10382_),
    .Y(_10383_));
 sky130_fd_sc_hd__and2_2 _32417_ (.A(_10381_),
    .B(_10382_),
    .X(_10384_));
 sky130_fd_sc_hd__nand2_2 _32418_ (.A(_19404_),
    .B(_19545_),
    .Y(_10385_));
 sky130_fd_sc_hd__inv_2 _32419_ (.A(_10385_),
    .Y(_10386_));
 sky130_fd_sc_hd__o21ai_2 _32420_ (.A1(_10383_),
    .A2(_10384_),
    .B1(_10386_),
    .Y(_10387_));
 sky130_fd_sc_hd__or2_2 _32421_ (.A(_10381_),
    .B(_10382_),
    .X(_10388_));
 sky130_fd_sc_hd__nand2_2 _32422_ (.A(_10381_),
    .B(_10382_),
    .Y(_10389_));
 sky130_fd_sc_hd__nand3_2 _32423_ (.A(_10388_),
    .B(_10385_),
    .C(_10389_),
    .Y(_10390_));
 sky130_fd_sc_hd__a21oi_2 _32424_ (.A1(_10040_),
    .A2(_10041_),
    .B1(_10035_),
    .Y(_10391_));
 sky130_fd_sc_hd__nand3_2 _32425_ (.A(_10387_),
    .B(_10390_),
    .C(_10391_),
    .Y(_10392_));
 sky130_fd_sc_hd__o21ai_2 _32426_ (.A1(_10383_),
    .A2(_10384_),
    .B1(_10385_),
    .Y(_10393_));
 sky130_fd_sc_hd__nand3_2 _32427_ (.A(_10388_),
    .B(_10386_),
    .C(_10389_),
    .Y(_10394_));
 sky130_fd_sc_hd__nand3b_2 _32428_ (.A_N(_10391_),
    .B(_10393_),
    .C(_10394_),
    .Y(_10395_));
 sky130_fd_sc_hd__nand3_2 _32429_ (.A(_10379_),
    .B(_10392_),
    .C(_10395_),
    .Y(_10396_));
 sky130_fd_sc_hd__a21o_2 _32430_ (.A1(_10395_),
    .A2(_10392_),
    .B1(_10379_),
    .X(_10397_));
 sky130_fd_sc_hd__and3_2 _32431_ (.A(_10045_),
    .B(_10046_),
    .C(_10047_),
    .X(_10398_));
 sky130_fd_sc_hd__and3_2 _32432_ (.A(_10038_),
    .B(_10042_),
    .C(_10043_),
    .X(_10399_));
 sky130_fd_sc_hd__nor2_2 _32433_ (.A(_10061_),
    .B(_10399_),
    .Y(_10400_));
 sky130_fd_sc_hd__o2bb2ai_2 _32434_ (.A1_N(_10396_),
    .A2_N(_10397_),
    .B1(_10398_),
    .B2(_10400_),
    .Y(_10401_));
 sky130_fd_sc_hd__o21ai_2 _32435_ (.A1(_10059_),
    .A2(_10398_),
    .B1(_10044_),
    .Y(_10402_));
 sky130_fd_sc_hd__nand3_2 _32436_ (.A(_10402_),
    .B(_10396_),
    .C(_10397_),
    .Y(_10403_));
 sky130_fd_sc_hd__or2_2 _32437_ (.A(_10051_),
    .B(_10053_),
    .X(_10404_));
 sky130_fd_sc_hd__nand2_2 _32438_ (.A(_10057_),
    .B(_10404_),
    .Y(_10405_));
 sky130_fd_sc_hd__and3_2 _32439_ (.A(_10401_),
    .B(_10403_),
    .C(_10405_),
    .X(_10406_));
 sky130_fd_sc_hd__a21oi_2 _32440_ (.A1(_10401_),
    .A2(_10403_),
    .B1(_10405_),
    .Y(_10407_));
 sky130_fd_sc_hd__o2bb2ai_2 _32441_ (.A1_N(_10366_),
    .A2_N(_10370_),
    .B1(_10406_),
    .B2(_10407_),
    .Y(_10408_));
 sky130_fd_sc_hd__nand2_2 _32442_ (.A(_10397_),
    .B(_10396_),
    .Y(_10409_));
 sky130_fd_sc_hd__a21oi_2 _32443_ (.A1(_10061_),
    .A2(_10048_),
    .B1(_10399_),
    .Y(_10410_));
 sky130_fd_sc_hd__inv_2 _32444_ (.A(_10405_),
    .Y(_10411_));
 sky130_fd_sc_hd__a21oi_2 _32445_ (.A1(_10409_),
    .A2(_10410_),
    .B1(_10411_),
    .Y(_10412_));
 sky130_fd_sc_hd__a21oi_2 _32446_ (.A1(_10403_),
    .A2(_10412_),
    .B1(_10407_),
    .Y(_10413_));
 sky130_fd_sc_hd__nand3_2 _32447_ (.A(_10413_),
    .B(_10366_),
    .C(_10370_),
    .Y(_10414_));
 sky130_fd_sc_hd__a22oi_2 _32448_ (.A1(_09972_),
    .A2(_10328_),
    .B1(_10408_),
    .B2(_10414_),
    .Y(_10415_));
 sky130_fd_sc_hd__o211a_2 _32449_ (.A1(_09979_),
    .A2(_09984_),
    .B1(_10414_),
    .C1(_10408_),
    .X(_10416_));
 sky130_fd_sc_hd__o22ai_2 _32450_ (.A1(_10325_),
    .A2(_10327_),
    .B1(_10415_),
    .B2(_10416_),
    .Y(_10417_));
 sky130_fd_sc_hd__nand2_2 _32451_ (.A(_09980_),
    .B(_09968_),
    .Y(_10418_));
 sky130_fd_sc_hd__a21o_2 _32452_ (.A1(_10408_),
    .A2(_10414_),
    .B1(_10418_),
    .X(_10419_));
 sky130_fd_sc_hd__nor2_2 _32453_ (.A(_10325_),
    .B(_10327_),
    .Y(_10420_));
 sky130_fd_sc_hd__nand3_2 _32454_ (.A(_10418_),
    .B(_10408_),
    .C(_10414_),
    .Y(_10421_));
 sky130_fd_sc_hd__nand3_2 _32455_ (.A(_10419_),
    .B(_10420_),
    .C(_10421_),
    .Y(_10422_));
 sky130_fd_sc_hd__nand2_2 _32456_ (.A(_10417_),
    .B(_10422_),
    .Y(_10423_));
 sky130_fd_sc_hd__o21ai_2 _32457_ (.A1(_10320_),
    .A2(_10324_),
    .B1(_10423_),
    .Y(_10424_));
 sky130_fd_sc_hd__nand2_2 _32458_ (.A(_10100_),
    .B(_10080_),
    .Y(_10425_));
 sky130_fd_sc_hd__nand3_2 _32459_ (.A(_09990_),
    .B(_10094_),
    .C(_10425_),
    .Y(_10426_));
 sky130_fd_sc_hd__nand2_2 _32460_ (.A(_10426_),
    .B(_09982_),
    .Y(_10427_));
 sky130_fd_sc_hd__nor2_2 _32461_ (.A(_10073_),
    .B(_10325_),
    .Y(_10428_));
 sky130_fd_sc_hd__o22ai_2 _32462_ (.A1(_10326_),
    .A2(_10428_),
    .B1(_10415_),
    .B2(_10416_),
    .Y(_10429_));
 sky130_fd_sc_hd__nor2_2 _32463_ (.A(_10326_),
    .B(_10428_),
    .Y(_10430_));
 sky130_fd_sc_hd__nand3_2 _32464_ (.A(_10419_),
    .B(_10430_),
    .C(_10421_),
    .Y(_10431_));
 sky130_fd_sc_hd__nand2_2 _32465_ (.A(_10429_),
    .B(_10431_),
    .Y(_10432_));
 sky130_fd_sc_hd__nand2_2 _32466_ (.A(_10323_),
    .B(_10322_),
    .Y(_10433_));
 sky130_fd_sc_hd__nand3_2 _32467_ (.A(_10319_),
    .B(_10313_),
    .C(_10317_),
    .Y(_10434_));
 sky130_fd_sc_hd__nand3_2 _32468_ (.A(_10432_),
    .B(_10433_),
    .C(_10434_),
    .Y(_10435_));
 sky130_fd_sc_hd__nand3_2 _32469_ (.A(_10424_),
    .B(_10427_),
    .C(_10435_),
    .Y(_10436_));
 sky130_fd_sc_hd__o21ai_2 _32470_ (.A1(_10320_),
    .A2(_10324_),
    .B1(_10432_),
    .Y(_10437_));
 sky130_fd_sc_hd__a21oi_2 _32471_ (.A1(_09987_),
    .A2(_09989_),
    .B1(_09988_),
    .Y(_10438_));
 sky130_fd_sc_hd__a31oi_2 _32472_ (.A1(_09990_),
    .A2(_10425_),
    .A3(_10094_),
    .B1(_10438_),
    .Y(_10439_));
 sky130_fd_sc_hd__nand3_2 _32473_ (.A(_10423_),
    .B(_10433_),
    .C(_10434_),
    .Y(_10440_));
 sky130_fd_sc_hd__nand3_2 _32474_ (.A(_10437_),
    .B(_10439_),
    .C(_10440_),
    .Y(_10441_));
 sky130_fd_sc_hd__a21boi_2 _32475_ (.A1(_10070_),
    .A2(_10066_),
    .B1_N(_10063_),
    .Y(_10442_));
 sky130_fd_sc_hd__nor2_2 _32476_ (.A(_10088_),
    .B(_10100_),
    .Y(_10443_));
 sky130_fd_sc_hd__nor2_2 _32477_ (.A(_10442_),
    .B(_10443_),
    .Y(_10444_));
 sky130_fd_sc_hd__and3_2 _32478_ (.A(_10089_),
    .B(_10080_),
    .C(_10442_),
    .X(_10445_));
 sky130_fd_sc_hd__o2bb2ai_2 _32479_ (.A1_N(_10436_),
    .A2_N(_10441_),
    .B1(_10444_),
    .B2(_10445_),
    .Y(_10446_));
 sky130_fd_sc_hd__nand2_2 _32480_ (.A(_10117_),
    .B(_10096_),
    .Y(_10447_));
 sky130_fd_sc_hd__nor2_2 _32481_ (.A(_10445_),
    .B(_10444_),
    .Y(_10448_));
 sky130_fd_sc_hd__nand3_2 _32482_ (.A(_10441_),
    .B(_10436_),
    .C(_10448_),
    .Y(_10449_));
 sky130_fd_sc_hd__nand3_2 _32483_ (.A(_10446_),
    .B(_10447_),
    .C(_10449_),
    .Y(_10450_));
 sky130_fd_sc_hd__o21a_2 _32484_ (.A1(_10088_),
    .A2(_10100_),
    .B1(_10442_),
    .X(_10451_));
 sky130_fd_sc_hd__and2b_2 _32485_ (.A_N(_10442_),
    .B(_10443_),
    .X(_10452_));
 sky130_fd_sc_hd__o2bb2ai_2 _32486_ (.A1_N(_10436_),
    .A2_N(_10441_),
    .B1(_10451_),
    .B2(_10452_),
    .Y(_10453_));
 sky130_fd_sc_hd__a21boi_2 _32487_ (.A1(_10104_),
    .A2(_10112_),
    .B1_N(_10096_),
    .Y(_10454_));
 sky130_fd_sc_hd__nand3b_2 _32488_ (.A_N(_10448_),
    .B(_10441_),
    .C(_10436_),
    .Y(_10455_));
 sky130_fd_sc_hd__nand3_2 _32489_ (.A(_10453_),
    .B(_10454_),
    .C(_10455_),
    .Y(_10456_));
 sky130_fd_sc_hd__a21oi_2 _32490_ (.A1(_10450_),
    .A2(_10456_),
    .B1(_10108_),
    .Y(_10457_));
 sky130_fd_sc_hd__and3_2 _32491_ (.A(_10450_),
    .B(_10456_),
    .C(_10108_),
    .X(_10458_));
 sky130_fd_sc_hd__o21ai_2 _32492_ (.A1(_09516_),
    .A2(_10115_),
    .B1(_10122_),
    .Y(_10459_));
 sky130_fd_sc_hd__o21bai_2 _32493_ (.A1(_10457_),
    .A2(_10458_),
    .B1_N(_10459_),
    .Y(_10460_));
 sky130_fd_sc_hd__nand2_2 _32494_ (.A(_10456_),
    .B(_10108_),
    .Y(_10461_));
 sky130_fd_sc_hd__inv_2 _32495_ (.A(_10450_),
    .Y(_10462_));
 sky130_fd_sc_hd__a21o_2 _32496_ (.A1(_10450_),
    .A2(_10456_),
    .B1(_10108_),
    .X(_10463_));
 sky130_fd_sc_hd__o211ai_2 _32497_ (.A1(_10461_),
    .A2(_10462_),
    .B1(_10459_),
    .C1(_10463_),
    .Y(_10464_));
 sky130_fd_sc_hd__nand2_2 _32498_ (.A(_10460_),
    .B(_10464_),
    .Y(_10465_));
 sky130_fd_sc_hd__a21oi_2 _32499_ (.A1(_10121_),
    .A2(_10122_),
    .B1(_09517_),
    .Y(_10466_));
 sky130_fd_sc_hd__nand2_2 _32500_ (.A(_10128_),
    .B(_10129_),
    .Y(_10467_));
 sky130_fd_sc_hd__o2111ai_2 _32501_ (.A1(_10466_),
    .A2(_10467_),
    .B1(_09806_),
    .C1(_10124_),
    .D1(_09805_),
    .Y(_10468_));
 sky130_fd_sc_hd__nand2_2 _32502_ (.A(_10130_),
    .B(_09806_),
    .Y(_10469_));
 sky130_fd_sc_hd__nand2_2 _32503_ (.A(_10469_),
    .B(_10124_),
    .Y(_10470_));
 sky130_fd_sc_hd__o21ai_2 _32504_ (.A1(_10468_),
    .A2(_09813_),
    .B1(_10470_),
    .Y(_10471_));
 sky130_fd_sc_hd__xnor2_2 _32505_ (.A(_10465_),
    .B(_10471_),
    .Y(_02649_));
 sky130_fd_sc_hd__nand2_2 _32506_ (.A(_10471_),
    .B(_10460_),
    .Y(_10472_));
 sky130_fd_sc_hd__a31o_2 _32507_ (.A1(_10402_),
    .A2(_10396_),
    .A3(_10397_),
    .B1(_10412_),
    .X(_10473_));
 sky130_fd_sc_hd__inv_2 _32508_ (.A(_10473_),
    .Y(_10474_));
 sky130_fd_sc_hd__a21oi_2 _32509_ (.A1(_10419_),
    .A2(_10420_),
    .B1(_10416_),
    .Y(_10475_));
 sky130_fd_sc_hd__nor2_2 _32510_ (.A(_10474_),
    .B(_10475_),
    .Y(_10476_));
 sky130_fd_sc_hd__and3_2 _32511_ (.A(_10422_),
    .B(_10421_),
    .C(_10474_),
    .X(_10477_));
 sky130_fd_sc_hd__inv_2 _32512_ (.A(_10345_),
    .Y(_10478_));
 sky130_fd_sc_hd__nor2_2 _32513_ (.A(_10348_),
    .B(_10353_),
    .Y(_10479_));
 sky130_fd_sc_hd__a22oi_2 _32514_ (.A1(_19381_),
    .A2(_19571_),
    .B1(_19384_),
    .B2(_19568_),
    .Y(_10480_));
 sky130_fd_sc_hd__nand3_2 _32515_ (.A(_08948_),
    .B(_08949_),
    .C(_08496_),
    .Y(_10481_));
 sky130_fd_sc_hd__nor2_2 _32516_ (.A(_08487_),
    .B(_10481_),
    .Y(_10482_));
 sky130_fd_sc_hd__nand2_2 _32517_ (.A(_05764_),
    .B(_08920_),
    .Y(_10483_));
 sky130_fd_sc_hd__o21ai_2 _32518_ (.A1(_10480_),
    .A2(_10482_),
    .B1(_10483_),
    .Y(_10484_));
 sky130_fd_sc_hd__buf_1 _32519_ (.A(_08487_),
    .X(_10485_));
 sky130_fd_sc_hd__inv_2 _32520_ (.A(_10483_),
    .Y(_10486_));
 sky130_fd_sc_hd__a22o_2 _32521_ (.A1(_19381_),
    .A2(_19571_),
    .B1(_19384_),
    .B2(_19568_),
    .X(_10487_));
 sky130_fd_sc_hd__o211ai_2 _32522_ (.A1(_10485_),
    .A2(_10481_),
    .B1(_10486_),
    .C1(_10487_),
    .Y(_10488_));
 sky130_fd_sc_hd__o22ai_2 _32523_ (.A1(_09263_),
    .A2(_10282_),
    .B1(_10285_),
    .B2(_10287_),
    .Y(_10489_));
 sky130_fd_sc_hd__nand3_2 _32524_ (.A(_10484_),
    .B(_10488_),
    .C(_10489_),
    .Y(_10490_));
 sky130_fd_sc_hd__o21ai_2 _32525_ (.A1(_10480_),
    .A2(_10482_),
    .B1(_10486_),
    .Y(_10491_));
 sky130_fd_sc_hd__o211ai_2 _32526_ (.A1(_09226_),
    .A2(_10481_),
    .B1(_10483_),
    .C1(_10487_),
    .Y(_10492_));
 sky130_fd_sc_hd__nand3b_2 _32527_ (.A_N(_10489_),
    .B(_10491_),
    .C(_10492_),
    .Y(_10493_));
 sky130_fd_sc_hd__nor2_2 _32528_ (.A(_10336_),
    .B(_10332_),
    .Y(_10494_));
 sky130_fd_sc_hd__o2bb2ai_2 _32529_ (.A1_N(_10490_),
    .A2_N(_10493_),
    .B1(_10333_),
    .B2(_10494_),
    .Y(_10495_));
 sky130_fd_sc_hd__nor2_2 _32530_ (.A(_10333_),
    .B(_10494_),
    .Y(_10496_));
 sky130_fd_sc_hd__nand3_2 _32531_ (.A(_10493_),
    .B(_10490_),
    .C(_10496_),
    .Y(_10497_));
 sky130_fd_sc_hd__nand2_2 _32532_ (.A(_10293_),
    .B(_10277_),
    .Y(_10498_));
 sky130_fd_sc_hd__a21oi_2 _32533_ (.A1(_10495_),
    .A2(_10497_),
    .B1(_10498_),
    .Y(_10499_));
 sky130_fd_sc_hd__inv_2 _32534_ (.A(_10490_),
    .Y(_10500_));
 sky130_fd_sc_hd__nand2_2 _32535_ (.A(_10493_),
    .B(_10496_),
    .Y(_10501_));
 sky130_fd_sc_hd__o211a_2 _32536_ (.A1(_10500_),
    .A2(_10501_),
    .B1(_10495_),
    .C1(_10498_),
    .X(_10502_));
 sky130_fd_sc_hd__o22ai_2 _32537_ (.A1(_10478_),
    .A2(_10479_),
    .B1(_10499_),
    .B2(_10502_),
    .Y(_10503_));
 sky130_fd_sc_hd__and2_2 _32538_ (.A(_10354_),
    .B(_10341_),
    .X(_10504_));
 sky130_fd_sc_hd__a21o_2 _32539_ (.A1(_10495_),
    .A2(_10497_),
    .B1(_10498_),
    .X(_10505_));
 sky130_fd_sc_hd__nand3_2 _32540_ (.A(_10498_),
    .B(_10495_),
    .C(_10497_),
    .Y(_10506_));
 sky130_fd_sc_hd__nand3b_2 _32541_ (.A_N(_10504_),
    .B(_10505_),
    .C(_10506_),
    .Y(_10507_));
 sky130_fd_sc_hd__o21ai_2 _32542_ (.A1(_10363_),
    .A2(_10352_),
    .B1(_10364_),
    .Y(_10508_));
 sky130_fd_sc_hd__a21oi_2 _32543_ (.A1(_10503_),
    .A2(_10507_),
    .B1(_10508_),
    .Y(_10509_));
 sky130_fd_sc_hd__a21boi_2 _32544_ (.A1(_10359_),
    .A2(_10360_),
    .B1_N(_10362_),
    .Y(_10510_));
 sky130_fd_sc_hd__o211a_2 _32545_ (.A1(_10355_),
    .A2(_10510_),
    .B1(_10507_),
    .C1(_10503_),
    .X(_10511_));
 sky130_fd_sc_hd__nor2_2 _32546_ (.A(_10372_),
    .B(_10374_),
    .Y(_10512_));
 sky130_fd_sc_hd__inv_2 _32547_ (.A(\pcpi_mul.rs1[26] ),
    .Y(_10513_));
 sky130_fd_sc_hd__buf_1 _32548_ (.A(_10513_),
    .X(_10514_));
 sky130_fd_sc_hd__nand3_2 _32549_ (.A(_19389_),
    .B(_05892_),
    .C(_19558_),
    .Y(_10515_));
 sky130_fd_sc_hd__nor2_2 _32550_ (.A(_10514_),
    .B(_10515_),
    .Y(_10516_));
 sky130_fd_sc_hd__a22o_2 _32551_ (.A1(_19389_),
    .A2(_19562_),
    .B1(_19392_),
    .B2(_19558_),
    .X(_10517_));
 sky130_fd_sc_hd__inv_2 _32552_ (.A(\pcpi_mul.rs1[31] ),
    .Y(_10518_));
 sky130_fd_sc_hd__buf_1 _32553_ (.A(_10518_),
    .X(_10519_));
 sky130_fd_sc_hd__buf_1 _32554_ (.A(_10519_),
    .X(_10520_));
 sky130_fd_sc_hd__nor2_2 _32555_ (.A(_04836_),
    .B(_10520_),
    .Y(_10521_));
 sky130_fd_sc_hd__nand3b_2 _32556_ (.A_N(_10516_),
    .B(_10517_),
    .C(_10521_),
    .Y(_10522_));
 sky130_fd_sc_hd__buf_1 _32557_ (.A(_10513_),
    .X(_10523_));
 sky130_fd_sc_hd__o21ai_2 _32558_ (.A1(_10523_),
    .A2(_10515_),
    .B1(_10517_),
    .Y(_10524_));
 sky130_fd_sc_hd__o21ai_2 _32559_ (.A1(_04836_),
    .A2(_10520_),
    .B1(_10524_),
    .Y(_10525_));
 sky130_fd_sc_hd__nor2_2 _32560_ (.A(_10386_),
    .B(_10383_),
    .Y(_10526_));
 sky130_fd_sc_hd__o2bb2ai_2 _32561_ (.A1_N(_10522_),
    .A2_N(_10525_),
    .B1(_10384_),
    .B2(_10526_),
    .Y(_10527_));
 sky130_fd_sc_hd__a21o_2 _32562_ (.A1(_10386_),
    .A2(_10389_),
    .B1(_10383_),
    .X(_10528_));
 sky130_fd_sc_hd__nand3_2 _32563_ (.A(_10525_),
    .B(_10522_),
    .C(_10528_),
    .Y(_10529_));
 sky130_fd_sc_hd__nand2_2 _32564_ (.A(_10527_),
    .B(_10529_),
    .Y(_10530_));
 sky130_fd_sc_hd__inv_2 _32565_ (.A(_05736_),
    .Y(_10531_));
 sky130_fd_sc_hd__inv_2 _32566_ (.A(\pcpi_mul.rs1[29] ),
    .Y(_10532_));
 sky130_fd_sc_hd__buf_1 _32567_ (.A(_10532_),
    .X(_10533_));
 sky130_fd_sc_hd__inv_2 _32568_ (.A(\pcpi_mul.rs1[30] ),
    .Y(_10534_));
 sky130_fd_sc_hd__buf_1 _32569_ (.A(_10534_),
    .X(_10535_));
 sky130_fd_sc_hd__o22a_2 _32570_ (.A1(_10531_),
    .A2(_10533_),
    .B1(_06394_),
    .B2(_10535_),
    .X(_10536_));
 sky130_fd_sc_hd__buf_1 _32571_ (.A(_19544_),
    .X(_10537_));
 sky130_fd_sc_hd__buf_1 _32572_ (.A(\pcpi_mul.rs1[29] ),
    .X(_10538_));
 sky130_fd_sc_hd__nand2_2 _32573_ (.A(_10537_),
    .B(_10538_),
    .Y(_10539_));
 sky130_fd_sc_hd__nor2_2 _32574_ (.A(_05102_),
    .B(_10539_),
    .Y(_10540_));
 sky130_fd_sc_hd__inv_2 _32575_ (.A(_10540_),
    .Y(_10541_));
 sky130_fd_sc_hd__inv_2 _32576_ (.A(\pcpi_mul.rs1[28] ),
    .Y(_10542_));
 sky130_fd_sc_hd__buf_1 _32577_ (.A(_10542_),
    .X(_10543_));
 sky130_fd_sc_hd__nor2_2 _32578_ (.A(_05151_),
    .B(_10543_),
    .Y(_10544_));
 sky130_fd_sc_hd__nand3b_2 _32579_ (.A_N(_10536_),
    .B(_10541_),
    .C(_10544_),
    .Y(_10545_));
 sky130_fd_sc_hd__o21bai_2 _32580_ (.A1(_10540_),
    .A2(_10536_),
    .B1_N(_10544_),
    .Y(_10546_));
 sky130_fd_sc_hd__and2_2 _32581_ (.A(_10545_),
    .B(_10546_),
    .X(_10547_));
 sky130_fd_sc_hd__nand2_2 _32582_ (.A(_10530_),
    .B(_10547_),
    .Y(_10548_));
 sky130_fd_sc_hd__a21boi_2 _32583_ (.A1(_10379_),
    .A2(_10392_),
    .B1_N(_10395_),
    .Y(_10549_));
 sky130_fd_sc_hd__nand2_2 _32584_ (.A(_10545_),
    .B(_10546_),
    .Y(_10550_));
 sky130_fd_sc_hd__nand3_2 _32585_ (.A(_10550_),
    .B(_10527_),
    .C(_10529_),
    .Y(_10551_));
 sky130_fd_sc_hd__nand3_2 _32586_ (.A(_10548_),
    .B(_10549_),
    .C(_10551_),
    .Y(_10552_));
 sky130_fd_sc_hd__o21a_2 _32587_ (.A1(_10512_),
    .A2(_10377_),
    .B1(_10552_),
    .X(_10553_));
 sky130_fd_sc_hd__a21bo_2 _32588_ (.A1(_10379_),
    .A2(_10392_),
    .B1_N(_10395_),
    .X(_10554_));
 sky130_fd_sc_hd__nand3_2 _32589_ (.A(_10547_),
    .B(_10529_),
    .C(_10527_),
    .Y(_10555_));
 sky130_fd_sc_hd__nand2_2 _32590_ (.A(_10530_),
    .B(_10550_),
    .Y(_10556_));
 sky130_fd_sc_hd__nand3_2 _32591_ (.A(_10554_),
    .B(_10555_),
    .C(_10556_),
    .Y(_10557_));
 sky130_fd_sc_hd__nor2_2 _32592_ (.A(_10512_),
    .B(_10377_),
    .Y(_10558_));
 sky130_fd_sc_hd__inv_2 _32593_ (.A(_10558_),
    .Y(_10559_));
 sky130_fd_sc_hd__a21oi_2 _32594_ (.A1(_10557_),
    .A2(_10552_),
    .B1(_10559_),
    .Y(_10560_));
 sky130_fd_sc_hd__a21oi_2 _32595_ (.A1(_10553_),
    .A2(_10557_),
    .B1(_10560_),
    .Y(_10561_));
 sky130_fd_sc_hd__o21ai_2 _32596_ (.A1(_10509_),
    .A2(_10511_),
    .B1(_10561_),
    .Y(_10562_));
 sky130_fd_sc_hd__a21boi_2 _32597_ (.A1(_10303_),
    .A2(_10309_),
    .B1_N(_10311_),
    .Y(_10563_));
 sky130_fd_sc_hd__a21o_2 _32598_ (.A1(_10553_),
    .A2(_10557_),
    .B1(_10560_),
    .X(_10564_));
 sky130_fd_sc_hd__a21o_2 _32599_ (.A1(_10503_),
    .A2(_10507_),
    .B1(_10508_),
    .X(_10565_));
 sky130_fd_sc_hd__nand3_2 _32600_ (.A(_10503_),
    .B(_10508_),
    .C(_10507_),
    .Y(_10566_));
 sky130_fd_sc_hd__nand3_2 _32601_ (.A(_10564_),
    .B(_10565_),
    .C(_10566_),
    .Y(_10567_));
 sky130_fd_sc_hd__nand3_2 _32602_ (.A(_10562_),
    .B(_10563_),
    .C(_10567_),
    .Y(_10568_));
 sky130_fd_sc_hd__buf_1 _32603_ (.A(_10568_),
    .X(_10569_));
 sky130_fd_sc_hd__nand2_2 _32604_ (.A(_10557_),
    .B(_10552_),
    .Y(_10570_));
 sky130_fd_sc_hd__nor2_2 _32605_ (.A(_10558_),
    .B(_10570_),
    .Y(_10571_));
 sky130_fd_sc_hd__o22ai_2 _32606_ (.A1(_10571_),
    .A2(_10560_),
    .B1(_10509_),
    .B2(_10511_),
    .Y(_10572_));
 sky130_fd_sc_hd__nand2_2 _32607_ (.A(_10314_),
    .B(_10311_),
    .Y(_10573_));
 sky130_fd_sc_hd__nand3_2 _32608_ (.A(_10565_),
    .B(_10561_),
    .C(_10566_),
    .Y(_10574_));
 sky130_fd_sc_hd__nand3_2 _32609_ (.A(_10572_),
    .B(_10573_),
    .C(_10574_),
    .Y(_10575_));
 sky130_fd_sc_hd__buf_1 _32610_ (.A(_10575_),
    .X(_10576_));
 sky130_fd_sc_hd__inv_2 _32611_ (.A(_10370_),
    .Y(_10577_));
 sky130_fd_sc_hd__a21o_2 _32612_ (.A1(_10366_),
    .A2(_10413_),
    .B1(_10577_),
    .X(_10578_));
 sky130_fd_sc_hd__a21oi_2 _32613_ (.A1(_10569_),
    .A2(_10576_),
    .B1(_10578_),
    .Y(_10579_));
 sky130_fd_sc_hd__and3_2 _32614_ (.A(_10568_),
    .B(_10575_),
    .C(_10578_),
    .X(_10580_));
 sky130_fd_sc_hd__nand3_2 _32615_ (.A(_09008_),
    .B(_09019_),
    .C(_06935_),
    .Y(_10581_));
 sky130_fd_sc_hd__nand2_2 _32616_ (.A(_19360_),
    .B(_06750_),
    .Y(_10582_));
 sky130_fd_sc_hd__a22oi_2 _32617_ (.A1(_09008_),
    .A2(_06935_),
    .B1(_09009_),
    .B2(_06557_),
    .Y(_10583_));
 sky130_fd_sc_hd__nor2_2 _32618_ (.A(_10582_),
    .B(_10583_),
    .Y(_10584_));
 sky130_fd_sc_hd__o21ai_2 _32619_ (.A1(_06959_),
    .A2(_10581_),
    .B1(_10584_),
    .Y(_10585_));
 sky130_fd_sc_hd__o21ai_2 _32620_ (.A1(_10212_),
    .A2(_10217_),
    .B1(_10209_),
    .Y(_10586_));
 sky130_fd_sc_hd__nor2_2 _32621_ (.A(_06959_),
    .B(_10581_),
    .Y(_10587_));
 sky130_fd_sc_hd__o21ai_2 _32622_ (.A1(_10583_),
    .A2(_10587_),
    .B1(_10582_),
    .Y(_10588_));
 sky130_fd_sc_hd__nand3_2 _32623_ (.A(_10585_),
    .B(_10586_),
    .C(_10588_),
    .Y(_10589_));
 sky130_fd_sc_hd__o21bai_2 _32624_ (.A1(_10583_),
    .A2(_10587_),
    .B1_N(_10582_),
    .Y(_10590_));
 sky130_fd_sc_hd__a21oi_2 _32625_ (.A1(_10211_),
    .A2(_10213_),
    .B1(_10218_),
    .Y(_10591_));
 sky130_fd_sc_hd__a22o_2 _32626_ (.A1(_19355_),
    .A2(_06388_),
    .B1(_19358_),
    .B2(_06954_),
    .X(_10592_));
 sky130_fd_sc_hd__o211ai_2 _32627_ (.A1(_06959_),
    .A2(_10581_),
    .B1(_10582_),
    .C1(_10592_),
    .Y(_10593_));
 sky130_fd_sc_hd__nand3_2 _32628_ (.A(_10590_),
    .B(_10591_),
    .C(_10593_),
    .Y(_10594_));
 sky130_fd_sc_hd__nand2_2 _32629_ (.A(_10589_),
    .B(_10594_),
    .Y(_10595_));
 sky130_fd_sc_hd__nor2_2 _32630_ (.A(_10245_),
    .B(_10242_),
    .Y(_10596_));
 sky130_fd_sc_hd__nor2_2 _32631_ (.A(_10244_),
    .B(_10596_),
    .Y(_10597_));
 sky130_fd_sc_hd__nand2_2 _32632_ (.A(_10595_),
    .B(_10597_),
    .Y(_10598_));
 sky130_fd_sc_hd__nand3b_2 _32633_ (.A_N(_10597_),
    .B(_10589_),
    .C(_10594_),
    .Y(_10599_));
 sky130_fd_sc_hd__nand2_2 _32634_ (.A(_10260_),
    .B(_10255_),
    .Y(_10600_));
 sky130_fd_sc_hd__a21oi_2 _32635_ (.A1(_10598_),
    .A2(_10599_),
    .B1(_10600_),
    .Y(_10601_));
 sky130_fd_sc_hd__inv_2 _32636_ (.A(_10255_),
    .Y(_10602_));
 sky130_fd_sc_hd__o21a_2 _32637_ (.A1(_09912_),
    .A2(_10257_),
    .B1(_10251_),
    .X(_10603_));
 sky130_fd_sc_hd__o211a_2 _32638_ (.A1(_10602_),
    .A2(_10603_),
    .B1(_10599_),
    .C1(_10598_),
    .X(_10604_));
 sky130_fd_sc_hd__nand2_2 _32639_ (.A(_07012_),
    .B(_19588_),
    .Y(_10605_));
 sky130_fd_sc_hd__nand2_2 _32640_ (.A(_06443_),
    .B(_07156_),
    .Y(_10606_));
 sky130_fd_sc_hd__nor2_2 _32641_ (.A(_10605_),
    .B(_10606_),
    .Y(_10607_));
 sky130_fd_sc_hd__and2_2 _32642_ (.A(_10605_),
    .B(_10606_),
    .X(_10608_));
 sky130_fd_sc_hd__nand2_2 _32643_ (.A(_06628_),
    .B(_19582_),
    .Y(_10609_));
 sky130_fd_sc_hd__inv_2 _32644_ (.A(_10609_),
    .Y(_10610_));
 sky130_fd_sc_hd__o21ai_2 _32645_ (.A1(_10607_),
    .A2(_10608_),
    .B1(_10610_),
    .Y(_10611_));
 sky130_fd_sc_hd__nand2_2 _32646_ (.A(_10605_),
    .B(_10606_),
    .Y(_10612_));
 sky130_fd_sc_hd__nand3b_2 _32647_ (.A_N(_10607_),
    .B(_10612_),
    .C(_10609_),
    .Y(_10613_));
 sky130_fd_sc_hd__a21oi_2 _32648_ (.A1(_10270_),
    .A2(_10275_),
    .B1(_10274_),
    .Y(_10614_));
 sky130_fd_sc_hd__a21oi_2 _32649_ (.A1(_10611_),
    .A2(_10613_),
    .B1(_10614_),
    .Y(_10615_));
 sky130_fd_sc_hd__nand3_2 _32650_ (.A(_10611_),
    .B(_10613_),
    .C(_10614_),
    .Y(_10616_));
 sky130_fd_sc_hd__inv_2 _32651_ (.A(_10616_),
    .Y(_10617_));
 sky130_fd_sc_hd__nand2_2 _32652_ (.A(_07203_),
    .B(_07594_),
    .Y(_10618_));
 sky130_fd_sc_hd__nand2_2 _32653_ (.A(_07034_),
    .B(_07605_),
    .Y(_10619_));
 sky130_fd_sc_hd__nor2_2 _32654_ (.A(_10618_),
    .B(_10619_),
    .Y(_10620_));
 sky130_fd_sc_hd__nand2_2 _32655_ (.A(_10618_),
    .B(_10619_),
    .Y(_10621_));
 sky130_fd_sc_hd__inv_2 _32656_ (.A(_10621_),
    .Y(_10622_));
 sky130_fd_sc_hd__nand2_2 _32657_ (.A(_19376_),
    .B(_09994_),
    .Y(_10623_));
 sky130_fd_sc_hd__inv_2 _32658_ (.A(_10623_),
    .Y(_10624_));
 sky130_fd_sc_hd__o21ai_2 _32659_ (.A1(_10620_),
    .A2(_10622_),
    .B1(_10624_),
    .Y(_10625_));
 sky130_fd_sc_hd__nand3b_2 _32660_ (.A_N(_10620_),
    .B(_10623_),
    .C(_10621_),
    .Y(_10626_));
 sky130_fd_sc_hd__nand2_2 _32661_ (.A(_10625_),
    .B(_10626_),
    .Y(_10627_));
 sky130_fd_sc_hd__o21ai_2 _32662_ (.A1(_10615_),
    .A2(_10617_),
    .B1(_10627_),
    .Y(_10628_));
 sky130_fd_sc_hd__inv_2 _32663_ (.A(_10627_),
    .Y(_10629_));
 sky130_fd_sc_hd__a21o_2 _32664_ (.A1(_10611_),
    .A2(_10613_),
    .B1(_10614_),
    .X(_10630_));
 sky130_fd_sc_hd__nand3_2 _32665_ (.A(_10629_),
    .B(_10616_),
    .C(_10630_),
    .Y(_10631_));
 sky130_fd_sc_hd__nand2_2 _32666_ (.A(_10628_),
    .B(_10631_),
    .Y(_10632_));
 sky130_fd_sc_hd__o21ai_2 _32667_ (.A1(_10601_),
    .A2(_10604_),
    .B1(_10632_),
    .Y(_10633_));
 sky130_fd_sc_hd__inv_2 _32668_ (.A(_10232_),
    .Y(_10634_));
 sky130_fd_sc_hd__o21a_2 _32669_ (.A1(_10634_),
    .A2(_10223_),
    .B1(_10230_),
    .X(_10635_));
 sky130_fd_sc_hd__nand2_2 _32670_ (.A(_10627_),
    .B(_10616_),
    .Y(_10636_));
 sky130_fd_sc_hd__o21ai_2 _32671_ (.A1(_10615_),
    .A2(_10617_),
    .B1(_10629_),
    .Y(_10637_));
 sky130_fd_sc_hd__o21ai_2 _32672_ (.A1(_10615_),
    .A2(_10636_),
    .B1(_10637_),
    .Y(_10638_));
 sky130_fd_sc_hd__a21o_2 _32673_ (.A1(_10598_),
    .A2(_10599_),
    .B1(_10600_),
    .X(_10639_));
 sky130_fd_sc_hd__nand3_2 _32674_ (.A(_10600_),
    .B(_10598_),
    .C(_10599_),
    .Y(_10640_));
 sky130_fd_sc_hd__nand3_2 _32675_ (.A(_10638_),
    .B(_10639_),
    .C(_10640_),
    .Y(_10641_));
 sky130_fd_sc_hd__nand3_2 _32676_ (.A(_10633_),
    .B(_10635_),
    .C(_10641_),
    .Y(_10642_));
 sky130_fd_sc_hd__a21oi_2 _32677_ (.A1(_10630_),
    .A2(_10616_),
    .B1(_10627_),
    .Y(_10643_));
 sky130_fd_sc_hd__nor2_2 _32678_ (.A(_10615_),
    .B(_10636_),
    .Y(_10644_));
 sky130_fd_sc_hd__o22ai_2 _32679_ (.A1(_10643_),
    .A2(_10644_),
    .B1(_10601_),
    .B2(_10604_),
    .Y(_10645_));
 sky130_fd_sc_hd__o21ai_2 _32680_ (.A1(_10634_),
    .A2(_10223_),
    .B1(_10230_),
    .Y(_10646_));
 sky130_fd_sc_hd__nand3_2 _32681_ (.A(_10639_),
    .B(_10632_),
    .C(_10640_),
    .Y(_10647_));
 sky130_fd_sc_hd__nand3_2 _32682_ (.A(_10645_),
    .B(_10646_),
    .C(_10647_),
    .Y(_10648_));
 sky130_fd_sc_hd__nand2_2 _32683_ (.A(_10301_),
    .B(_10295_),
    .Y(_10649_));
 sky130_fd_sc_hd__nand2_2 _32684_ (.A(_10649_),
    .B(_10300_),
    .Y(_10650_));
 sky130_fd_sc_hd__a21oi_2 _32685_ (.A1(_10642_),
    .A2(_10648_),
    .B1(_10650_),
    .Y(_10651_));
 sky130_fd_sc_hd__inv_2 _32686_ (.A(_10650_),
    .Y(_10652_));
 sky130_fd_sc_hd__nand2_2 _32687_ (.A(_10642_),
    .B(_10648_),
    .Y(_10653_));
 sky130_fd_sc_hd__nor2_2 _32688_ (.A(_10652_),
    .B(_10653_),
    .Y(_10654_));
 sky130_fd_sc_hd__buf_1 _32689_ (.A(_09094_),
    .X(_10655_));
 sky130_fd_sc_hd__buf_1 _32690_ (.A(_08791_),
    .X(_10656_));
 sky130_fd_sc_hd__a22oi_2 _32691_ (.A1(_10655_),
    .A2(_19617_),
    .B1(_10656_),
    .B2(_19614_),
    .Y(_10657_));
 sky130_fd_sc_hd__nand3_2 _32692_ (.A(_08391_),
    .B(_09614_),
    .C(_06162_),
    .Y(_10658_));
 sky130_fd_sc_hd__nor2_2 _32693_ (.A(_06494_),
    .B(_10658_),
    .Y(_10659_));
 sky130_fd_sc_hd__nand2_2 _32694_ (.A(_08388_),
    .B(_05598_),
    .Y(_10660_));
 sky130_fd_sc_hd__inv_2 _32695_ (.A(_10660_),
    .Y(_10661_));
 sky130_fd_sc_hd__o21ai_2 _32696_ (.A1(_10657_),
    .A2(_10659_),
    .B1(_10661_),
    .Y(_10662_));
 sky130_fd_sc_hd__a21oi_2 _32697_ (.A1(_10201_),
    .A2(_10200_),
    .B1(_10196_),
    .Y(_10663_));
 sky130_fd_sc_hd__a22o_2 _32698_ (.A1(_08396_),
    .A2(_05613_),
    .B1(_08383_),
    .B2(_07210_),
    .X(_10664_));
 sky130_fd_sc_hd__o211ai_2 _32699_ (.A1(_06505_),
    .A2(_10658_),
    .B1(_10660_),
    .C1(_10664_),
    .Y(_10665_));
 sky130_fd_sc_hd__nand3_2 _32700_ (.A(_10662_),
    .B(_10663_),
    .C(_10665_),
    .Y(_10666_));
 sky130_fd_sc_hd__nor2_2 _32701_ (.A(_10197_),
    .B(_10194_),
    .Y(_10667_));
 sky130_fd_sc_hd__o211ai_2 _32702_ (.A1(_06505_),
    .A2(_10658_),
    .B1(_10661_),
    .C1(_10664_),
    .Y(_10668_));
 sky130_fd_sc_hd__o21ai_2 _32703_ (.A1(_10657_),
    .A2(_10659_),
    .B1(_10660_),
    .Y(_10669_));
 sky130_fd_sc_hd__o211ai_2 _32704_ (.A1(_10196_),
    .A2(_10667_),
    .B1(_10668_),
    .C1(_10669_),
    .Y(_10670_));
 sky130_fd_sc_hd__nand2_2 _32705_ (.A(_09101_),
    .B(_05911_),
    .Y(_10671_));
 sky130_fd_sc_hd__nand2_2 _32706_ (.A(_19350_),
    .B(_06726_),
    .Y(_10672_));
 sky130_fd_sc_hd__nor2_2 _32707_ (.A(_10671_),
    .B(_10672_),
    .Y(_10673_));
 sky130_fd_sc_hd__and2_2 _32708_ (.A(_10671_),
    .B(_10672_),
    .X(_10674_));
 sky130_fd_sc_hd__nand2_2 _32709_ (.A(_08407_),
    .B(_06724_),
    .Y(_10675_));
 sky130_fd_sc_hd__o21a_2 _32710_ (.A1(_10673_),
    .A2(_10674_),
    .B1(_10675_),
    .X(_10676_));
 sky130_fd_sc_hd__or2_2 _32711_ (.A(_10671_),
    .B(_10672_),
    .X(_10677_));
 sky130_fd_sc_hd__inv_2 _32712_ (.A(_10675_),
    .Y(_10678_));
 sky130_fd_sc_hd__nand2_2 _32713_ (.A(_10671_),
    .B(_10672_),
    .Y(_10679_));
 sky130_fd_sc_hd__and3_2 _32714_ (.A(_10677_),
    .B(_10678_),
    .C(_10679_),
    .X(_10680_));
 sky130_fd_sc_hd__o2bb2ai_2 _32715_ (.A1_N(_10666_),
    .A2_N(_10670_),
    .B1(_10676_),
    .B2(_10680_),
    .Y(_10681_));
 sky130_fd_sc_hd__o21ai_2 _32716_ (.A1(_10673_),
    .A2(_10674_),
    .B1(_10678_),
    .Y(_10682_));
 sky130_fd_sc_hd__nand3_2 _32717_ (.A(_10677_),
    .B(_10675_),
    .C(_10679_),
    .Y(_10683_));
 sky130_fd_sc_hd__nand2_2 _32718_ (.A(_10682_),
    .B(_10683_),
    .Y(_10684_));
 sky130_fd_sc_hd__nand3_2 _32719_ (.A(_10684_),
    .B(_10670_),
    .C(_10666_),
    .Y(_10685_));
 sky130_fd_sc_hd__nand2_2 _32720_ (.A(_10179_),
    .B(_10174_),
    .Y(_10686_));
 sky130_fd_sc_hd__a21oi_2 _32721_ (.A1(_10681_),
    .A2(_10685_),
    .B1(_10686_),
    .Y(_10687_));
 sky130_fd_sc_hd__a31oi_2 _32722_ (.A1(_10163_),
    .A2(_10165_),
    .A3(_10168_),
    .B1(_10176_),
    .Y(_10688_));
 sky130_fd_sc_hd__inv_2 _32723_ (.A(_10174_),
    .Y(_10689_));
 sky130_fd_sc_hd__o211a_2 _32724_ (.A1(_10688_),
    .A2(_10689_),
    .B1(_10685_),
    .C1(_10681_),
    .X(_10690_));
 sky130_fd_sc_hd__nand2_2 _32725_ (.A(_10207_),
    .B(_10221_),
    .Y(_10691_));
 sky130_fd_sc_hd__nand2_2 _32726_ (.A(_10691_),
    .B(_10203_),
    .Y(_10692_));
 sky130_fd_sc_hd__o21bai_2 _32727_ (.A1(_10687_),
    .A2(_10690_),
    .B1_N(_10692_),
    .Y(_10693_));
 sky130_fd_sc_hd__nand2_2 _32728_ (.A(_10681_),
    .B(_10685_),
    .Y(_10694_));
 sky130_fd_sc_hd__nor2_2 _32729_ (.A(_10688_),
    .B(_10689_),
    .Y(_10695_));
 sky130_fd_sc_hd__nand2_2 _32730_ (.A(_10694_),
    .B(_10695_),
    .Y(_10696_));
 sky130_fd_sc_hd__nand3_2 _32731_ (.A(_10686_),
    .B(_10685_),
    .C(_10681_),
    .Y(_10697_));
 sky130_fd_sc_hd__nand3_2 _32732_ (.A(_10696_),
    .B(_10697_),
    .C(_10692_),
    .Y(_10698_));
 sky130_fd_sc_hd__buf_1 _32733_ (.A(\pcpi_mul.rs2[31] ),
    .X(_10699_));
 sky130_fd_sc_hd__buf_1 _32734_ (.A(_10699_),
    .X(_10700_));
 sky130_fd_sc_hd__a22oi_2 _32735_ (.A1(_10700_),
    .A2(_19641_),
    .B1(_19312_),
    .B2(_19637_),
    .Y(_10701_));
 sky130_fd_sc_hd__and4_2 _32736_ (.A(_10700_),
    .B(_19312_),
    .C(_05124_),
    .D(_06598_),
    .X(_10702_));
 sky130_fd_sc_hd__nand2_2 _32737_ (.A(_09841_),
    .B(\pcpi_mul.rs2[28] ),
    .Y(_10703_));
 sky130_fd_sc_hd__buf_1 _32738_ (.A(_10703_),
    .X(_10704_));
 sky130_fd_sc_hd__buf_1 _32739_ (.A(_10704_),
    .X(_10705_));
 sky130_fd_sc_hd__nand2_2 _32740_ (.A(_19323_),
    .B(_06501_),
    .Y(_10706_));
 sky130_fd_sc_hd__a22o_2 _32741_ (.A1(_10146_),
    .A2(_05120_),
    .B1(_09838_),
    .B2(_06622_),
    .X(_10707_));
 sky130_fd_sc_hd__o211ai_2 _32742_ (.A1(_05147_),
    .A2(_10705_),
    .B1(_10706_),
    .C1(_10707_),
    .Y(_10708_));
 sky130_fd_sc_hd__a22oi_2 _32743_ (.A1(_10139_),
    .A2(_19634_),
    .B1(_19320_),
    .B2(_19631_),
    .Y(_10709_));
 sky130_fd_sc_hd__nor2_2 _32744_ (.A(_05147_),
    .B(_10704_),
    .Y(_10710_));
 sky130_fd_sc_hd__inv_2 _32745_ (.A(_10706_),
    .Y(_10711_));
 sky130_fd_sc_hd__o21ai_2 _32746_ (.A1(_10709_),
    .A2(_10710_),
    .B1(_10711_),
    .Y(_10712_));
 sky130_fd_sc_hd__o211ai_2 _32747_ (.A1(_10701_),
    .A2(_10702_),
    .B1(_10708_),
    .C1(_10712_),
    .Y(_10713_));
 sky130_fd_sc_hd__nand2_2 _32748_ (.A(_10707_),
    .B(_10711_),
    .Y(_10714_));
 sky130_fd_sc_hd__nor2_2 _32749_ (.A(_10701_),
    .B(_10702_),
    .Y(_10715_));
 sky130_fd_sc_hd__o21ai_2 _32750_ (.A1(_10709_),
    .A2(_10710_),
    .B1(_10706_),
    .Y(_10716_));
 sky130_fd_sc_hd__o211ai_2 _32751_ (.A1(_10710_),
    .A2(_10714_),
    .B1(_10715_),
    .C1(_10716_),
    .Y(_10717_));
 sky130_fd_sc_hd__inv_2 _32752_ (.A(_10154_),
    .Y(_10718_));
 sky130_fd_sc_hd__nand2_2 _32753_ (.A(_10149_),
    .B(_10145_),
    .Y(_10719_));
 sky130_fd_sc_hd__o2bb2ai_2 _32754_ (.A1_N(_10713_),
    .A2_N(_10717_),
    .B1(_10718_),
    .B2(_10719_),
    .Y(_10720_));
 sky130_fd_sc_hd__nand2_2 _32755_ (.A(_10142_),
    .B(_10144_),
    .Y(_10721_));
 sky130_fd_sc_hd__o211a_2 _32756_ (.A1(_10148_),
    .A2(_10721_),
    .B1(_10154_),
    .C1(_10149_),
    .X(_10722_));
 sky130_fd_sc_hd__nand3_2 _32757_ (.A(_10722_),
    .B(_10713_),
    .C(_10717_),
    .Y(_10723_));
 sky130_fd_sc_hd__nand3_2 _32758_ (.A(_09339_),
    .B(_09120_),
    .C(_05345_),
    .Y(_10724_));
 sky130_fd_sc_hd__nor2_2 _32759_ (.A(_05261_),
    .B(_10724_),
    .Y(_10725_));
 sky130_fd_sc_hd__a22o_2 _32760_ (.A1(_09819_),
    .A2(_05269_),
    .B1(_09827_),
    .B2(_06606_),
    .X(_10726_));
 sky130_fd_sc_hd__nand2_2 _32761_ (.A(\pcpi_mul.rs2[24] ),
    .B(_06808_),
    .Y(_10727_));
 sky130_fd_sc_hd__inv_2 _32762_ (.A(_10727_),
    .Y(_10728_));
 sky130_fd_sc_hd__nand2_2 _32763_ (.A(_10726_),
    .B(_10728_),
    .Y(_10729_));
 sky130_fd_sc_hd__o21ai_2 _32764_ (.A1(_10143_),
    .A2(_10147_),
    .B1(_10140_),
    .Y(_10730_));
 sky130_fd_sc_hd__a22oi_2 _32765_ (.A1(_09819_),
    .A2(_06502_),
    .B1(_19331_),
    .B2(_06614_),
    .Y(_10731_));
 sky130_fd_sc_hd__o21ai_2 _32766_ (.A1(_10731_),
    .A2(_10725_),
    .B1(_10727_),
    .Y(_10732_));
 sky130_fd_sc_hd__o211ai_2 _32767_ (.A1(_10725_),
    .A2(_10729_),
    .B1(_10730_),
    .C1(_10732_),
    .Y(_10733_));
 sky130_fd_sc_hd__o21ai_2 _32768_ (.A1(_10731_),
    .A2(_10725_),
    .B1(_10728_),
    .Y(_10734_));
 sky130_fd_sc_hd__a21oi_2 _32769_ (.A1(_10142_),
    .A2(_10144_),
    .B1(_10148_),
    .Y(_10735_));
 sky130_fd_sc_hd__o211ai_2 _32770_ (.A1(_05501_),
    .A2(_10724_),
    .B1(_10727_),
    .C1(_10726_),
    .Y(_10736_));
 sky130_fd_sc_hd__nand3_2 _32771_ (.A(_10734_),
    .B(_10735_),
    .C(_10736_),
    .Y(_10737_));
 sky130_fd_sc_hd__a21o_2 _32772_ (.A1(_10167_),
    .A2(_10162_),
    .B1(_10160_),
    .X(_10738_));
 sky130_fd_sc_hd__a21oi_2 _32773_ (.A1(_10733_),
    .A2(_10737_),
    .B1(_10738_),
    .Y(_10739_));
 sky130_fd_sc_hd__a21oi_2 _32774_ (.A1(_10734_),
    .A2(_10736_),
    .B1(_10735_),
    .Y(_10740_));
 sky130_fd_sc_hd__nand2_2 _32775_ (.A(_10737_),
    .B(_10738_),
    .Y(_10741_));
 sky130_fd_sc_hd__nor2_2 _32776_ (.A(_10740_),
    .B(_10741_),
    .Y(_10742_));
 sky130_fd_sc_hd__o2bb2ai_2 _32777_ (.A1_N(_10720_),
    .A2_N(_10723_),
    .B1(_10739_),
    .B2(_10742_),
    .Y(_10743_));
 sky130_fd_sc_hd__a21o_2 _32778_ (.A1(_10733_),
    .A2(_10737_),
    .B1(_10738_),
    .X(_10744_));
 sky130_fd_sc_hd__o2111ai_2 _32779_ (.A1(_10740_),
    .A2(_10741_),
    .B1(_10723_),
    .C1(_10720_),
    .D1(_10744_),
    .Y(_10745_));
 sky130_fd_sc_hd__a21oi_2 _32780_ (.A1(_10743_),
    .A2(_10745_),
    .B1(_10183_),
    .Y(_10746_));
 sky130_fd_sc_hd__nor2_2 _32781_ (.A(_10181_),
    .B(_10182_),
    .Y(_10747_));
 sky130_fd_sc_hd__o2111a_2 _32782_ (.A1(_10175_),
    .A2(_10176_),
    .B1(_10747_),
    .C1(_10745_),
    .D1(_10743_),
    .X(_10748_));
 sky130_fd_sc_hd__o2bb2ai_2 _32783_ (.A1_N(_10693_),
    .A2_N(_10698_),
    .B1(_10746_),
    .B2(_10748_),
    .Y(_10749_));
 sky130_fd_sc_hd__nand2_2 _32784_ (.A(_10696_),
    .B(_10692_),
    .Y(_10750_));
 sky130_fd_sc_hd__nand3_2 _32785_ (.A(_10743_),
    .B(_10183_),
    .C(_10745_),
    .Y(_10751_));
 sky130_fd_sc_hd__o2bb2ai_2 _32786_ (.A1_N(_10745_),
    .A2_N(_10743_),
    .B1(_10181_),
    .B2(_10185_),
    .Y(_10752_));
 sky130_fd_sc_hd__o2111ai_2 _32787_ (.A1(_10690_),
    .A2(_10750_),
    .B1(_10751_),
    .C1(_10693_),
    .D1(_10752_),
    .Y(_10753_));
 sky130_fd_sc_hd__nand3_2 _32788_ (.A(_10184_),
    .B(_10227_),
    .C(_10233_),
    .Y(_10754_));
 sky130_fd_sc_hd__nand2_2 _32789_ (.A(_10754_),
    .B(_10188_),
    .Y(_10755_));
 sky130_fd_sc_hd__a21oi_2 _32790_ (.A1(_10749_),
    .A2(_10753_),
    .B1(_10755_),
    .Y(_10756_));
 sky130_fd_sc_hd__nand3_2 _32791_ (.A(_10693_),
    .B(_10698_),
    .C(_10751_),
    .Y(_10757_));
 sky130_fd_sc_hd__o211a_2 _32792_ (.A1(_10746_),
    .A2(_10757_),
    .B1(_10749_),
    .C1(_10755_),
    .X(_10758_));
 sky130_fd_sc_hd__o22ai_2 _32793_ (.A1(_10651_),
    .A2(_10654_),
    .B1(_10756_),
    .B2(_10758_),
    .Y(_10759_));
 sky130_fd_sc_hd__a22oi_2 _32794_ (.A1(_10693_),
    .A2(_10698_),
    .B1(_10752_),
    .B2(_10751_),
    .Y(_10760_));
 sky130_fd_sc_hd__o2bb2ai_2 _32795_ (.A1_N(_10188_),
    .A2_N(_10754_),
    .B1(_10746_),
    .B2(_10757_),
    .Y(_10761_));
 sky130_fd_sc_hd__nand2_2 _32796_ (.A(_10653_),
    .B(_10652_),
    .Y(_10762_));
 sky130_fd_sc_hd__nand3_2 _32797_ (.A(_10642_),
    .B(_10648_),
    .C(_10650_),
    .Y(_10763_));
 sky130_fd_sc_hd__o2111a_2 _32798_ (.A1(_10690_),
    .A2(_10750_),
    .B1(_10751_),
    .C1(_10693_),
    .D1(_10752_),
    .X(_10764_));
 sky130_fd_sc_hd__o21bai_2 _32799_ (.A1(_10760_),
    .A2(_10764_),
    .B1_N(_10755_),
    .Y(_10765_));
 sky130_fd_sc_hd__o2111ai_2 _32800_ (.A1(_10760_),
    .A2(_10761_),
    .B1(_10762_),
    .C1(_10763_),
    .D1(_10765_),
    .Y(_10766_));
 sky130_fd_sc_hd__inv_2 _32801_ (.A(_10235_),
    .Y(_10767_));
 sky130_fd_sc_hd__nand2_2 _32802_ (.A(_10135_),
    .B(_10237_),
    .Y(_10768_));
 sky130_fd_sc_hd__a21oi_2 _32803_ (.A1(_10235_),
    .A2(_10237_),
    .B1(_10135_),
    .Y(_10769_));
 sky130_fd_sc_hd__nand3_2 _32804_ (.A(_10303_),
    .B(_10311_),
    .C(_10309_),
    .Y(_10770_));
 sky130_fd_sc_hd__nand2_2 _32805_ (.A(_10316_),
    .B(_10770_),
    .Y(_10771_));
 sky130_fd_sc_hd__o22ai_2 _32806_ (.A1(_10767_),
    .A2(_10768_),
    .B1(_10769_),
    .B2(_10771_),
    .Y(_10772_));
 sky130_fd_sc_hd__a21oi_2 _32807_ (.A1(_10759_),
    .A2(_10766_),
    .B1(_10772_),
    .Y(_10773_));
 sky130_fd_sc_hd__nand3_2 _32808_ (.A(_10755_),
    .B(_10749_),
    .C(_10753_),
    .Y(_10774_));
 sky130_fd_sc_hd__nand3_2 _32809_ (.A(_10762_),
    .B(_10774_),
    .C(_10763_),
    .Y(_10775_));
 sky130_fd_sc_hd__o211a_2 _32810_ (.A1(_10756_),
    .A2(_10775_),
    .B1(_10772_),
    .C1(_10759_),
    .X(_10776_));
 sky130_fd_sc_hd__o22ai_2 _32811_ (.A1(_10579_),
    .A2(_10580_),
    .B1(_10773_),
    .B2(_10776_),
    .Y(_10777_));
 sky130_fd_sc_hd__a21oi_2 _32812_ (.A1(_10413_),
    .A2(_10366_),
    .B1(_10577_),
    .Y(_10778_));
 sky130_fd_sc_hd__a21oi_2 _32813_ (.A1(_10569_),
    .A2(_10575_),
    .B1(_10778_),
    .Y(_10779_));
 sky130_fd_sc_hd__inv_2 _32814_ (.A(_10366_),
    .Y(_10780_));
 sky130_fd_sc_hd__nor2_2 _32815_ (.A(_10413_),
    .B(_10577_),
    .Y(_10781_));
 sky130_fd_sc_hd__o211a_2 _32816_ (.A1(_10780_),
    .A2(_10781_),
    .B1(_10575_),
    .C1(_10568_),
    .X(_10782_));
 sky130_fd_sc_hd__nand3_2 _32817_ (.A(_10759_),
    .B(_10772_),
    .C(_10766_),
    .Y(_10783_));
 sky130_fd_sc_hd__a22oi_2 _32818_ (.A1(_10762_),
    .A2(_10763_),
    .B1(_10765_),
    .B2(_10774_),
    .Y(_10784_));
 sky130_fd_sc_hd__nor2_2 _32819_ (.A(_10756_),
    .B(_10775_),
    .Y(_10785_));
 sky130_fd_sc_hd__o21bai_2 _32820_ (.A1(_10784_),
    .A2(_10785_),
    .B1_N(_10772_),
    .Y(_10786_));
 sky130_fd_sc_hd__o211ai_2 _32821_ (.A1(_10779_),
    .A2(_10782_),
    .B1(_10783_),
    .C1(_10786_),
    .Y(_10787_));
 sky130_fd_sc_hd__inv_2 _32822_ (.A(_10313_),
    .Y(_10788_));
 sky130_fd_sc_hd__nand2_2 _32823_ (.A(_10319_),
    .B(_10317_),
    .Y(_10789_));
 sky130_fd_sc_hd__o22ai_2 _32824_ (.A1(_10788_),
    .A2(_10789_),
    .B1(_10320_),
    .B2(_10423_),
    .Y(_10790_));
 sky130_fd_sc_hd__a21oi_2 _32825_ (.A1(_10777_),
    .A2(_10787_),
    .B1(_10790_),
    .Y(_10791_));
 sky130_fd_sc_hd__a22oi_2 _32826_ (.A1(_10323_),
    .A2(_10322_),
    .B1(_10429_),
    .B2(_10431_),
    .Y(_10792_));
 sky130_fd_sc_hd__o211a_2 _32827_ (.A1(_10324_),
    .A2(_10792_),
    .B1(_10787_),
    .C1(_10777_),
    .X(_10793_));
 sky130_fd_sc_hd__o22ai_2 _32828_ (.A1(_10476_),
    .A2(_10477_),
    .B1(_10791_),
    .B2(_10793_),
    .Y(_10794_));
 sky130_fd_sc_hd__a21oi_2 _32829_ (.A1(_10433_),
    .A2(_10434_),
    .B1(_10432_),
    .Y(_10795_));
 sky130_fd_sc_hd__nand2_2 _32830_ (.A(_10427_),
    .B(_10435_),
    .Y(_10796_));
 sky130_fd_sc_hd__o2bb2ai_2 _32831_ (.A1_N(_10441_),
    .A2_N(_10448_),
    .B1(_10795_),
    .B2(_10796_),
    .Y(_10797_));
 sky130_fd_sc_hd__a21o_2 _32832_ (.A1(_10777_),
    .A2(_10787_),
    .B1(_10790_),
    .X(_10798_));
 sky130_fd_sc_hd__nand3_2 _32833_ (.A(_10790_),
    .B(_10787_),
    .C(_10777_),
    .Y(_10799_));
 sky130_fd_sc_hd__nor2_2 _32834_ (.A(_10476_),
    .B(_10477_),
    .Y(_10800_));
 sky130_fd_sc_hd__nand3_2 _32835_ (.A(_10798_),
    .B(_10799_),
    .C(_10800_),
    .Y(_10801_));
 sky130_fd_sc_hd__nand3_2 _32836_ (.A(_10794_),
    .B(_10797_),
    .C(_10801_),
    .Y(_10802_));
 sky130_fd_sc_hd__o21ai_2 _32837_ (.A1(_10791_),
    .A2(_10793_),
    .B1(_10800_),
    .Y(_10803_));
 sky130_fd_sc_hd__a21boi_2 _32838_ (.A1(_10448_),
    .A2(_10441_),
    .B1_N(_10436_),
    .Y(_10804_));
 sky130_fd_sc_hd__o211ai_2 _32839_ (.A1(_10476_),
    .A2(_10477_),
    .B1(_10799_),
    .C1(_10798_),
    .Y(_10805_));
 sky130_fd_sc_hd__nand3_2 _32840_ (.A(_10803_),
    .B(_10804_),
    .C(_10805_),
    .Y(_10806_));
 sky130_fd_sc_hd__o2bb2ai_2 _32841_ (.A1_N(_10802_),
    .A2_N(_10806_),
    .B1(_10442_),
    .B2(_10443_),
    .Y(_10807_));
 sky130_fd_sc_hd__nand3_2 _32842_ (.A(_10806_),
    .B(_10802_),
    .C(_10444_),
    .Y(_10808_));
 sky130_fd_sc_hd__nand2_2 _32843_ (.A(_10461_),
    .B(_10450_),
    .Y(_10809_));
 sky130_fd_sc_hd__a21o_2 _32844_ (.A1(_10807_),
    .A2(_10808_),
    .B1(_10809_),
    .X(_10810_));
 sky130_fd_sc_hd__nand3_2 _32845_ (.A(_10807_),
    .B(_10809_),
    .C(_10808_),
    .Y(_10811_));
 sky130_fd_sc_hd__nand2_2 _32846_ (.A(_10810_),
    .B(_10811_),
    .Y(_10812_));
 sky130_fd_sc_hd__a21bo_2 _32847_ (.A1(_10472_),
    .A2(_10464_),
    .B1_N(_10812_),
    .X(_10813_));
 sky130_fd_sc_hd__nand3b_2 _32848_ (.A_N(_10812_),
    .B(_10472_),
    .C(_10464_),
    .Y(_10814_));
 sky130_fd_sc_hd__nand2_2 _32849_ (.A(_10813_),
    .B(_10814_),
    .Y(_02650_));
 sky130_fd_sc_hd__a21bo_2 _32850_ (.A1(_10444_),
    .A2(_10806_),
    .B1_N(_10802_),
    .X(_10815_));
 sky130_fd_sc_hd__nand2_2 _32851_ (.A(_19311_),
    .B(_08393_),
    .Y(_10816_));
 sky130_fd_sc_hd__buf_1 _32852_ (.A(\pcpi_mul.rs2[32] ),
    .X(_10817_));
 sky130_fd_sc_hd__buf_1 _32853_ (.A(_10817_),
    .X(_10818_));
 sky130_fd_sc_hd__nand3_2 _32854_ (.A(_10818_),
    .B(_19307_),
    .C(_07904_),
    .Y(_10819_));
 sky130_fd_sc_hd__nor2_2 _32855_ (.A(_05805_),
    .B(_10819_),
    .Y(_10820_));
 sky130_fd_sc_hd__nor2_2 _32856_ (.A(_10816_),
    .B(_10820_),
    .Y(_10821_));
 sky130_fd_sc_hd__buf_1 _32857_ (.A(\pcpi_mul.rs2[31] ),
    .X(_10822_));
 sky130_fd_sc_hd__buf_1 _32858_ (.A(_10822_),
    .X(_10823_));
 sky130_fd_sc_hd__buf_1 _32859_ (.A(_10817_),
    .X(_10824_));
 sky130_fd_sc_hd__a22o_2 _32860_ (.A1(_10823_),
    .A2(_05804_),
    .B1(_04838_),
    .B2(_10824_),
    .X(_10825_));
 sky130_fd_sc_hd__nand2_2 _32861_ (.A(_19308_),
    .B(_06598_),
    .Y(_10826_));
 sky130_fd_sc_hd__buf_1 _32862_ (.A(_19312_),
    .X(_10827_));
 sky130_fd_sc_hd__nand3b_2 _32863_ (.A_N(_10826_),
    .B(_10827_),
    .C(_19637_),
    .Y(_10828_));
 sky130_fd_sc_hd__a21o_2 _32864_ (.A1(_10821_),
    .A2(_10825_),
    .B1(_10828_),
    .X(_10829_));
 sky130_fd_sc_hd__buf_1 _32865_ (.A(_18181_),
    .X(_10830_));
 sky130_fd_sc_hd__inv_2 _32866_ (.A(\pcpi_mul.rs2[31] ),
    .Y(_10831_));
 sky130_fd_sc_hd__buf_1 _32867_ (.A(_10831_),
    .X(_10832_));
 sky130_fd_sc_hd__o22a_2 _32868_ (.A1(_06598_),
    .A2(_10830_),
    .B1(_10832_),
    .B2(_05106_),
    .X(_10833_));
 sky130_fd_sc_hd__o21bai_2 _32869_ (.A1(_10820_),
    .A2(_10833_),
    .B1_N(_10816_),
    .Y(_10834_));
 sky130_fd_sc_hd__nand3b_2 _32870_ (.A_N(_10820_),
    .B(_10825_),
    .C(_10816_),
    .Y(_10835_));
 sky130_fd_sc_hd__nand3_2 _32871_ (.A(_10834_),
    .B(_10828_),
    .C(_10835_),
    .Y(_10836_));
 sky130_fd_sc_hd__nand2_2 _32872_ (.A(_19323_),
    .B(_05765_),
    .Y(_10837_));
 sky130_fd_sc_hd__inv_2 _32873_ (.A(_10837_),
    .Y(_10838_));
 sky130_fd_sc_hd__nand2_2 _32874_ (.A(_09841_),
    .B(_06792_),
    .Y(_10839_));
 sky130_fd_sc_hd__nand2_2 _32875_ (.A(_19319_),
    .B(_05206_),
    .Y(_10840_));
 sky130_fd_sc_hd__nor2_2 _32876_ (.A(_10839_),
    .B(_10840_),
    .Y(_10841_));
 sky130_fd_sc_hd__nand2_2 _32877_ (.A(_10839_),
    .B(_10840_),
    .Y(_10842_));
 sky130_fd_sc_hd__inv_2 _32878_ (.A(_10842_),
    .Y(_10843_));
 sky130_fd_sc_hd__nor2_2 _32879_ (.A(_10841_),
    .B(_10843_),
    .Y(_10844_));
 sky130_fd_sc_hd__nor2_2 _32880_ (.A(_10838_),
    .B(_10844_),
    .Y(_10845_));
 sky130_fd_sc_hd__and2_2 _32881_ (.A(_10844_),
    .B(_10838_),
    .X(_10846_));
 sky130_fd_sc_hd__o2bb2ai_2 _32882_ (.A1_N(_10829_),
    .A2_N(_10836_),
    .B1(_10845_),
    .B2(_10846_),
    .Y(_10847_));
 sky130_fd_sc_hd__inv_2 _32883_ (.A(_10717_),
    .Y(_10848_));
 sky130_fd_sc_hd__o21ai_2 _32884_ (.A1(_10841_),
    .A2(_10843_),
    .B1(_10838_),
    .Y(_10849_));
 sky130_fd_sc_hd__nand3b_2 _32885_ (.A_N(_10841_),
    .B(_10837_),
    .C(_10842_),
    .Y(_10850_));
 sky130_fd_sc_hd__nand2_2 _32886_ (.A(_10849_),
    .B(_10850_),
    .Y(_10851_));
 sky130_fd_sc_hd__nand3_2 _32887_ (.A(_10836_),
    .B(_10851_),
    .C(_10829_),
    .Y(_10852_));
 sky130_fd_sc_hd__nand3_2 _32888_ (.A(_10847_),
    .B(_10848_),
    .C(_10852_),
    .Y(_10853_));
 sky130_fd_sc_hd__nand2_2 _32889_ (.A(_10836_),
    .B(_10829_),
    .Y(_10854_));
 sky130_fd_sc_hd__nand2_2 _32890_ (.A(_10854_),
    .B(_10851_),
    .Y(_10855_));
 sky130_fd_sc_hd__nand3b_2 _32891_ (.A_N(_10851_),
    .B(_10836_),
    .C(_10829_),
    .Y(_10856_));
 sky130_fd_sc_hd__nand3_2 _32892_ (.A(_10855_),
    .B(_10717_),
    .C(_10856_),
    .Y(_10857_));
 sky130_fd_sc_hd__a21oi_2 _32893_ (.A1(_10707_),
    .A2(_10711_),
    .B1(_10710_),
    .Y(_10858_));
 sky130_fd_sc_hd__nand2_2 _32894_ (.A(_09826_),
    .B(_05422_),
    .Y(_10859_));
 sky130_fd_sc_hd__nand2_2 _32895_ (.A(_09827_),
    .B(_05426_),
    .Y(_10860_));
 sky130_fd_sc_hd__nor2_2 _32896_ (.A(_10859_),
    .B(_10860_),
    .Y(_10861_));
 sky130_fd_sc_hd__buf_1 _32897_ (.A(\pcpi_mul.rs2[24] ),
    .X(_10862_));
 sky130_fd_sc_hd__nand2_2 _32898_ (.A(_10862_),
    .B(_19616_),
    .Y(_10863_));
 sky130_fd_sc_hd__inv_2 _32899_ (.A(_10863_),
    .Y(_10864_));
 sky130_fd_sc_hd__nand2_2 _32900_ (.A(_10859_),
    .B(_10860_),
    .Y(_10865_));
 sky130_fd_sc_hd__nand3b_2 _32901_ (.A_N(_10861_),
    .B(_10864_),
    .C(_10865_),
    .Y(_10866_));
 sky130_fd_sc_hd__buf_1 _32902_ (.A(_09120_),
    .X(_10867_));
 sky130_fd_sc_hd__a21o_2 _32903_ (.A1(_10867_),
    .A2(_05713_),
    .B1(_10859_),
    .X(_10868_));
 sky130_fd_sc_hd__a21o_2 _32904_ (.A1(_19328_),
    .A2(_05343_),
    .B1(_10860_),
    .X(_10869_));
 sky130_fd_sc_hd__nand3_2 _32905_ (.A(_10868_),
    .B(_10869_),
    .C(_10863_),
    .Y(_10870_));
 sky130_fd_sc_hd__nand2_2 _32906_ (.A(_10866_),
    .B(_10870_),
    .Y(_10871_));
 sky130_fd_sc_hd__nor2_2 _32907_ (.A(_10858_),
    .B(_10871_),
    .Y(_10872_));
 sky130_fd_sc_hd__nand2_2 _32908_ (.A(_10871_),
    .B(_10858_),
    .Y(_10873_));
 sky130_fd_sc_hd__nor2_2 _32909_ (.A(_10727_),
    .B(_10731_),
    .Y(_10874_));
 sky130_fd_sc_hd__nor2_2 _32910_ (.A(_10725_),
    .B(_10874_),
    .Y(_10875_));
 sky130_fd_sc_hd__inv_2 _32911_ (.A(_10875_),
    .Y(_10876_));
 sky130_fd_sc_hd__nand2_2 _32912_ (.A(_10873_),
    .B(_10876_),
    .Y(_10877_));
 sky130_fd_sc_hd__nor2_2 _32913_ (.A(_10872_),
    .B(_10877_),
    .Y(_10878_));
 sky130_fd_sc_hd__a21o_2 _32914_ (.A1(_10707_),
    .A2(_10711_),
    .B1(_10710_),
    .X(_10879_));
 sky130_fd_sc_hd__nand3_2 _32915_ (.A(_10879_),
    .B(_10866_),
    .C(_10870_),
    .Y(_10880_));
 sky130_fd_sc_hd__a21oi_2 _32916_ (.A1(_10873_),
    .A2(_10880_),
    .B1(_10876_),
    .Y(_10881_));
 sky130_fd_sc_hd__o2bb2ai_2 _32917_ (.A1_N(_10853_),
    .A2_N(_10857_),
    .B1(_10878_),
    .B2(_10881_),
    .Y(_10882_));
 sky130_fd_sc_hd__a21oi_2 _32918_ (.A1(_10866_),
    .A2(_10870_),
    .B1(_10879_),
    .Y(_10883_));
 sky130_fd_sc_hd__nor2_2 _32919_ (.A(_10875_),
    .B(_10883_),
    .Y(_10884_));
 sky130_fd_sc_hd__a21oi_2 _32920_ (.A1(_10880_),
    .A2(_10884_),
    .B1(_10881_),
    .Y(_10885_));
 sky130_fd_sc_hd__nand3_2 _32921_ (.A(_10885_),
    .B(_10857_),
    .C(_10853_),
    .Y(_10886_));
 sky130_fd_sc_hd__nand2_2 _32922_ (.A(_10745_),
    .B(_10723_),
    .Y(_10887_));
 sky130_fd_sc_hd__nand3_2 _32923_ (.A(_10882_),
    .B(_10886_),
    .C(_10887_),
    .Y(_10888_));
 sky130_fd_sc_hd__nand2_2 _32924_ (.A(_10857_),
    .B(_10853_),
    .Y(_10889_));
 sky130_fd_sc_hd__nand2_2 _32925_ (.A(_10889_),
    .B(_10885_),
    .Y(_10890_));
 sky130_fd_sc_hd__and2_2 _32926_ (.A(_10745_),
    .B(_10723_),
    .X(_10891_));
 sky130_fd_sc_hd__o211ai_2 _32927_ (.A1(_10881_),
    .A2(_10878_),
    .B1(_10857_),
    .C1(_10853_),
    .Y(_10892_));
 sky130_fd_sc_hd__nand3_2 _32928_ (.A(_10890_),
    .B(_10891_),
    .C(_10892_),
    .Y(_10893_));
 sky130_fd_sc_hd__a21oi_2 _32929_ (.A1(_10664_),
    .A2(_10661_),
    .B1(_10659_),
    .Y(_10894_));
 sky130_fd_sc_hd__nand2_2 _32930_ (.A(_19336_),
    .B(_05614_),
    .Y(_10895_));
 sky130_fd_sc_hd__nand2_2 _32931_ (.A(_19339_),
    .B(_06497_),
    .Y(_10896_));
 sky130_fd_sc_hd__nor2_2 _32932_ (.A(_10895_),
    .B(_10896_),
    .Y(_10897_));
 sky130_fd_sc_hd__nand2_2 _32933_ (.A(_10895_),
    .B(_10896_),
    .Y(_10898_));
 sky130_fd_sc_hd__nand2_2 _32934_ (.A(_19342_),
    .B(_05717_),
    .Y(_10899_));
 sky130_fd_sc_hd__inv_2 _32935_ (.A(_10899_),
    .Y(_10900_));
 sky130_fd_sc_hd__nand3b_2 _32936_ (.A_N(_10897_),
    .B(_10898_),
    .C(_10900_),
    .Y(_10901_));
 sky130_fd_sc_hd__and2_2 _32937_ (.A(_10895_),
    .B(_10896_),
    .X(_10902_));
 sky130_fd_sc_hd__o21ai_2 _32938_ (.A1(_10897_),
    .A2(_10902_),
    .B1(_10899_),
    .Y(_10903_));
 sky130_fd_sc_hd__nand3b_2 _32939_ (.A_N(_10894_),
    .B(_10901_),
    .C(_10903_),
    .Y(_10904_));
 sky130_fd_sc_hd__o21ai_2 _32940_ (.A1(_10897_),
    .A2(_10902_),
    .B1(_10900_),
    .Y(_10905_));
 sky130_fd_sc_hd__nand3b_2 _32941_ (.A_N(_10897_),
    .B(_10898_),
    .C(_10899_),
    .Y(_10906_));
 sky130_fd_sc_hd__nand3_2 _32942_ (.A(_10905_),
    .B(_10906_),
    .C(_10894_),
    .Y(_10907_));
 sky130_fd_sc_hd__nand2_2 _32943_ (.A(_07480_),
    .B(_07109_),
    .Y(_10908_));
 sky130_fd_sc_hd__nand2_2 _32944_ (.A(_07906_),
    .B(_08218_),
    .Y(_10909_));
 sky130_fd_sc_hd__nor2_2 _32945_ (.A(_10908_),
    .B(_10909_),
    .Y(_10910_));
 sky130_fd_sc_hd__nand2_2 _32946_ (.A(_10908_),
    .B(_10909_),
    .Y(_10911_));
 sky130_fd_sc_hd__inv_2 _32947_ (.A(_10911_),
    .Y(_10912_));
 sky130_fd_sc_hd__nand2_2 _32948_ (.A(_08407_),
    .B(_08761_),
    .Y(_10913_));
 sky130_fd_sc_hd__inv_2 _32949_ (.A(_10913_),
    .Y(_10914_));
 sky130_fd_sc_hd__o21ai_2 _32950_ (.A1(_10910_),
    .A2(_10912_),
    .B1(_10914_),
    .Y(_10915_));
 sky130_fd_sc_hd__nand3b_2 _32951_ (.A_N(_10910_),
    .B(_10913_),
    .C(_10911_),
    .Y(_10916_));
 sky130_fd_sc_hd__nand2_2 _32952_ (.A(_10915_),
    .B(_10916_),
    .Y(_10917_));
 sky130_fd_sc_hd__a21oi_2 _32953_ (.A1(_10904_),
    .A2(_10907_),
    .B1(_10917_),
    .Y(_10918_));
 sky130_fd_sc_hd__nor3_2 _32954_ (.A(_10910_),
    .B(_10914_),
    .C(_10912_),
    .Y(_10919_));
 sky130_fd_sc_hd__o21a_2 _32955_ (.A1(_10910_),
    .A2(_10912_),
    .B1(_10914_),
    .X(_10920_));
 sky130_fd_sc_hd__o211a_2 _32956_ (.A1(_10919_),
    .A2(_10920_),
    .B1(_10907_),
    .C1(_10904_),
    .X(_10921_));
 sky130_fd_sc_hd__nand2_2 _32957_ (.A(_10741_),
    .B(_10733_),
    .Y(_10922_));
 sky130_fd_sc_hd__o21bai_2 _32958_ (.A1(_10918_),
    .A2(_10921_),
    .B1_N(_10922_),
    .Y(_10923_));
 sky130_fd_sc_hd__a21o_2 _32959_ (.A1(_10904_),
    .A2(_10907_),
    .B1(_10917_),
    .X(_10924_));
 sky130_fd_sc_hd__nand3_2 _32960_ (.A(_10904_),
    .B(_10917_),
    .C(_10907_),
    .Y(_10925_));
 sky130_fd_sc_hd__nand3_2 _32961_ (.A(_10924_),
    .B(_10922_),
    .C(_10925_),
    .Y(_10926_));
 sky130_fd_sc_hd__nand2_2 _32962_ (.A(_10684_),
    .B(_10666_),
    .Y(_10927_));
 sky130_fd_sc_hd__nand2_2 _32963_ (.A(_10927_),
    .B(_10670_),
    .Y(_10928_));
 sky130_fd_sc_hd__a21oi_2 _32964_ (.A1(_10923_),
    .A2(_10926_),
    .B1(_10928_),
    .Y(_10929_));
 sky130_fd_sc_hd__nand3_2 _32965_ (.A(_10923_),
    .B(_10926_),
    .C(_10928_),
    .Y(_10930_));
 sky130_fd_sc_hd__inv_2 _32966_ (.A(_10930_),
    .Y(_10931_));
 sky130_fd_sc_hd__o2bb2ai_2 _32967_ (.A1_N(_10888_),
    .A2_N(_10893_),
    .B1(_10929_),
    .B2(_10931_),
    .Y(_10932_));
 sky130_fd_sc_hd__inv_2 _32968_ (.A(_10928_),
    .Y(_10933_));
 sky130_fd_sc_hd__a21oi_2 _32969_ (.A1(_10924_),
    .A2(_10925_),
    .B1(_10922_),
    .Y(_10934_));
 sky130_fd_sc_hd__nor2_2 _32970_ (.A(_10933_),
    .B(_10934_),
    .Y(_10935_));
 sky130_fd_sc_hd__a21oi_2 _32971_ (.A1(_10935_),
    .A2(_10926_),
    .B1(_10929_),
    .Y(_10936_));
 sky130_fd_sc_hd__nand3_2 _32972_ (.A(_10936_),
    .B(_10888_),
    .C(_10893_),
    .Y(_10937_));
 sky130_fd_sc_hd__nand2_2 _32973_ (.A(_10753_),
    .B(_10751_),
    .Y(_10938_));
 sky130_fd_sc_hd__a21o_2 _32974_ (.A1(_10932_),
    .A2(_10937_),
    .B1(_10938_),
    .X(_10939_));
 sky130_fd_sc_hd__a21oi_2 _32975_ (.A1(_10678_),
    .A2(_10679_),
    .B1(_10673_),
    .Y(_10940_));
 sky130_fd_sc_hd__nand3_2 _32976_ (.A(_06822_),
    .B(_06824_),
    .C(_06748_),
    .Y(_10941_));
 sky130_fd_sc_hd__a22o_2 _32977_ (.A1(_09018_),
    .A2(_07798_),
    .B1(_09019_),
    .B2(_19590_),
    .X(_10942_));
 sky130_fd_sc_hd__o21ai_2 _32978_ (.A1(_10268_),
    .A2(_10941_),
    .B1(_10942_),
    .Y(_10943_));
 sky130_fd_sc_hd__nand2_2 _32979_ (.A(_09386_),
    .B(_08447_),
    .Y(_10944_));
 sky130_fd_sc_hd__nand2_2 _32980_ (.A(_10943_),
    .B(_10944_),
    .Y(_10945_));
 sky130_fd_sc_hd__nor2_2 _32981_ (.A(_08053_),
    .B(_10941_),
    .Y(_10946_));
 sky130_fd_sc_hd__inv_2 _32982_ (.A(_10944_),
    .Y(_10947_));
 sky130_fd_sc_hd__nand3b_2 _32983_ (.A_N(_10946_),
    .B(_10942_),
    .C(_10947_),
    .Y(_10948_));
 sky130_fd_sc_hd__nand3b_2 _32984_ (.A_N(_10940_),
    .B(_10945_),
    .C(_10948_),
    .Y(_10949_));
 sky130_fd_sc_hd__nand2_2 _32985_ (.A(_10943_),
    .B(_10947_),
    .Y(_10950_));
 sky130_fd_sc_hd__nand3b_2 _32986_ (.A_N(_10946_),
    .B(_10942_),
    .C(_10944_),
    .Y(_10951_));
 sky130_fd_sc_hd__nand3_2 _32987_ (.A(_10950_),
    .B(_10951_),
    .C(_10940_),
    .Y(_10952_));
 sky130_fd_sc_hd__or2_2 _32988_ (.A(_10587_),
    .B(_10584_),
    .X(_10953_));
 sky130_fd_sc_hd__a21o_2 _32989_ (.A1(_10949_),
    .A2(_10952_),
    .B1(_10953_),
    .X(_10954_));
 sky130_fd_sc_hd__nand3_2 _32990_ (.A(_10949_),
    .B(_10952_),
    .C(_10953_),
    .Y(_10955_));
 sky130_fd_sc_hd__nand2_2 _32991_ (.A(_10599_),
    .B(_10589_),
    .Y(_10956_));
 sky130_fd_sc_hd__a21oi_2 _32992_ (.A1(_10954_),
    .A2(_10955_),
    .B1(_10956_),
    .Y(_10957_));
 sky130_fd_sc_hd__a21oi_2 _32993_ (.A1(_10950_),
    .A2(_10951_),
    .B1(_10940_),
    .Y(_10958_));
 sky130_fd_sc_hd__nand2_2 _32994_ (.A(_10952_),
    .B(_10953_),
    .Y(_10959_));
 sky130_fd_sc_hd__o211a_2 _32995_ (.A1(_10958_),
    .A2(_10959_),
    .B1(_10956_),
    .C1(_10954_),
    .X(_10960_));
 sky130_fd_sc_hd__nand2_2 _32996_ (.A(_09051_),
    .B(_09250_),
    .Y(_10961_));
 sky130_fd_sc_hd__nand2_2 _32997_ (.A(_06605_),
    .B(_08103_),
    .Y(_10962_));
 sky130_fd_sc_hd__nor2_2 _32998_ (.A(_10961_),
    .B(_10962_),
    .Y(_10963_));
 sky130_fd_sc_hd__nand2_2 _32999_ (.A(_10961_),
    .B(_10962_),
    .Y(_10964_));
 sky130_fd_sc_hd__inv_2 _33000_ (.A(_10964_),
    .Y(_10965_));
 sky130_fd_sc_hd__buf_1 _33001_ (.A(_09199_),
    .X(_10966_));
 sky130_fd_sc_hd__nand2_2 _33002_ (.A(_06020_),
    .B(_10966_),
    .Y(_10967_));
 sky130_fd_sc_hd__o21bai_2 _33003_ (.A1(_10963_),
    .A2(_10965_),
    .B1_N(_10967_),
    .Y(_10968_));
 sky130_fd_sc_hd__nand3b_2 _33004_ (.A_N(_10963_),
    .B(_10967_),
    .C(_10964_),
    .Y(_10969_));
 sky130_fd_sc_hd__nand2_2 _33005_ (.A(_10968_),
    .B(_10969_),
    .Y(_10970_));
 sky130_fd_sc_hd__nand3_2 _33006_ (.A(_06271_),
    .B(_08320_),
    .C(_08950_),
    .Y(_10971_));
 sky130_fd_sc_hd__nor2_2 _33007_ (.A(_08947_),
    .B(_10971_),
    .Y(_10972_));
 sky130_fd_sc_hd__a22o_2 _33008_ (.A1(_19364_),
    .A2(_08959_),
    .B1(_06273_),
    .B2(_09933_),
    .X(_10973_));
 sky130_fd_sc_hd__nand2_2 _33009_ (.A(_06628_),
    .B(_07590_),
    .Y(_10974_));
 sky130_fd_sc_hd__inv_2 _33010_ (.A(_10974_),
    .Y(_10975_));
 sky130_fd_sc_hd__nand2_2 _33011_ (.A(_10973_),
    .B(_10975_),
    .Y(_10976_));
 sky130_fd_sc_hd__a21o_2 _33012_ (.A1(_10610_),
    .A2(_10612_),
    .B1(_10607_),
    .X(_10977_));
 sky130_fd_sc_hd__o21ai_2 _33013_ (.A1(_08957_),
    .A2(_10971_),
    .B1(_10973_),
    .Y(_10978_));
 sky130_fd_sc_hd__nand2_2 _33014_ (.A(_10978_),
    .B(_10974_),
    .Y(_10979_));
 sky130_fd_sc_hd__o211ai_2 _33015_ (.A1(_10972_),
    .A2(_10976_),
    .B1(_10977_),
    .C1(_10979_),
    .Y(_10980_));
 sky130_fd_sc_hd__nand2_2 _33016_ (.A(_10978_),
    .B(_10975_),
    .Y(_10981_));
 sky130_fd_sc_hd__nand3b_2 _33017_ (.A_N(_10972_),
    .B(_10973_),
    .C(_10974_),
    .Y(_10982_));
 sky130_fd_sc_hd__a21oi_2 _33018_ (.A1(_10610_),
    .A2(_10612_),
    .B1(_10607_),
    .Y(_10983_));
 sky130_fd_sc_hd__nand3_2 _33019_ (.A(_10981_),
    .B(_10982_),
    .C(_10983_),
    .Y(_10984_));
 sky130_fd_sc_hd__nand2_2 _33020_ (.A(_10980_),
    .B(_10984_),
    .Y(_10985_));
 sky130_fd_sc_hd__xor2_2 _33021_ (.A(_10970_),
    .B(_10985_),
    .X(_10986_));
 sky130_fd_sc_hd__o21ai_2 _33022_ (.A1(_10957_),
    .A2(_10960_),
    .B1(_10986_),
    .Y(_10987_));
 sky130_fd_sc_hd__nand2_2 _33023_ (.A(_10750_),
    .B(_10697_),
    .Y(_10988_));
 sky130_fd_sc_hd__a21o_2 _33024_ (.A1(_10954_),
    .A2(_10955_),
    .B1(_10956_),
    .X(_10989_));
 sky130_fd_sc_hd__xnor2_2 _33025_ (.A(_10970_),
    .B(_10985_),
    .Y(_10990_));
 sky130_fd_sc_hd__nand3_2 _33026_ (.A(_10956_),
    .B(_10954_),
    .C(_10955_),
    .Y(_10991_));
 sky130_fd_sc_hd__nand3_2 _33027_ (.A(_10989_),
    .B(_10990_),
    .C(_10991_),
    .Y(_10992_));
 sky130_fd_sc_hd__nand3_2 _33028_ (.A(_10987_),
    .B(_10988_),
    .C(_10992_),
    .Y(_10993_));
 sky130_fd_sc_hd__o21ai_2 _33029_ (.A1(_10957_),
    .A2(_10960_),
    .B1(_10990_),
    .Y(_10994_));
 sky130_fd_sc_hd__nand3_2 _33030_ (.A(_10989_),
    .B(_10986_),
    .C(_10991_),
    .Y(_10995_));
 sky130_fd_sc_hd__a21oi_2 _33031_ (.A1(_10696_),
    .A2(_10692_),
    .B1(_10690_),
    .Y(_10996_));
 sky130_fd_sc_hd__a21oi_2 _33032_ (.A1(_10639_),
    .A2(_10632_),
    .B1(_10604_),
    .Y(_10997_));
 sky130_fd_sc_hd__a31oi_2 _33033_ (.A1(_10994_),
    .A2(_10995_),
    .A3(_10996_),
    .B1(_10997_),
    .Y(_10998_));
 sky130_fd_sc_hd__nand3_2 _33034_ (.A(_10994_),
    .B(_10996_),
    .C(_10995_),
    .Y(_10999_));
 sky130_fd_sc_hd__inv_2 _33035_ (.A(_10997_),
    .Y(_11000_));
 sky130_fd_sc_hd__a21oi_2 _33036_ (.A1(_10999_),
    .A2(_10993_),
    .B1(_11000_),
    .Y(_11001_));
 sky130_fd_sc_hd__a21oi_2 _33037_ (.A1(_10993_),
    .A2(_10998_),
    .B1(_11001_),
    .Y(_11002_));
 sky130_fd_sc_hd__nand3_2 _33038_ (.A(_10932_),
    .B(_10938_),
    .C(_10937_),
    .Y(_11003_));
 sky130_fd_sc_hd__nand3_2 _33039_ (.A(_10939_),
    .B(_11002_),
    .C(_11003_),
    .Y(_11004_));
 sky130_fd_sc_hd__a21oi_2 _33040_ (.A1(_10932_),
    .A2(_10937_),
    .B1(_10938_),
    .Y(_11005_));
 sky130_fd_sc_hd__o211a_2 _33041_ (.A1(_10748_),
    .A2(_10764_),
    .B1(_10937_),
    .C1(_10932_),
    .X(_11006_));
 sky130_fd_sc_hd__a21o_2 _33042_ (.A1(_10993_),
    .A2(_10999_),
    .B1(_11000_),
    .X(_11007_));
 sky130_fd_sc_hd__nand2_2 _33043_ (.A(_10998_),
    .B(_10993_),
    .Y(_11008_));
 sky130_fd_sc_hd__nand2_2 _33044_ (.A(_11007_),
    .B(_11008_),
    .Y(_11009_));
 sky130_fd_sc_hd__o21ai_2 _33045_ (.A1(_11005_),
    .A2(_11006_),
    .B1(_11009_),
    .Y(_11010_));
 sky130_fd_sc_hd__o211ai_2 _33046_ (.A1(_10758_),
    .A2(_10785_),
    .B1(_11004_),
    .C1(_11010_),
    .Y(_11011_));
 sky130_fd_sc_hd__o21ai_2 _33047_ (.A1(_11005_),
    .A2(_11006_),
    .B1(_11002_),
    .Y(_11012_));
 sky130_fd_sc_hd__o21a_2 _33048_ (.A1(_10756_),
    .A2(_10775_),
    .B1(_10774_),
    .X(_11013_));
 sky130_fd_sc_hd__nand3_2 _33049_ (.A(_10939_),
    .B(_11003_),
    .C(_11009_),
    .Y(_11014_));
 sky130_fd_sc_hd__nand3_2 _33050_ (.A(_11012_),
    .B(_11013_),
    .C(_11014_),
    .Y(_11015_));
 sky130_fd_sc_hd__nand2_2 _33051_ (.A(_11011_),
    .B(_11015_),
    .Y(_11016_));
 sky130_fd_sc_hd__a21oi_2 _33052_ (.A1(_10521_),
    .A2(_10517_),
    .B1(_10516_),
    .Y(_11017_));
 sky130_fd_sc_hd__nand2_2 _33053_ (.A(_06735_),
    .B(_09736_),
    .Y(_11018_));
 sky130_fd_sc_hd__nand2_2 _33054_ (.A(_05403_),
    .B(_09722_),
    .Y(_11019_));
 sky130_fd_sc_hd__nor2_2 _33055_ (.A(_11018_),
    .B(_11019_),
    .Y(_11020_));
 sky130_fd_sc_hd__inv_2 _33056_ (.A(_11020_),
    .Y(_11021_));
 sky130_fd_sc_hd__nand2_2 _33057_ (.A(_11018_),
    .B(_11019_),
    .Y(_11022_));
 sky130_fd_sc_hd__buf_1 _33058_ (.A(\pcpi_mul.rs1[32] ),
    .X(_11023_));
 sky130_fd_sc_hd__nand2_2 _33059_ (.A(_11023_),
    .B(_19403_),
    .Y(_11024_));
 sky130_fd_sc_hd__inv_2 _33060_ (.A(_11024_),
    .Y(_11025_));
 sky130_fd_sc_hd__buf_1 _33061_ (.A(_11025_),
    .X(_11026_));
 sky130_fd_sc_hd__nand3_2 _33062_ (.A(_11021_),
    .B(_11022_),
    .C(_11026_),
    .Y(_11027_));
 sky130_fd_sc_hd__and2_2 _33063_ (.A(_11018_),
    .B(_11019_),
    .X(_11028_));
 sky130_fd_sc_hd__buf_1 _33064_ (.A(_11024_),
    .X(_11029_));
 sky130_fd_sc_hd__buf_1 _33065_ (.A(_11029_),
    .X(_11030_));
 sky130_fd_sc_hd__o21ai_2 _33066_ (.A1(_11020_),
    .A2(_11028_),
    .B1(_11030_),
    .Y(_11031_));
 sky130_fd_sc_hd__nand3b_2 _33067_ (.A_N(_11017_),
    .B(_11027_),
    .C(_11031_),
    .Y(_11032_));
 sky130_fd_sc_hd__nand3_2 _33068_ (.A(_11021_),
    .B(_11022_),
    .C(_11030_),
    .Y(_11033_));
 sky130_fd_sc_hd__o21ai_2 _33069_ (.A1(_11020_),
    .A2(_11028_),
    .B1(_11026_),
    .Y(_11034_));
 sky130_fd_sc_hd__nand3_2 _33070_ (.A(_11033_),
    .B(_11034_),
    .C(_11017_),
    .Y(_11035_));
 sky130_fd_sc_hd__buf_1 _33071_ (.A(_10532_),
    .X(_11036_));
 sky130_fd_sc_hd__buf_1 _33072_ (.A(_19544_),
    .X(_11037_));
 sky130_fd_sc_hd__buf_1 _33073_ (.A(_11037_),
    .X(_11038_));
 sky130_fd_sc_hd__a22oi_2 _33074_ (.A1(_19399_),
    .A2(_11038_),
    .B1(_19402_),
    .B2(_19541_),
    .Y(_11039_));
 sky130_fd_sc_hd__and4_2 _33075_ (.A(_05141_),
    .B(_05144_),
    .C(_19541_),
    .D(_11038_),
    .X(_11040_));
 sky130_fd_sc_hd__nor2_2 _33076_ (.A(_11039_),
    .B(_11040_),
    .Y(_11041_));
 sky130_fd_sc_hd__o21ai_2 _33077_ (.A1(_05151_),
    .A2(_11036_),
    .B1(_11041_),
    .Y(_11042_));
 sky130_fd_sc_hd__nor2_2 _33078_ (.A(_05151_),
    .B(_11036_),
    .Y(_11043_));
 sky130_fd_sc_hd__o21ai_2 _33079_ (.A1(_11039_),
    .A2(_11040_),
    .B1(_11043_),
    .Y(_11044_));
 sky130_fd_sc_hd__nand2_2 _33080_ (.A(_11042_),
    .B(_11044_),
    .Y(_11045_));
 sky130_fd_sc_hd__a21o_2 _33081_ (.A1(_11032_),
    .A2(_11035_),
    .B1(_11045_),
    .X(_11046_));
 sky130_fd_sc_hd__nand3_2 _33082_ (.A(_11032_),
    .B(_11045_),
    .C(_11035_),
    .Y(_11047_));
 sky130_fd_sc_hd__a21oi_2 _33083_ (.A1(_10525_),
    .A2(_10522_),
    .B1(_10528_),
    .Y(_11048_));
 sky130_fd_sc_hd__o21ai_2 _33084_ (.A1(_11048_),
    .A2(_10550_),
    .B1(_10529_),
    .Y(_11049_));
 sky130_fd_sc_hd__a21o_2 _33085_ (.A1(_11046_),
    .A2(_11047_),
    .B1(_11049_),
    .X(_11050_));
 sky130_fd_sc_hd__nand3_2 _33086_ (.A(_11046_),
    .B(_11049_),
    .C(_11047_),
    .Y(_11051_));
 sky130_fd_sc_hd__nand2_2 _33087_ (.A(_10545_),
    .B(_10541_),
    .Y(_11052_));
 sky130_fd_sc_hd__a21oi_2 _33088_ (.A1(_11050_),
    .A2(_11051_),
    .B1(_11052_),
    .Y(_11053_));
 sky130_fd_sc_hd__and3_2 _33089_ (.A(_11050_),
    .B(_11052_),
    .C(_11051_),
    .X(_11054_));
 sky130_fd_sc_hd__nand3_2 _33090_ (.A(_08948_),
    .B(_09254_),
    .C(_10380_),
    .Y(_11055_));
 sky130_fd_sc_hd__a22o_2 _33091_ (.A1(_19381_),
    .A2(_08922_),
    .B1(_09254_),
    .B2(_19565_),
    .X(_11056_));
 sky130_fd_sc_hd__o21ai_2 _33092_ (.A1(_10485_),
    .A2(_11055_),
    .B1(_11056_),
    .Y(_11057_));
 sky130_fd_sc_hd__nand2_2 _33093_ (.A(_19386_),
    .B(_09220_),
    .Y(_11058_));
 sky130_fd_sc_hd__nand2_2 _33094_ (.A(_11057_),
    .B(_11058_),
    .Y(_11059_));
 sky130_fd_sc_hd__nor2_2 _33095_ (.A(_08487_),
    .B(_11055_),
    .Y(_11060_));
 sky130_fd_sc_hd__inv_2 _33096_ (.A(_11058_),
    .Y(_11061_));
 sky130_fd_sc_hd__nand3b_2 _33097_ (.A_N(_11060_),
    .B(_11056_),
    .C(_11061_),
    .Y(_11062_));
 sky130_fd_sc_hd__a21o_2 _33098_ (.A1(_10624_),
    .A2(_10621_),
    .B1(_10620_),
    .X(_11063_));
 sky130_fd_sc_hd__nand3_2 _33099_ (.A(_11059_),
    .B(_11062_),
    .C(_11063_),
    .Y(_11064_));
 sky130_fd_sc_hd__nand2_2 _33100_ (.A(_11057_),
    .B(_11061_),
    .Y(_11065_));
 sky130_fd_sc_hd__nand3b_2 _33101_ (.A_N(_11060_),
    .B(_11056_),
    .C(_11058_),
    .Y(_11066_));
 sky130_fd_sc_hd__a21oi_2 _33102_ (.A1(_10624_),
    .A2(_10621_),
    .B1(_10620_),
    .Y(_11067_));
 sky130_fd_sc_hd__nand3_2 _33103_ (.A(_11065_),
    .B(_11066_),
    .C(_11067_),
    .Y(_11068_));
 sky130_fd_sc_hd__nor2_2 _33104_ (.A(_10483_),
    .B(_10480_),
    .Y(_11069_));
 sky130_fd_sc_hd__nor2_2 _33105_ (.A(_10482_),
    .B(_11069_),
    .Y(_11070_));
 sky130_fd_sc_hd__inv_2 _33106_ (.A(_11070_),
    .Y(_11071_));
 sky130_fd_sc_hd__a21o_2 _33107_ (.A1(_11064_),
    .A2(_11068_),
    .B1(_11071_),
    .X(_11072_));
 sky130_fd_sc_hd__nand3_2 _33108_ (.A(_11071_),
    .B(_11064_),
    .C(_11068_),
    .Y(_11073_));
 sky130_fd_sc_hd__nand2_2 _33109_ (.A(_10636_),
    .B(_10630_),
    .Y(_11074_));
 sky130_fd_sc_hd__a21oi_2 _33110_ (.A1(_11072_),
    .A2(_11073_),
    .B1(_11074_),
    .Y(_11075_));
 sky130_fd_sc_hd__inv_2 _33111_ (.A(_11064_),
    .Y(_11076_));
 sky130_fd_sc_hd__nand2_2 _33112_ (.A(_11071_),
    .B(_11068_),
    .Y(_11077_));
 sky130_fd_sc_hd__o211a_2 _33113_ (.A1(_11076_),
    .A2(_11077_),
    .B1(_11074_),
    .C1(_11072_),
    .X(_11078_));
 sky130_fd_sc_hd__nand2_2 _33114_ (.A(_10501_),
    .B(_10490_),
    .Y(_11079_));
 sky130_fd_sc_hd__inv_2 _33115_ (.A(_11079_),
    .Y(_11080_));
 sky130_fd_sc_hd__o21ai_2 _33116_ (.A1(_11075_),
    .A2(_11078_),
    .B1(_11080_),
    .Y(_11081_));
 sky130_fd_sc_hd__a21o_2 _33117_ (.A1(_11072_),
    .A2(_11073_),
    .B1(_11074_),
    .X(_11082_));
 sky130_fd_sc_hd__nand3_2 _33118_ (.A(_11072_),
    .B(_11074_),
    .C(_11073_),
    .Y(_11083_));
 sky130_fd_sc_hd__nand3_2 _33119_ (.A(_11082_),
    .B(_11083_),
    .C(_11079_),
    .Y(_11084_));
 sky130_fd_sc_hd__nand2_2 _33120_ (.A(_10507_),
    .B(_10506_),
    .Y(_11085_));
 sky130_fd_sc_hd__a21oi_2 _33121_ (.A1(_11081_),
    .A2(_11084_),
    .B1(_11085_),
    .Y(_11086_));
 sky130_fd_sc_hd__nor2_2 _33122_ (.A(_10504_),
    .B(_10499_),
    .Y(_11087_));
 sky130_fd_sc_hd__o211a_2 _33123_ (.A1(_10502_),
    .A2(_11087_),
    .B1(_11084_),
    .C1(_11081_),
    .X(_11088_));
 sky130_fd_sc_hd__o22ai_2 _33124_ (.A1(_11053_),
    .A2(_11054_),
    .B1(_11086_),
    .B2(_11088_),
    .Y(_11089_));
 sky130_fd_sc_hd__nor2_2 _33125_ (.A(_11053_),
    .B(_11054_),
    .Y(_11090_));
 sky130_fd_sc_hd__a21o_2 _33126_ (.A1(_11081_),
    .A2(_11084_),
    .B1(_11085_),
    .X(_11091_));
 sky130_fd_sc_hd__nand3_2 _33127_ (.A(_11085_),
    .B(_11081_),
    .C(_11084_),
    .Y(_11092_));
 sky130_fd_sc_hd__nand3_2 _33128_ (.A(_11090_),
    .B(_11091_),
    .C(_11092_),
    .Y(_11093_));
 sky130_fd_sc_hd__nand2_2 _33129_ (.A(_10763_),
    .B(_10648_),
    .Y(_11094_));
 sky130_fd_sc_hd__a21oi_2 _33130_ (.A1(_11089_),
    .A2(_11093_),
    .B1(_11094_),
    .Y(_11095_));
 sky130_fd_sc_hd__and3_2 _33131_ (.A(_11089_),
    .B(_11093_),
    .C(_11094_),
    .X(_11096_));
 sky130_fd_sc_hd__nor2_2 _33132_ (.A(_10509_),
    .B(_10564_),
    .Y(_11097_));
 sky130_fd_sc_hd__nor2_2 _33133_ (.A(_10511_),
    .B(_11097_),
    .Y(_11098_));
 sky130_fd_sc_hd__o21ai_2 _33134_ (.A1(_11095_),
    .A2(_11096_),
    .B1(_11098_),
    .Y(_11099_));
 sky130_fd_sc_hd__a21o_2 _33135_ (.A1(_11089_),
    .A2(_11093_),
    .B1(_11094_),
    .X(_11100_));
 sky130_fd_sc_hd__inv_2 _33136_ (.A(_11098_),
    .Y(_11101_));
 sky130_fd_sc_hd__nand3_2 _33137_ (.A(_11089_),
    .B(_11093_),
    .C(_11094_),
    .Y(_11102_));
 sky130_fd_sc_hd__nand3_2 _33138_ (.A(_11100_),
    .B(_11101_),
    .C(_11102_),
    .Y(_11103_));
 sky130_fd_sc_hd__nand2_2 _33139_ (.A(_11099_),
    .B(_11103_),
    .Y(_11104_));
 sky130_fd_sc_hd__nand2_2 _33140_ (.A(_11016_),
    .B(_11104_),
    .Y(_11105_));
 sky130_fd_sc_hd__a21o_2 _33141_ (.A1(_10569_),
    .A2(_10576_),
    .B1(_10778_),
    .X(_11106_));
 sky130_fd_sc_hd__nand3_2 _33142_ (.A(_10569_),
    .B(_10576_),
    .C(_10778_),
    .Y(_11107_));
 sky130_fd_sc_hd__nand2_2 _33143_ (.A(_11106_),
    .B(_11107_),
    .Y(_11108_));
 sky130_fd_sc_hd__a21o_2 _33144_ (.A1(_11108_),
    .A2(_10786_),
    .B1(_10776_),
    .X(_11109_));
 sky130_fd_sc_hd__nand2_2 _33145_ (.A(_11100_),
    .B(_11101_),
    .Y(_11110_));
 sky130_fd_sc_hd__o2111ai_2 _33146_ (.A1(_11096_),
    .A2(_11110_),
    .B1(_11099_),
    .C1(_11015_),
    .D1(_11011_),
    .Y(_11111_));
 sky130_fd_sc_hd__nand3_2 _33147_ (.A(_11105_),
    .B(_11109_),
    .C(_11111_),
    .Y(_11112_));
 sky130_fd_sc_hd__nand3_2 _33148_ (.A(_11016_),
    .B(_11103_),
    .C(_11099_),
    .Y(_11113_));
 sky130_fd_sc_hd__a21oi_2 _33149_ (.A1(_11108_),
    .A2(_10786_),
    .B1(_10776_),
    .Y(_11114_));
 sky130_fd_sc_hd__nand3_2 _33150_ (.A(_11104_),
    .B(_11011_),
    .C(_11015_),
    .Y(_11115_));
 sky130_fd_sc_hd__nand3_2 _33151_ (.A(_11113_),
    .B(_11114_),
    .C(_11115_),
    .Y(_11116_));
 sky130_fd_sc_hd__nand2_2 _33152_ (.A(_10569_),
    .B(_10578_),
    .Y(_11117_));
 sky130_fd_sc_hd__and2b_2 _33153_ (.A_N(_10553_),
    .B(_10557_),
    .X(_11118_));
 sky130_fd_sc_hd__a21o_2 _33154_ (.A1(_11117_),
    .A2(_10576_),
    .B1(_11118_),
    .X(_11119_));
 sky130_fd_sc_hd__nand2_2 _33155_ (.A(_10575_),
    .B(_11118_),
    .Y(_11120_));
 sky130_fd_sc_hd__a21o_2 _33156_ (.A1(_10569_),
    .A2(_10578_),
    .B1(_11120_),
    .X(_11121_));
 sky130_fd_sc_hd__buf_1 _33157_ (.A(_10818_),
    .X(_11122_));
 sky130_fd_sc_hd__buf_1 _33158_ (.A(_11122_),
    .X(_11123_));
 sky130_fd_sc_hd__buf_1 _33159_ (.A(_11123_),
    .X(_11124_));
 sky130_fd_sc_hd__a21oi_2 _33160_ (.A1(_11119_),
    .A2(_11121_),
    .B1(_11124_),
    .Y(_11125_));
 sky130_fd_sc_hd__a21oi_2 _33161_ (.A1(_11117_),
    .A2(_10576_),
    .B1(_11118_),
    .Y(_11126_));
 sky130_fd_sc_hd__nand2_2 _33162_ (.A(_11121_),
    .B(_11124_),
    .Y(_11127_));
 sky130_fd_sc_hd__nor2_2 _33163_ (.A(_11126_),
    .B(_11127_),
    .Y(_11128_));
 sky130_fd_sc_hd__o2bb2ai_2 _33164_ (.A1_N(_11112_),
    .A2_N(_11116_),
    .B1(_11125_),
    .B2(_11128_),
    .Y(_11129_));
 sky130_fd_sc_hd__nor2_2 _33165_ (.A(_11125_),
    .B(_11128_),
    .Y(_11130_));
 sky130_fd_sc_hd__nand3_2 _33166_ (.A(_11116_),
    .B(_11112_),
    .C(_11130_),
    .Y(_11131_));
 sky130_fd_sc_hd__a21o_2 _33167_ (.A1(_10798_),
    .A2(_10800_),
    .B1(_10793_),
    .X(_11132_));
 sky130_fd_sc_hd__a21o_2 _33168_ (.A1(_11129_),
    .A2(_11131_),
    .B1(_11132_),
    .X(_11133_));
 sky130_fd_sc_hd__nand3_2 _33169_ (.A(_11129_),
    .B(_11132_),
    .C(_11131_),
    .Y(_11134_));
 sky130_fd_sc_hd__inv_2 _33170_ (.A(_10476_),
    .Y(_11135_));
 sky130_fd_sc_hd__a21o_2 _33171_ (.A1(_11133_),
    .A2(_11134_),
    .B1(_11135_),
    .X(_11136_));
 sky130_fd_sc_hd__nand3_2 _33172_ (.A(_11133_),
    .B(_11135_),
    .C(_11134_),
    .Y(_11137_));
 sky130_fd_sc_hd__nand3b_2 _33173_ (.A_N(_10815_),
    .B(_11136_),
    .C(_11137_),
    .Y(_11138_));
 sky130_fd_sc_hd__o2bb2ai_2 _33174_ (.A1_N(_11134_),
    .A2_N(_11133_),
    .B1(_10475_),
    .B2(_10474_),
    .Y(_11139_));
 sky130_fd_sc_hd__nand3_2 _33175_ (.A(_11133_),
    .B(_10476_),
    .C(_11134_),
    .Y(_11140_));
 sky130_fd_sc_hd__nand3_2 _33176_ (.A(_11139_),
    .B(_11140_),
    .C(_10815_),
    .Y(_11141_));
 sky130_fd_sc_hd__nand2_2 _33177_ (.A(_11138_),
    .B(_11141_),
    .Y(_11142_));
 sky130_fd_sc_hd__a21o_2 _33178_ (.A1(_08035_),
    .A2(_08028_),
    .B1(_08031_),
    .X(_11143_));
 sky130_fd_sc_hd__o2111ai_2 _33179_ (.A1(_08293_),
    .A2(_08296_),
    .B1(_08302_),
    .C1(_08300_),
    .D1(_11143_),
    .Y(_11144_));
 sky130_fd_sc_hd__nor3_2 _33180_ (.A(_08041_),
    .B(_11144_),
    .C(_07544_),
    .Y(_11145_));
 sky130_fd_sc_hd__inv_2 _33181_ (.A(_10808_),
    .Y(_11146_));
 sky130_fd_sc_hd__nand2_2 _33182_ (.A(_10807_),
    .B(_10809_),
    .Y(_11147_));
 sky130_fd_sc_hd__o2111ai_2 _33183_ (.A1(_11146_),
    .A2(_11147_),
    .B1(_10464_),
    .C1(_10460_),
    .D1(_10810_),
    .Y(_11148_));
 sky130_fd_sc_hd__nor3_2 _33184_ (.A(_10468_),
    .B(_11148_),
    .C(_09811_),
    .Y(_11149_));
 sky130_fd_sc_hd__o2111ai_2 _33185_ (.A1(_06318_),
    .A2(_06485_),
    .B1(_11145_),
    .C1(_06490_),
    .D1(_11149_),
    .Y(_11150_));
 sky130_fd_sc_hd__nand2_2 _33186_ (.A(_08587_),
    .B(_11149_),
    .Y(_11151_));
 sky130_fd_sc_hd__nor2_2 _33187_ (.A(_10468_),
    .B(_11148_),
    .Y(_11152_));
 sky130_fd_sc_hd__a21oi_2 _33188_ (.A1(_10807_),
    .A2(_10808_),
    .B1(_10809_),
    .Y(_11153_));
 sky130_fd_sc_hd__o21a_2 _33189_ (.A1(_10464_),
    .A2(_11153_),
    .B1(_10811_),
    .X(_11154_));
 sky130_fd_sc_hd__o21ai_2 _33190_ (.A1(_10470_),
    .A2(_11148_),
    .B1(_11154_),
    .Y(_11155_));
 sky130_fd_sc_hd__a21oi_2 _33191_ (.A1(_09810_),
    .A2(_11152_),
    .B1(_11155_),
    .Y(_11156_));
 sky130_fd_sc_hd__nand3_2 _33192_ (.A(_11150_),
    .B(_11151_),
    .C(_11156_),
    .Y(_11157_));
 sky130_fd_sc_hd__xnor2_2 _33193_ (.A(_11142_),
    .B(_11157_),
    .Y(_02651_));
 sky130_fd_sc_hd__and3_2 _33194_ (.A(_11117_),
    .B(_10576_),
    .C(_11118_),
    .X(_11158_));
 sky130_fd_sc_hd__nor2_2 _33195_ (.A(_11124_),
    .B(_11126_),
    .Y(_11159_));
 sky130_fd_sc_hd__nand3_2 _33196_ (.A(_11015_),
    .B(_11099_),
    .C(_11103_),
    .Y(_11160_));
 sky130_fd_sc_hd__nand2_2 _33197_ (.A(_11160_),
    .B(_11011_),
    .Y(_11161_));
 sky130_fd_sc_hd__o21ai_2 _33198_ (.A1(_11005_),
    .A2(_11009_),
    .B1(_11003_),
    .Y(_11162_));
 sky130_fd_sc_hd__and4b_2 _33199_ (.A_N(_05105_),
    .B(_10817_),
    .C(_10822_),
    .D(_05248_),
    .X(_11163_));
 sky130_fd_sc_hd__buf_1 _33200_ (.A(_10831_),
    .X(_11164_));
 sky130_fd_sc_hd__o22a_2 _33201_ (.A1(_07904_),
    .A2(_18181_),
    .B1(_11164_),
    .B2(_05100_),
    .X(_11165_));
 sky130_fd_sc_hd__nand2_2 _33202_ (.A(_19311_),
    .B(_06447_),
    .Y(_11166_));
 sky130_fd_sc_hd__inv_2 _33203_ (.A(_11166_),
    .Y(_11167_));
 sky130_fd_sc_hd__o21ai_2 _33204_ (.A1(_11163_),
    .A2(_11165_),
    .B1(_11167_),
    .Y(_11168_));
 sky130_fd_sc_hd__buf_1 _33205_ (.A(_10817_),
    .X(_11169_));
 sky130_fd_sc_hd__a22o_2 _33206_ (.A1(_10823_),
    .A2(_08393_),
    .B1(_05106_),
    .B2(_11169_),
    .X(_11170_));
 sky130_fd_sc_hd__nand3b_2 _33207_ (.A_N(_11163_),
    .B(_11170_),
    .C(_11166_),
    .Y(_11171_));
 sky130_fd_sc_hd__o21ai_2 _33208_ (.A1(_19641_),
    .A2(_10819_),
    .B1(_10816_),
    .Y(_11172_));
 sky130_fd_sc_hd__nand2_2 _33209_ (.A(_10825_),
    .B(_11172_),
    .Y(_11173_));
 sky130_fd_sc_hd__nand3_2 _33210_ (.A(_11168_),
    .B(_11171_),
    .C(_11173_),
    .Y(_11174_));
 sky130_fd_sc_hd__o21ai_2 _33211_ (.A1(_11163_),
    .A2(_11165_),
    .B1(_11166_),
    .Y(_11175_));
 sky130_fd_sc_hd__nand3b_2 _33212_ (.A_N(_11163_),
    .B(_11170_),
    .C(_11167_),
    .Y(_11176_));
 sky130_fd_sc_hd__nand3b_2 _33213_ (.A_N(_11173_),
    .B(_11175_),
    .C(_11176_),
    .Y(_11177_));
 sky130_fd_sc_hd__buf_1 _33214_ (.A(_10703_),
    .X(_11178_));
 sky130_fd_sc_hd__a22o_2 _33215_ (.A1(_10138_),
    .A2(_05222_),
    .B1(_10141_),
    .B2(_05269_),
    .X(_11179_));
 sky130_fd_sc_hd__o21ai_2 _33216_ (.A1(_07651_),
    .A2(_11178_),
    .B1(_11179_),
    .Y(_11180_));
 sky130_fd_sc_hd__nor2_2 _33217_ (.A(_09356_),
    .B(_05260_),
    .Y(_11181_));
 sky130_fd_sc_hd__nand2_2 _33218_ (.A(_11180_),
    .B(_11181_),
    .Y(_11182_));
 sky130_fd_sc_hd__inv_2 _33219_ (.A(_11182_),
    .Y(_11183_));
 sky130_fd_sc_hd__o21a_2 _33220_ (.A1(_07651_),
    .A2(_10704_),
    .B1(_11179_),
    .X(_11184_));
 sky130_fd_sc_hd__inv_2 _33221_ (.A(_11181_),
    .Y(_11185_));
 sky130_fd_sc_hd__nand2_2 _33222_ (.A(_11184_),
    .B(_11185_),
    .Y(_11186_));
 sky130_fd_sc_hd__inv_2 _33223_ (.A(_11186_),
    .Y(_11187_));
 sky130_fd_sc_hd__o2bb2ai_2 _33224_ (.A1_N(_11174_),
    .A2_N(_11177_),
    .B1(_11183_),
    .B2(_11187_),
    .Y(_11188_));
 sky130_fd_sc_hd__a21oi_2 _33225_ (.A1(_10821_),
    .A2(_10825_),
    .B1(_10828_),
    .Y(_11189_));
 sky130_fd_sc_hd__a21oi_2 _33226_ (.A1(_10836_),
    .A2(_10851_),
    .B1(_11189_),
    .Y(_11190_));
 sky130_fd_sc_hd__nand2_2 _33227_ (.A(_11186_),
    .B(_11182_),
    .Y(_11191_));
 sky130_fd_sc_hd__nand3b_2 _33228_ (.A_N(_11191_),
    .B(_11174_),
    .C(_11177_),
    .Y(_11192_));
 sky130_fd_sc_hd__nand3_2 _33229_ (.A(_11188_),
    .B(_11190_),
    .C(_11192_),
    .Y(_11193_));
 sky130_fd_sc_hd__nor2_2 _33230_ (.A(_11181_),
    .B(_11184_),
    .Y(_11194_));
 sky130_fd_sc_hd__nor2_2 _33231_ (.A(_11180_),
    .B(_11185_),
    .Y(_11195_));
 sky130_fd_sc_hd__o2bb2ai_2 _33232_ (.A1_N(_11174_),
    .A2_N(_11177_),
    .B1(_11194_),
    .B2(_11195_),
    .Y(_11196_));
 sky130_fd_sc_hd__a21o_2 _33233_ (.A1(_10836_),
    .A2(_10851_),
    .B1(_11189_),
    .X(_11197_));
 sky130_fd_sc_hd__nand3_2 _33234_ (.A(_11177_),
    .B(_11174_),
    .C(_11191_),
    .Y(_11198_));
 sky130_fd_sc_hd__nand3_2 _33235_ (.A(_11196_),
    .B(_11197_),
    .C(_11198_),
    .Y(_11199_));
 sky130_fd_sc_hd__a21oi_2 _33236_ (.A1(_10838_),
    .A2(_10842_),
    .B1(_10841_),
    .Y(_11200_));
 sky130_fd_sc_hd__a22oi_2 _33237_ (.A1(_09819_),
    .A2(_05505_),
    .B1(_19331_),
    .B2(_05613_),
    .Y(_11201_));
 sky130_fd_sc_hd__and4_2 _33238_ (.A(_10166_),
    .B(_09827_),
    .C(_06052_),
    .D(_05505_),
    .X(_11202_));
 sky130_fd_sc_hd__nand2_2 _33239_ (.A(_10862_),
    .B(_05615_),
    .Y(_11203_));
 sky130_fd_sc_hd__o21ai_2 _33240_ (.A1(_11201_),
    .A2(_11202_),
    .B1(_11203_),
    .Y(_11204_));
 sky130_fd_sc_hd__buf_1 _33241_ (.A(_19327_),
    .X(_11205_));
 sky130_fd_sc_hd__a22o_2 _33242_ (.A1(_11205_),
    .A2(_19620_),
    .B1(_10867_),
    .B2(_19617_),
    .X(_11206_));
 sky130_fd_sc_hd__inv_2 _33243_ (.A(_11203_),
    .Y(_11207_));
 sky130_fd_sc_hd__nand3b_2 _33244_ (.A_N(_11202_),
    .B(_11206_),
    .C(_11207_),
    .Y(_11208_));
 sky130_fd_sc_hd__nand3b_2 _33245_ (.A_N(_11200_),
    .B(_11204_),
    .C(_11208_),
    .Y(_11209_));
 sky130_fd_sc_hd__nand3b_2 _33246_ (.A_N(_11202_),
    .B(_11206_),
    .C(_11203_),
    .Y(_11210_));
 sky130_fd_sc_hd__o21ai_2 _33247_ (.A1(_11201_),
    .A2(_11202_),
    .B1(_11207_),
    .Y(_11211_));
 sky130_fd_sc_hd__nand3_2 _33248_ (.A(_11210_),
    .B(_11200_),
    .C(_11211_),
    .Y(_11212_));
 sky130_fd_sc_hd__a21oi_2 _33249_ (.A1(_10864_),
    .A2(_10865_),
    .B1(_10861_),
    .Y(_11213_));
 sky130_fd_sc_hd__inv_2 _33250_ (.A(_11213_),
    .Y(_11214_));
 sky130_fd_sc_hd__a21oi_2 _33251_ (.A1(_11209_),
    .A2(_11212_),
    .B1(_11214_),
    .Y(_11215_));
 sky130_fd_sc_hd__and3_2 _33252_ (.A(_11209_),
    .B(_11212_),
    .C(_11214_),
    .X(_11216_));
 sky130_fd_sc_hd__o2bb2ai_2 _33253_ (.A1_N(_11193_),
    .A2_N(_11199_),
    .B1(_11215_),
    .B2(_11216_),
    .Y(_11217_));
 sky130_fd_sc_hd__inv_2 _33254_ (.A(_10852_),
    .Y(_11218_));
 sky130_fd_sc_hd__nand2_2 _33255_ (.A(_10847_),
    .B(_10848_),
    .Y(_11219_));
 sky130_fd_sc_hd__o2bb2ai_2 _33256_ (.A1_N(_10857_),
    .A2_N(_10885_),
    .B1(_11218_),
    .B2(_11219_),
    .Y(_11220_));
 sky130_fd_sc_hd__nor2_2 _33257_ (.A(_11215_),
    .B(_11216_),
    .Y(_11221_));
 sky130_fd_sc_hd__nand3_2 _33258_ (.A(_11199_),
    .B(_11193_),
    .C(_11221_),
    .Y(_11222_));
 sky130_fd_sc_hd__nand3_2 _33259_ (.A(_11217_),
    .B(_11220_),
    .C(_11222_),
    .Y(_11223_));
 sky130_fd_sc_hd__buf_1 _33260_ (.A(_11223_),
    .X(_11224_));
 sky130_fd_sc_hd__and2_2 _33261_ (.A(_11212_),
    .B(_11214_),
    .X(_11225_));
 sky130_fd_sc_hd__a21o_2 _33262_ (.A1(_11225_),
    .A2(_11209_),
    .B1(_11215_),
    .X(_11226_));
 sky130_fd_sc_hd__a21o_2 _33263_ (.A1(_11199_),
    .A2(_11193_),
    .B1(_11226_),
    .X(_11227_));
 sky130_fd_sc_hd__a21boi_2 _33264_ (.A1(_10885_),
    .A2(_10857_),
    .B1_N(_10853_),
    .Y(_11228_));
 sky130_fd_sc_hd__nand3_2 _33265_ (.A(_11199_),
    .B(_11226_),
    .C(_11193_),
    .Y(_11229_));
 sky130_fd_sc_hd__nand3_2 _33266_ (.A(_11227_),
    .B(_11228_),
    .C(_11229_),
    .Y(_11230_));
 sky130_fd_sc_hd__nand2_2 _33267_ (.A(_08385_),
    .B(_19609_),
    .Y(_11231_));
 sky130_fd_sc_hd__nand2_2 _33268_ (.A(_08386_),
    .B(_19606_),
    .Y(_11232_));
 sky130_fd_sc_hd__nor2_2 _33269_ (.A(_11231_),
    .B(_11232_),
    .Y(_11233_));
 sky130_fd_sc_hd__nand2_2 _33270_ (.A(_07976_),
    .B(_05897_),
    .Y(_11234_));
 sky130_fd_sc_hd__inv_2 _33271_ (.A(_11234_),
    .Y(_11235_));
 sky130_fd_sc_hd__nand2_2 _33272_ (.A(_11231_),
    .B(_11232_),
    .Y(_11236_));
 sky130_fd_sc_hd__nand2_2 _33273_ (.A(_11235_),
    .B(_11236_),
    .Y(_11237_));
 sky130_fd_sc_hd__a21o_2 _33274_ (.A1(_10900_),
    .A2(_10898_),
    .B1(_10897_),
    .X(_11238_));
 sky130_fd_sc_hd__and2_2 _33275_ (.A(_11231_),
    .B(_11232_),
    .X(_11239_));
 sky130_fd_sc_hd__o21ai_2 _33276_ (.A1(_11233_),
    .A2(_11239_),
    .B1(_11234_),
    .Y(_11240_));
 sky130_fd_sc_hd__o211ai_2 _33277_ (.A1(_11233_),
    .A2(_11237_),
    .B1(_11238_),
    .C1(_11240_),
    .Y(_11241_));
 sky130_fd_sc_hd__o21ai_2 _33278_ (.A1(_11233_),
    .A2(_11239_),
    .B1(_11235_),
    .Y(_11242_));
 sky130_fd_sc_hd__nand3b_2 _33279_ (.A_N(_11233_),
    .B(_11236_),
    .C(_11234_),
    .Y(_11243_));
 sky130_fd_sc_hd__a21oi_2 _33280_ (.A1(_10900_),
    .A2(_10898_),
    .B1(_10897_),
    .Y(_11244_));
 sky130_fd_sc_hd__nand3_2 _33281_ (.A(_11242_),
    .B(_11243_),
    .C(_11244_),
    .Y(_11245_));
 sky130_fd_sc_hd__nand2_2 _33282_ (.A(_08808_),
    .B(_06736_),
    .Y(_11246_));
 sky130_fd_sc_hd__nand2_2 _33283_ (.A(_08185_),
    .B(_06935_),
    .Y(_11247_));
 sky130_fd_sc_hd__nor2_2 _33284_ (.A(_11246_),
    .B(_11247_),
    .Y(_11248_));
 sky130_fd_sc_hd__and2_2 _33285_ (.A(_11246_),
    .B(_11247_),
    .X(_11249_));
 sky130_fd_sc_hd__nor2_2 _33286_ (.A(_11248_),
    .B(_11249_),
    .Y(_11250_));
 sky130_fd_sc_hd__buf_1 _33287_ (.A(_07052_),
    .X(_11251_));
 sky130_fd_sc_hd__nor2_2 _33288_ (.A(_11251_),
    .B(_06958_),
    .Y(_11252_));
 sky130_fd_sc_hd__inv_2 _33289_ (.A(_11252_),
    .Y(_11253_));
 sky130_fd_sc_hd__nand2_2 _33290_ (.A(_11250_),
    .B(_11253_),
    .Y(_11254_));
 sky130_fd_sc_hd__o21ai_2 _33291_ (.A1(_11248_),
    .A2(_11249_),
    .B1(_11252_),
    .Y(_11255_));
 sky130_fd_sc_hd__nand2_2 _33292_ (.A(_11254_),
    .B(_11255_),
    .Y(_11256_));
 sky130_fd_sc_hd__a21o_2 _33293_ (.A1(_11241_),
    .A2(_11245_),
    .B1(_11256_),
    .X(_11257_));
 sky130_fd_sc_hd__nand3_2 _33294_ (.A(_11256_),
    .B(_11241_),
    .C(_11245_),
    .Y(_11258_));
 sky130_fd_sc_hd__nand2_2 _33295_ (.A(_11257_),
    .B(_11258_),
    .Y(_11259_));
 sky130_fd_sc_hd__nor2_2 _33296_ (.A(_10872_),
    .B(_10884_),
    .Y(_11260_));
 sky130_fd_sc_hd__nand2_2 _33297_ (.A(_11259_),
    .B(_11260_),
    .Y(_11261_));
 sky130_fd_sc_hd__nand2_2 _33298_ (.A(_10877_),
    .B(_10880_),
    .Y(_11262_));
 sky130_fd_sc_hd__nand3_2 _33299_ (.A(_11262_),
    .B(_11258_),
    .C(_11257_),
    .Y(_11263_));
 sky130_fd_sc_hd__nand2_2 _33300_ (.A(_10917_),
    .B(_10907_),
    .Y(_11264_));
 sky130_fd_sc_hd__nand2_2 _33301_ (.A(_11264_),
    .B(_10904_),
    .Y(_11265_));
 sky130_fd_sc_hd__nand3_2 _33302_ (.A(_11261_),
    .B(_11263_),
    .C(_11265_),
    .Y(_11266_));
 sky130_fd_sc_hd__inv_2 _33303_ (.A(_11266_),
    .Y(_11267_));
 sky130_fd_sc_hd__a21oi_2 _33304_ (.A1(_11261_),
    .A2(_11263_),
    .B1(_11265_),
    .Y(_11268_));
 sky130_fd_sc_hd__o2bb2ai_2 _33305_ (.A1_N(_11224_),
    .A2_N(_11230_),
    .B1(_11267_),
    .B2(_11268_),
    .Y(_11269_));
 sky130_fd_sc_hd__inv_2 _33306_ (.A(_10886_),
    .Y(_11270_));
 sky130_fd_sc_hd__nand2_2 _33307_ (.A(_10882_),
    .B(_10887_),
    .Y(_11271_));
 sky130_fd_sc_hd__nand2_2 _33308_ (.A(_10923_),
    .B(_10926_),
    .Y(_11272_));
 sky130_fd_sc_hd__nand2_2 _33309_ (.A(_11272_),
    .B(_10933_),
    .Y(_11273_));
 sky130_fd_sc_hd__nand2_2 _33310_ (.A(_11273_),
    .B(_10930_),
    .Y(_11274_));
 sky130_fd_sc_hd__a21oi_2 _33311_ (.A1(_10882_),
    .A2(_10886_),
    .B1(_10887_),
    .Y(_11275_));
 sky130_fd_sc_hd__o22ai_2 _33312_ (.A1(_11270_),
    .A2(_11271_),
    .B1(_11274_),
    .B2(_11275_),
    .Y(_11276_));
 sky130_fd_sc_hd__inv_2 _33313_ (.A(_11265_),
    .Y(_11277_));
 sky130_fd_sc_hd__a21oi_2 _33314_ (.A1(_11257_),
    .A2(_11258_),
    .B1(_11262_),
    .Y(_11278_));
 sky130_fd_sc_hd__nor2_2 _33315_ (.A(_11277_),
    .B(_11278_),
    .Y(_11279_));
 sky130_fd_sc_hd__a21oi_2 _33316_ (.A1(_11263_),
    .A2(_11279_),
    .B1(_11268_),
    .Y(_11280_));
 sky130_fd_sc_hd__nand3_2 _33317_ (.A(_11280_),
    .B(_11230_),
    .C(_11224_),
    .Y(_11281_));
 sky130_fd_sc_hd__nand3_2 _33318_ (.A(_11269_),
    .B(_11276_),
    .C(_11281_),
    .Y(_11282_));
 sky130_fd_sc_hd__nand2_2 _33319_ (.A(_11230_),
    .B(_11223_),
    .Y(_11283_));
 sky130_fd_sc_hd__nand2_2 _33320_ (.A(_11283_),
    .B(_11280_),
    .Y(_11284_));
 sky130_fd_sc_hd__a21boi_2 _33321_ (.A1(_10936_),
    .A2(_10893_),
    .B1_N(_10888_),
    .Y(_11285_));
 sky130_fd_sc_hd__inv_2 _33322_ (.A(_10907_),
    .Y(_11286_));
 sky130_fd_sc_hd__and3_2 _33323_ (.A(_10904_),
    .B(_10915_),
    .C(_10916_),
    .X(_11287_));
 sky130_fd_sc_hd__o2bb2ai_2 _33324_ (.A1_N(_11263_),
    .A2_N(_11261_),
    .B1(_11286_),
    .B2(_11287_),
    .Y(_11288_));
 sky130_fd_sc_hd__nand2_2 _33325_ (.A(_11288_),
    .B(_11266_),
    .Y(_11289_));
 sky130_fd_sc_hd__nand3_2 _33326_ (.A(_11289_),
    .B(_11230_),
    .C(_11224_),
    .Y(_11290_));
 sky130_fd_sc_hd__nand3_2 _33327_ (.A(_11284_),
    .B(_11285_),
    .C(_11290_),
    .Y(_11291_));
 sky130_fd_sc_hd__a21oi_2 _33328_ (.A1(_10989_),
    .A2(_10990_),
    .B1(_10960_),
    .Y(_11292_));
 sky130_fd_sc_hd__inv_2 _33329_ (.A(_11292_),
    .Y(_11293_));
 sky130_fd_sc_hd__nand2_2 _33330_ (.A(_08182_),
    .B(_06542_),
    .Y(_11294_));
 sky130_fd_sc_hd__nand2_2 _33331_ (.A(_19357_),
    .B(_19588_),
    .Y(_11295_));
 sky130_fd_sc_hd__nor2_2 _33332_ (.A(_11294_),
    .B(_11295_),
    .Y(_11296_));
 sky130_fd_sc_hd__nor2_2 _33333_ (.A(_08352_),
    .B(_08598_),
    .Y(_11297_));
 sky130_fd_sc_hd__nand2_2 _33334_ (.A(_11294_),
    .B(_11295_),
    .Y(_11298_));
 sky130_fd_sc_hd__nand3b_2 _33335_ (.A_N(_11296_),
    .B(_11297_),
    .C(_11298_),
    .Y(_11299_));
 sky130_fd_sc_hd__buf_1 _33336_ (.A(_06831_),
    .X(_11300_));
 sky130_fd_sc_hd__a21o_2 _33337_ (.A1(_09019_),
    .A2(_06945_),
    .B1(_11294_),
    .X(_11301_));
 sky130_fd_sc_hd__a21o_2 _33338_ (.A1(_09018_),
    .A2(_06950_),
    .B1(_11295_),
    .X(_11302_));
 sky130_fd_sc_hd__o211ai_2 _33339_ (.A1(_11300_),
    .A2(_08611_),
    .B1(_11301_),
    .C1(_11302_),
    .Y(_11303_));
 sky130_fd_sc_hd__a21o_2 _33340_ (.A1(_10914_),
    .A2(_10911_),
    .B1(_10910_),
    .X(_11304_));
 sky130_fd_sc_hd__a21oi_2 _33341_ (.A1(_11299_),
    .A2(_11303_),
    .B1(_11304_),
    .Y(_11305_));
 sky130_fd_sc_hd__nand3_2 _33342_ (.A(_11299_),
    .B(_11304_),
    .C(_11303_),
    .Y(_11306_));
 sky130_fd_sc_hd__a21oi_2 _33343_ (.A1(_10942_),
    .A2(_10947_),
    .B1(_10946_),
    .Y(_11307_));
 sky130_fd_sc_hd__nand2_2 _33344_ (.A(_11306_),
    .B(_11307_),
    .Y(_11308_));
 sky130_fd_sc_hd__a21oi_2 _33345_ (.A1(_10952_),
    .A2(_10953_),
    .B1(_10958_),
    .Y(_11309_));
 sky130_fd_sc_hd__and3_2 _33346_ (.A(_11299_),
    .B(_11304_),
    .C(_11303_),
    .X(_11310_));
 sky130_fd_sc_hd__inv_2 _33347_ (.A(_11307_),
    .Y(_11311_));
 sky130_fd_sc_hd__o21ai_2 _33348_ (.A1(_11305_),
    .A2(_11310_),
    .B1(_11311_),
    .Y(_11312_));
 sky130_fd_sc_hd__o211ai_2 _33349_ (.A1(_11305_),
    .A2(_11308_),
    .B1(_11309_),
    .C1(_11312_),
    .Y(_11313_));
 sky130_fd_sc_hd__o21ai_2 _33350_ (.A1(_11305_),
    .A2(_11310_),
    .B1(_11307_),
    .Y(_11314_));
 sky130_fd_sc_hd__nand3b_2 _33351_ (.A_N(_11305_),
    .B(_11306_),
    .C(_11311_),
    .Y(_11315_));
 sky130_fd_sc_hd__nand2_2 _33352_ (.A(_10959_),
    .B(_10949_),
    .Y(_11316_));
 sky130_fd_sc_hd__nand3_2 _33353_ (.A(_11314_),
    .B(_11315_),
    .C(_11316_),
    .Y(_11317_));
 sky130_fd_sc_hd__nand2_2 _33354_ (.A(_11313_),
    .B(_11317_),
    .Y(_11318_));
 sky130_fd_sc_hd__nand2_2 _33355_ (.A(_09051_),
    .B(_08103_),
    .Y(_11319_));
 sky130_fd_sc_hd__nand2_2 _33356_ (.A(_06433_),
    .B(_09199_),
    .Y(_11320_));
 sky130_fd_sc_hd__nor2_2 _33357_ (.A(_11319_),
    .B(_11320_),
    .Y(_11321_));
 sky130_fd_sc_hd__and2_2 _33358_ (.A(_11319_),
    .B(_11320_),
    .X(_11322_));
 sky130_fd_sc_hd__nand2_2 _33359_ (.A(_06616_),
    .B(_19567_),
    .Y(_11323_));
 sky130_fd_sc_hd__inv_2 _33360_ (.A(_11323_),
    .Y(_11324_));
 sky130_fd_sc_hd__o21ai_2 _33361_ (.A1(_11321_),
    .A2(_11322_),
    .B1(_11324_),
    .Y(_11325_));
 sky130_fd_sc_hd__nand2_2 _33362_ (.A(_11319_),
    .B(_11320_),
    .Y(_11326_));
 sky130_fd_sc_hd__nand3b_2 _33363_ (.A_N(_11321_),
    .B(_11323_),
    .C(_11326_),
    .Y(_11327_));
 sky130_fd_sc_hd__nand2_2 _33364_ (.A(_11325_),
    .B(_11327_),
    .Y(_11328_));
 sky130_fd_sc_hd__nand3_2 _33365_ (.A(_08315_),
    .B(_07934_),
    .C(_19582_),
    .Y(_11329_));
 sky130_fd_sc_hd__nor2_2 _33366_ (.A(_09246_),
    .B(_11329_),
    .Y(_11330_));
 sky130_fd_sc_hd__a22o_2 _33367_ (.A1(_06271_),
    .A2(_08490_),
    .B1(_06273_),
    .B2(_08108_),
    .X(_11331_));
 sky130_fd_sc_hd__nand2_2 _33368_ (.A(_19368_),
    .B(_08651_),
    .Y(_11332_));
 sky130_fd_sc_hd__inv_2 _33369_ (.A(_11332_),
    .Y(_11333_));
 sky130_fd_sc_hd__nand2_2 _33370_ (.A(_11331_),
    .B(_11333_),
    .Y(_11334_));
 sky130_fd_sc_hd__a21o_2 _33371_ (.A1(_10973_),
    .A2(_10975_),
    .B1(_10972_),
    .X(_11335_));
 sky130_fd_sc_hd__o21ai_2 _33372_ (.A1(_09263_),
    .A2(_11329_),
    .B1(_11331_),
    .Y(_11336_));
 sky130_fd_sc_hd__nand2_2 _33373_ (.A(_11336_),
    .B(_11332_),
    .Y(_11337_));
 sky130_fd_sc_hd__o211ai_2 _33374_ (.A1(_11330_),
    .A2(_11334_),
    .B1(_11335_),
    .C1(_11337_),
    .Y(_11338_));
 sky130_fd_sc_hd__nand2_2 _33375_ (.A(_11336_),
    .B(_11333_),
    .Y(_11339_));
 sky130_fd_sc_hd__nand3b_2 _33376_ (.A_N(_11330_),
    .B(_11331_),
    .C(_11332_),
    .Y(_11340_));
 sky130_fd_sc_hd__a21oi_2 _33377_ (.A1(_10973_),
    .A2(_10975_),
    .B1(_10972_),
    .Y(_11341_));
 sky130_fd_sc_hd__nand3_2 _33378_ (.A(_11339_),
    .B(_11340_),
    .C(_11341_),
    .Y(_11342_));
 sky130_fd_sc_hd__nand2_2 _33379_ (.A(_11338_),
    .B(_11342_),
    .Y(_11343_));
 sky130_fd_sc_hd__xnor2_2 _33380_ (.A(_11328_),
    .B(_11343_),
    .Y(_11344_));
 sky130_fd_sc_hd__nand2_2 _33381_ (.A(_11318_),
    .B(_11344_),
    .Y(_11345_));
 sky130_fd_sc_hd__a21boi_2 _33382_ (.A1(_10923_),
    .A2(_10928_),
    .B1_N(_10926_),
    .Y(_11346_));
 sky130_fd_sc_hd__xor2_2 _33383_ (.A(_11328_),
    .B(_11343_),
    .X(_11347_));
 sky130_fd_sc_hd__nand3_2 _33384_ (.A(_11347_),
    .B(_11313_),
    .C(_11317_),
    .Y(_11348_));
 sky130_fd_sc_hd__nand3_2 _33385_ (.A(_11345_),
    .B(_11346_),
    .C(_11348_),
    .Y(_11349_));
 sky130_fd_sc_hd__nand2_2 _33386_ (.A(_11293_),
    .B(_11349_),
    .Y(_11350_));
 sky130_fd_sc_hd__nand2_2 _33387_ (.A(_10930_),
    .B(_10926_),
    .Y(_11351_));
 sky130_fd_sc_hd__nand3_2 _33388_ (.A(_11344_),
    .B(_11313_),
    .C(_11317_),
    .Y(_11352_));
 sky130_fd_sc_hd__nand2_2 _33389_ (.A(_11318_),
    .B(_11347_),
    .Y(_11353_));
 sky130_fd_sc_hd__nand3_2 _33390_ (.A(_11351_),
    .B(_11352_),
    .C(_11353_),
    .Y(_11354_));
 sky130_fd_sc_hd__inv_2 _33391_ (.A(_11354_),
    .Y(_11355_));
 sky130_fd_sc_hd__nor2_2 _33392_ (.A(_11350_),
    .B(_11355_),
    .Y(_11356_));
 sky130_fd_sc_hd__a21oi_2 _33393_ (.A1(_11354_),
    .A2(_11349_),
    .B1(_11293_),
    .Y(_11357_));
 sky130_fd_sc_hd__o2bb2ai_2 _33394_ (.A1_N(_11282_),
    .A2_N(_11291_),
    .B1(_11356_),
    .B2(_11357_),
    .Y(_11358_));
 sky130_fd_sc_hd__a31oi_2 _33395_ (.A1(_11345_),
    .A2(_11346_),
    .A3(_11348_),
    .B1(_11292_),
    .Y(_11359_));
 sky130_fd_sc_hd__a21oi_2 _33396_ (.A1(_11354_),
    .A2(_11359_),
    .B1(_11357_),
    .Y(_11360_));
 sky130_fd_sc_hd__nand3_2 _33397_ (.A(_11360_),
    .B(_11291_),
    .C(_11282_),
    .Y(_11361_));
 sky130_fd_sc_hd__nand3_2 _33398_ (.A(_11162_),
    .B(_11358_),
    .C(_11361_),
    .Y(_11362_));
 sky130_fd_sc_hd__a21oi_2 _33399_ (.A1(_10939_),
    .A2(_11002_),
    .B1(_11006_),
    .Y(_11363_));
 sky130_fd_sc_hd__nand2_2 _33400_ (.A(_11291_),
    .B(_11282_),
    .Y(_11364_));
 sky130_fd_sc_hd__nand2_2 _33401_ (.A(_11364_),
    .B(_11360_),
    .Y(_11365_));
 sky130_fd_sc_hd__a21o_2 _33402_ (.A1(_11354_),
    .A2(_11349_),
    .B1(_11293_),
    .X(_11366_));
 sky130_fd_sc_hd__o21ai_2 _33403_ (.A1(_11350_),
    .A2(_11355_),
    .B1(_11366_),
    .Y(_11367_));
 sky130_fd_sc_hd__nand3_2 _33404_ (.A(_11367_),
    .B(_11291_),
    .C(_11282_),
    .Y(_11368_));
 sky130_fd_sc_hd__nand3_2 _33405_ (.A(_11363_),
    .B(_11365_),
    .C(_11368_),
    .Y(_11369_));
 sky130_fd_sc_hd__nand2_2 _33406_ (.A(_19380_),
    .B(_19564_),
    .Y(_11370_));
 sky130_fd_sc_hd__nand2_2 _33407_ (.A(_09247_),
    .B(_19561_),
    .Y(_11371_));
 sky130_fd_sc_hd__nor2_2 _33408_ (.A(_11370_),
    .B(_11371_),
    .Y(_11372_));
 sky130_fd_sc_hd__and2_2 _33409_ (.A(_11370_),
    .B(_11371_),
    .X(_11373_));
 sky130_fd_sc_hd__inv_2 _33410_ (.A(_19557_),
    .Y(_11374_));
 sky130_fd_sc_hd__nor2_2 _33411_ (.A(_05244_),
    .B(_11374_),
    .Y(_11375_));
 sky130_fd_sc_hd__o21bai_2 _33412_ (.A1(_11372_),
    .A2(_11373_),
    .B1_N(_11375_),
    .Y(_11376_));
 sky130_fd_sc_hd__or2_2 _33413_ (.A(_11370_),
    .B(_11371_),
    .X(_11377_));
 sky130_fd_sc_hd__nand2_2 _33414_ (.A(_11370_),
    .B(_11371_),
    .Y(_11378_));
 sky130_fd_sc_hd__nand3_2 _33415_ (.A(_11377_),
    .B(_11375_),
    .C(_11378_),
    .Y(_11379_));
 sky130_fd_sc_hd__a31o_2 _33416_ (.A1(_10964_),
    .A2(_19377_),
    .A3(_19572_),
    .B1(_10963_),
    .X(_11380_));
 sky130_fd_sc_hd__a21oi_2 _33417_ (.A1(_11376_),
    .A2(_11379_),
    .B1(_11380_),
    .Y(_11381_));
 sky130_fd_sc_hd__and3_2 _33418_ (.A(_10964_),
    .B(_19377_),
    .C(_10966_),
    .X(_11382_));
 sky130_fd_sc_hd__o211a_2 _33419_ (.A1(_10963_),
    .A2(_11382_),
    .B1(_11376_),
    .C1(_11379_),
    .X(_11383_));
 sky130_fd_sc_hd__a21oi_2 _33420_ (.A1(_11056_),
    .A2(_11061_),
    .B1(_11060_),
    .Y(_11384_));
 sky130_fd_sc_hd__inv_2 _33421_ (.A(_11384_),
    .Y(_11385_));
 sky130_fd_sc_hd__o21ai_2 _33422_ (.A1(_11381_),
    .A2(_11383_),
    .B1(_11385_),
    .Y(_11386_));
 sky130_fd_sc_hd__a21boi_2 _33423_ (.A1(_10970_),
    .A2(_10984_),
    .B1_N(_10980_),
    .Y(_11387_));
 sky130_fd_sc_hd__a21o_2 _33424_ (.A1(_11376_),
    .A2(_11379_),
    .B1(_11380_),
    .X(_11388_));
 sky130_fd_sc_hd__nand3_2 _33425_ (.A(_11376_),
    .B(_11379_),
    .C(_11380_),
    .Y(_11389_));
 sky130_fd_sc_hd__nand3_2 _33426_ (.A(_11388_),
    .B(_11389_),
    .C(_11384_),
    .Y(_11390_));
 sky130_fd_sc_hd__nand3_2 _33427_ (.A(_11386_),
    .B(_11387_),
    .C(_11390_),
    .Y(_11391_));
 sky130_fd_sc_hd__o21ai_2 _33428_ (.A1(_11381_),
    .A2(_11383_),
    .B1(_11384_),
    .Y(_11392_));
 sky130_fd_sc_hd__nand3_2 _33429_ (.A(_11388_),
    .B(_11389_),
    .C(_11385_),
    .Y(_11393_));
 sky130_fd_sc_hd__nand2_2 _33430_ (.A(_10970_),
    .B(_10984_),
    .Y(_11394_));
 sky130_fd_sc_hd__nand2_2 _33431_ (.A(_11394_),
    .B(_10980_),
    .Y(_11395_));
 sky130_fd_sc_hd__nand3_2 _33432_ (.A(_11392_),
    .B(_11393_),
    .C(_11395_),
    .Y(_11396_));
 sky130_fd_sc_hd__nand2_2 _33433_ (.A(_11391_),
    .B(_11396_),
    .Y(_11397_));
 sky130_fd_sc_hd__nand2_2 _33434_ (.A(_11077_),
    .B(_11064_),
    .Y(_11398_));
 sky130_fd_sc_hd__nand2_2 _33435_ (.A(_11397_),
    .B(_11398_),
    .Y(_11399_));
 sky130_fd_sc_hd__nand2_2 _33436_ (.A(_11083_),
    .B(_11080_),
    .Y(_11400_));
 sky130_fd_sc_hd__nand2_2 _33437_ (.A(_11400_),
    .B(_11082_),
    .Y(_11401_));
 sky130_fd_sc_hd__a21oi_2 _33438_ (.A1(_11068_),
    .A2(_11071_),
    .B1(_11076_),
    .Y(_11402_));
 sky130_fd_sc_hd__nand3_2 _33439_ (.A(_11391_),
    .B(_11396_),
    .C(_11402_),
    .Y(_11403_));
 sky130_fd_sc_hd__nand3_2 _33440_ (.A(_11399_),
    .B(_11401_),
    .C(_11403_),
    .Y(_11404_));
 sky130_fd_sc_hd__nand2_2 _33441_ (.A(_11397_),
    .B(_11402_),
    .Y(_11405_));
 sky130_fd_sc_hd__o21ai_2 _33442_ (.A1(_11080_),
    .A2(_11075_),
    .B1(_11083_),
    .Y(_11406_));
 sky130_fd_sc_hd__nand3_2 _33443_ (.A(_11391_),
    .B(_11396_),
    .C(_11398_),
    .Y(_11407_));
 sky130_fd_sc_hd__nand3_2 _33444_ (.A(_11405_),
    .B(_11406_),
    .C(_11407_),
    .Y(_11408_));
 sky130_fd_sc_hd__nand2_2 _33445_ (.A(_11404_),
    .B(_11408_),
    .Y(_11409_));
 sky130_fd_sc_hd__buf_1 _33446_ (.A(\pcpi_mul.rs1[28] ),
    .X(_11410_));
 sky130_fd_sc_hd__nand2_2 _33447_ (.A(_06199_),
    .B(_11410_),
    .Y(_11411_));
 sky130_fd_sc_hd__nand2_2 _33448_ (.A(_06201_),
    .B(_10538_),
    .Y(_11412_));
 sky130_fd_sc_hd__nor2_2 _33449_ (.A(_11411_),
    .B(_11412_),
    .Y(_11413_));
 sky130_fd_sc_hd__nand2_2 _33450_ (.A(_11411_),
    .B(_11412_),
    .Y(_11414_));
 sky130_fd_sc_hd__inv_2 _33451_ (.A(_11414_),
    .Y(_11415_));
 sky130_fd_sc_hd__o21ai_2 _33452_ (.A1(_11413_),
    .A2(_11415_),
    .B1(_11030_),
    .Y(_11416_));
 sky130_fd_sc_hd__or2_2 _33453_ (.A(_11411_),
    .B(_11412_),
    .X(_11417_));
 sky130_fd_sc_hd__buf_1 _33454_ (.A(_11025_),
    .X(_11418_));
 sky130_fd_sc_hd__nand3_2 _33455_ (.A(_11417_),
    .B(_11418_),
    .C(_11414_),
    .Y(_11419_));
 sky130_fd_sc_hd__a21o_2 _33456_ (.A1(_11418_),
    .A2(_11022_),
    .B1(_11020_),
    .X(_11420_));
 sky130_fd_sc_hd__nand3_2 _33457_ (.A(_11416_),
    .B(_11419_),
    .C(_11420_),
    .Y(_11421_));
 sky130_fd_sc_hd__o21ai_2 _33458_ (.A1(_11413_),
    .A2(_11415_),
    .B1(_11026_),
    .Y(_11422_));
 sky130_fd_sc_hd__nand3_2 _33459_ (.A(_11417_),
    .B(_11029_),
    .C(_11414_),
    .Y(_11423_));
 sky130_fd_sc_hd__a21oi_2 _33460_ (.A1(_11026_),
    .A2(_11022_),
    .B1(_11020_),
    .Y(_11424_));
 sky130_fd_sc_hd__nand3_2 _33461_ (.A(_11422_),
    .B(_11423_),
    .C(_11424_),
    .Y(_11425_));
 sky130_fd_sc_hd__nand2_2 _33462_ (.A(_11421_),
    .B(_11425_),
    .Y(_11426_));
 sky130_fd_sc_hd__buf_1 _33463_ (.A(\pcpi_mul.rs1[31] ),
    .X(_11427_));
 sky130_fd_sc_hd__nand2_2 _33464_ (.A(_06072_),
    .B(_11427_),
    .Y(_11428_));
 sky130_fd_sc_hd__buf_1 _33465_ (.A(_11023_),
    .X(_11429_));
 sky130_fd_sc_hd__nand2_2 _33466_ (.A(_11429_),
    .B(_05118_),
    .Y(_11430_));
 sky130_fd_sc_hd__nor2_2 _33467_ (.A(_11428_),
    .B(_11430_),
    .Y(_11431_));
 sky130_fd_sc_hd__nand2_2 _33468_ (.A(_11428_),
    .B(_11430_),
    .Y(_11432_));
 sky130_fd_sc_hd__inv_2 _33469_ (.A(_11432_),
    .Y(_11433_));
 sky130_fd_sc_hd__nor2_2 _33470_ (.A(_05150_),
    .B(_10535_),
    .Y(_11434_));
 sky130_fd_sc_hd__inv_2 _33471_ (.A(_11434_),
    .Y(_11435_));
 sky130_fd_sc_hd__o21ai_2 _33472_ (.A1(_11431_),
    .A2(_11433_),
    .B1(_11435_),
    .Y(_11436_));
 sky130_fd_sc_hd__nand3b_2 _33473_ (.A_N(_11431_),
    .B(_11434_),
    .C(_11432_),
    .Y(_11437_));
 sky130_fd_sc_hd__nand2_2 _33474_ (.A(_11436_),
    .B(_11437_),
    .Y(_11438_));
 sky130_fd_sc_hd__nand2_2 _33475_ (.A(_11426_),
    .B(_11438_),
    .Y(_11439_));
 sky130_fd_sc_hd__nand3b_2 _33476_ (.A_N(_11438_),
    .B(_11421_),
    .C(_11425_),
    .Y(_11440_));
 sky130_fd_sc_hd__nand2_2 _33477_ (.A(_11035_),
    .B(_11045_),
    .Y(_11441_));
 sky130_fd_sc_hd__nand2_2 _33478_ (.A(_11441_),
    .B(_11032_),
    .Y(_11442_));
 sky130_fd_sc_hd__a21oi_2 _33479_ (.A1(_11439_),
    .A2(_11440_),
    .B1(_11442_),
    .Y(_11443_));
 sky130_fd_sc_hd__nand3_2 _33480_ (.A(_11439_),
    .B(_11442_),
    .C(_11440_),
    .Y(_11444_));
 sky130_fd_sc_hd__a21o_2 _33481_ (.A1(_11041_),
    .A2(_11043_),
    .B1(_11040_),
    .X(_11445_));
 sky130_fd_sc_hd__nand2_2 _33482_ (.A(_11444_),
    .B(_11445_),
    .Y(_11446_));
 sky130_fd_sc_hd__nor2_2 _33483_ (.A(_11443_),
    .B(_11446_),
    .Y(_11447_));
 sky130_fd_sc_hd__a21o_2 _33484_ (.A1(_11439_),
    .A2(_11440_),
    .B1(_11442_),
    .X(_11448_));
 sky130_fd_sc_hd__a21oi_2 _33485_ (.A1(_11448_),
    .A2(_11444_),
    .B1(_11445_),
    .Y(_11449_));
 sky130_fd_sc_hd__nor2_2 _33486_ (.A(_11447_),
    .B(_11449_),
    .Y(_11450_));
 sky130_fd_sc_hd__nand2_2 _33487_ (.A(_11409_),
    .B(_11450_),
    .Y(_11451_));
 sky130_fd_sc_hd__a21oi_2 _33488_ (.A1(_10994_),
    .A2(_10995_),
    .B1(_10996_),
    .Y(_11452_));
 sky130_fd_sc_hd__a21oi_2 _33489_ (.A1(_10999_),
    .A2(_11000_),
    .B1(_11452_),
    .Y(_11453_));
 sky130_fd_sc_hd__o211ai_2 _33490_ (.A1(_11447_),
    .A2(_11449_),
    .B1(_11404_),
    .C1(_11408_),
    .Y(_11454_));
 sky130_fd_sc_hd__nand3_2 _33491_ (.A(_11451_),
    .B(_11453_),
    .C(_11454_),
    .Y(_11455_));
 sky130_fd_sc_hd__nand3_2 _33492_ (.A(_11450_),
    .B(_11404_),
    .C(_11408_),
    .Y(_11456_));
 sky130_fd_sc_hd__o2bb2ai_2 _33493_ (.A1_N(_11408_),
    .A2_N(_11404_),
    .B1(_11447_),
    .B2(_11449_),
    .Y(_11457_));
 sky130_fd_sc_hd__o211ai_2 _33494_ (.A1(_11452_),
    .A2(_10998_),
    .B1(_11456_),
    .C1(_11457_),
    .Y(_11458_));
 sky130_fd_sc_hd__nand2_2 _33495_ (.A(_11093_),
    .B(_11092_),
    .Y(_11459_));
 sky130_fd_sc_hd__a21oi_2 _33496_ (.A1(_11455_),
    .A2(_11458_),
    .B1(_11459_),
    .Y(_11460_));
 sky130_fd_sc_hd__nand2_2 _33497_ (.A(_11455_),
    .B(_11459_),
    .Y(_11461_));
 sky130_fd_sc_hd__inv_2 _33498_ (.A(_11458_),
    .Y(_11462_));
 sky130_fd_sc_hd__nor2_2 _33499_ (.A(_11461_),
    .B(_11462_),
    .Y(_11463_));
 sky130_fd_sc_hd__o2bb2ai_2 _33500_ (.A1_N(_11362_),
    .A2_N(_11369_),
    .B1(_11460_),
    .B2(_11463_),
    .Y(_11464_));
 sky130_fd_sc_hd__a32oi_2 _33501_ (.A1(_11451_),
    .A2(_11453_),
    .A3(_11454_),
    .B1(_11092_),
    .B2(_11093_),
    .Y(_11465_));
 sky130_fd_sc_hd__a21oi_2 _33502_ (.A1(_11458_),
    .A2(_11465_),
    .B1(_11460_),
    .Y(_11466_));
 sky130_fd_sc_hd__nand3_2 _33503_ (.A(_11466_),
    .B(_11369_),
    .C(_11362_),
    .Y(_11467_));
 sky130_fd_sc_hd__nand3_2 _33504_ (.A(_11161_),
    .B(_11464_),
    .C(_11467_),
    .Y(_11468_));
 sky130_fd_sc_hd__a21oi_2 _33505_ (.A1(_11012_),
    .A2(_11014_),
    .B1(_11013_),
    .Y(_11469_));
 sky130_fd_sc_hd__a31oi_2 _33506_ (.A1(_11015_),
    .A2(_11099_),
    .A3(_11103_),
    .B1(_11469_),
    .Y(_11470_));
 sky130_fd_sc_hd__nand2_2 _33507_ (.A(_11369_),
    .B(_11362_),
    .Y(_11471_));
 sky130_fd_sc_hd__nand2_2 _33508_ (.A(_11471_),
    .B(_11466_),
    .Y(_11472_));
 sky130_fd_sc_hd__a21o_2 _33509_ (.A1(_11455_),
    .A2(_11458_),
    .B1(_11459_),
    .X(_11473_));
 sky130_fd_sc_hd__o21ai_2 _33510_ (.A1(_11462_),
    .A2(_11461_),
    .B1(_11473_),
    .Y(_11474_));
 sky130_fd_sc_hd__nand3_2 _33511_ (.A(_11474_),
    .B(_11369_),
    .C(_11362_),
    .Y(_11475_));
 sky130_fd_sc_hd__nand3_2 _33512_ (.A(_11470_),
    .B(_11472_),
    .C(_11475_),
    .Y(_11476_));
 sky130_fd_sc_hd__nand2_2 _33513_ (.A(_11110_),
    .B(_11102_),
    .Y(_11477_));
 sky130_fd_sc_hd__inv_2 _33514_ (.A(_11054_),
    .Y(_11478_));
 sky130_fd_sc_hd__nand2_2 _33515_ (.A(_11478_),
    .B(_11051_),
    .Y(_11479_));
 sky130_fd_sc_hd__nand2_2 _33516_ (.A(_11477_),
    .B(_11479_),
    .Y(_11480_));
 sky130_fd_sc_hd__inv_2 _33517_ (.A(_11480_),
    .Y(_11481_));
 sky130_fd_sc_hd__nor2_2 _33518_ (.A(_11479_),
    .B(_11477_),
    .Y(_11482_));
 sky130_fd_sc_hd__o2bb2ai_2 _33519_ (.A1_N(_11468_),
    .A2_N(_11476_),
    .B1(_11481_),
    .B2(_11482_),
    .Y(_11483_));
 sky130_fd_sc_hd__nor2_2 _33520_ (.A(_11482_),
    .B(_11481_),
    .Y(_11484_));
 sky130_fd_sc_hd__nand3_2 _33521_ (.A(_11484_),
    .B(_11476_),
    .C(_11468_),
    .Y(_11485_));
 sky130_fd_sc_hd__nand2_2 _33522_ (.A(_11116_),
    .B(_11130_),
    .Y(_11486_));
 sky130_fd_sc_hd__nand2_2 _33523_ (.A(_11486_),
    .B(_11112_),
    .Y(_11487_));
 sky130_fd_sc_hd__a21oi_2 _33524_ (.A1(_11483_),
    .A2(_11485_),
    .B1(_11487_),
    .Y(_11488_));
 sky130_fd_sc_hd__and3_2 _33525_ (.A(_11105_),
    .B(_11109_),
    .C(_11111_),
    .X(_11489_));
 sky130_fd_sc_hd__o21ai_2 _33526_ (.A1(_11126_),
    .A2(_11158_),
    .B1(_18184_),
    .Y(_11490_));
 sky130_fd_sc_hd__o21ai_2 _33527_ (.A1(_11126_),
    .A2(_11127_),
    .B1(_11490_),
    .Y(_11491_));
 sky130_fd_sc_hd__a31oi_2 _33528_ (.A1(_11113_),
    .A2(_11115_),
    .A3(_11114_),
    .B1(_11491_),
    .Y(_11492_));
 sky130_fd_sc_hd__o211a_2 _33529_ (.A1(_11489_),
    .A2(_11492_),
    .B1(_11485_),
    .C1(_11483_),
    .X(_11493_));
 sky130_fd_sc_hd__o22ai_2 _33530_ (.A1(_11158_),
    .A2(_11159_),
    .B1(_11488_),
    .B2(_11493_),
    .Y(_11494_));
 sky130_fd_sc_hd__a21o_2 _33531_ (.A1(_11483_),
    .A2(_11485_),
    .B1(_11487_),
    .X(_11495_));
 sky130_fd_sc_hd__nand3_2 _33532_ (.A(_11487_),
    .B(_11483_),
    .C(_11485_),
    .Y(_11496_));
 sky130_fd_sc_hd__nand2_2 _33533_ (.A(_11127_),
    .B(_11119_),
    .Y(_11497_));
 sky130_fd_sc_hd__nand3_2 _33534_ (.A(_11495_),
    .B(_11496_),
    .C(_11497_),
    .Y(_11498_));
 sky130_fd_sc_hd__a21oi_2 _33535_ (.A1(_11129_),
    .A2(_11131_),
    .B1(_11132_),
    .Y(_11499_));
 sky130_fd_sc_hd__o21ai_2 _33536_ (.A1(_11135_),
    .A2(_11499_),
    .B1(_11134_),
    .Y(_11500_));
 sky130_fd_sc_hd__a21oi_2 _33537_ (.A1(_11494_),
    .A2(_11498_),
    .B1(_11500_),
    .Y(_11501_));
 sky130_fd_sc_hd__nand3_2 _33538_ (.A(_11494_),
    .B(_11500_),
    .C(_11498_),
    .Y(_11502_));
 sky130_fd_sc_hd__inv_2 _33539_ (.A(_11502_),
    .Y(_11503_));
 sky130_fd_sc_hd__nor2_2 _33540_ (.A(_11501_),
    .B(_11503_),
    .Y(_11504_));
 sky130_fd_sc_hd__a21bo_2 _33541_ (.A1(_11157_),
    .A2(_11138_),
    .B1_N(_11141_),
    .X(_11505_));
 sky130_fd_sc_hd__xor2_2 _33542_ (.A(_11504_),
    .B(_11505_),
    .X(_02652_));
 sky130_fd_sc_hd__nand2_2 _33543_ (.A(_11174_),
    .B(_11191_),
    .Y(_11506_));
 sky130_fd_sc_hd__nand2_2 _33544_ (.A(_11506_),
    .B(_11177_),
    .Y(_11507_));
 sky130_fd_sc_hd__and4b_2 _33545_ (.A_N(_05323_),
    .B(_10817_),
    .C(_10822_),
    .D(_05271_),
    .X(_11508_));
 sky130_fd_sc_hd__buf_1 _33546_ (.A(_18181_),
    .X(_11509_));
 sky130_fd_sc_hd__o22a_2 _33547_ (.A1(_05215_),
    .A2(_11509_),
    .B1(_11164_),
    .B2(_05320_),
    .X(_11510_));
 sky130_fd_sc_hd__nand2_2 _33548_ (.A(\pcpi_mul.rs2[30] ),
    .B(_05158_),
    .Y(_11511_));
 sky130_fd_sc_hd__inv_2 _33549_ (.A(_11511_),
    .Y(_11512_));
 sky130_fd_sc_hd__o21ai_2 _33550_ (.A1(_11508_),
    .A2(_11510_),
    .B1(_11512_),
    .Y(_11513_));
 sky130_fd_sc_hd__buf_1 _33551_ (.A(\pcpi_mul.rs2[32] ),
    .X(_11514_));
 sky130_fd_sc_hd__a22o_2 _33552_ (.A1(_10699_),
    .A2(_05213_),
    .B1(_05100_),
    .B2(_11514_),
    .X(_11515_));
 sky130_fd_sc_hd__nand3b_2 _33553_ (.A_N(_11508_),
    .B(_11515_),
    .C(_11511_),
    .Y(_11516_));
 sky130_fd_sc_hd__a21oi_2 _33554_ (.A1(_11170_),
    .A2(_11167_),
    .B1(_11163_),
    .Y(_11517_));
 sky130_fd_sc_hd__nand3_2 _33555_ (.A(_11513_),
    .B(_11516_),
    .C(_11517_),
    .Y(_11518_));
 sky130_fd_sc_hd__o21ai_2 _33556_ (.A1(_11508_),
    .A2(_11510_),
    .B1(_11511_),
    .Y(_11519_));
 sky130_fd_sc_hd__o21bai_2 _33557_ (.A1(_11166_),
    .A2(_11165_),
    .B1_N(_11163_),
    .Y(_11520_));
 sky130_fd_sc_hd__nand3b_2 _33558_ (.A_N(_11508_),
    .B(_11515_),
    .C(_11512_),
    .Y(_11521_));
 sky130_fd_sc_hd__nand3_2 _33559_ (.A(_11519_),
    .B(_11520_),
    .C(_11521_),
    .Y(_11522_));
 sky130_fd_sc_hd__nor2_2 _33560_ (.A(_09356_),
    .B(_06332_),
    .Y(_11523_));
 sky130_fd_sc_hd__a22oi_2 _33561_ (.A1(_09842_),
    .A2(_06502_),
    .B1(_10136_),
    .B2(_06614_),
    .Y(_11524_));
 sky130_fd_sc_hd__and4_2 _33562_ (.A(_19315_),
    .B(_19319_),
    .C(_19622_),
    .D(_19625_),
    .X(_11525_));
 sky130_fd_sc_hd__nor2_2 _33563_ (.A(_11524_),
    .B(_11525_),
    .Y(_11526_));
 sky130_fd_sc_hd__nor2_2 _33564_ (.A(_11523_),
    .B(_11526_),
    .Y(_11527_));
 sky130_fd_sc_hd__inv_2 _33565_ (.A(_11523_),
    .Y(_11528_));
 sky130_fd_sc_hd__inv_2 _33566_ (.A(_11526_),
    .Y(_11529_));
 sky130_fd_sc_hd__nor2_2 _33567_ (.A(_11528_),
    .B(_11529_),
    .Y(_11530_));
 sky130_fd_sc_hd__o2bb2ai_2 _33568_ (.A1_N(_11518_),
    .A2_N(_11522_),
    .B1(_11527_),
    .B2(_11530_),
    .Y(_11531_));
 sky130_fd_sc_hd__nand2_2 _33569_ (.A(_11526_),
    .B(_11528_),
    .Y(_11532_));
 sky130_fd_sc_hd__o21ai_2 _33570_ (.A1(_11524_),
    .A2(_11525_),
    .B1(_11523_),
    .Y(_11533_));
 sky130_fd_sc_hd__nand2_2 _33571_ (.A(_11532_),
    .B(_11533_),
    .Y(_11534_));
 sky130_fd_sc_hd__nand3_2 _33572_ (.A(_11522_),
    .B(_11518_),
    .C(_11534_),
    .Y(_11535_));
 sky130_fd_sc_hd__nand3_2 _33573_ (.A(_11507_),
    .B(_11531_),
    .C(_11535_),
    .Y(_11536_));
 sky130_fd_sc_hd__a21boi_2 _33574_ (.A1(_11191_),
    .A2(_11174_),
    .B1_N(_11177_),
    .Y(_11537_));
 sky130_fd_sc_hd__inv_2 _33575_ (.A(_11533_),
    .Y(_11538_));
 sky130_fd_sc_hd__inv_2 _33576_ (.A(_11532_),
    .Y(_11539_));
 sky130_fd_sc_hd__o2bb2ai_2 _33577_ (.A1_N(_11518_),
    .A2_N(_11522_),
    .B1(_11538_),
    .B2(_11539_),
    .Y(_11540_));
 sky130_fd_sc_hd__nand3b_2 _33578_ (.A_N(_11534_),
    .B(_11522_),
    .C(_11518_),
    .Y(_11541_));
 sky130_fd_sc_hd__nand3_2 _33579_ (.A(_11537_),
    .B(_11540_),
    .C(_11541_),
    .Y(_11542_));
 sky130_fd_sc_hd__nor2_2 _33580_ (.A(_07651_),
    .B(_11178_),
    .Y(_11543_));
 sky130_fd_sc_hd__a21o_2 _33581_ (.A1(_11181_),
    .A2(_11179_),
    .B1(_11543_),
    .X(_11544_));
 sky130_fd_sc_hd__nand2_2 _33582_ (.A(_09826_),
    .B(_06507_),
    .Y(_11545_));
 sky130_fd_sc_hd__nand2_2 _33583_ (.A(_09827_),
    .B(_05734_),
    .Y(_11546_));
 sky130_fd_sc_hd__nor2_2 _33584_ (.A(_11545_),
    .B(_11546_),
    .Y(_11547_));
 sky130_fd_sc_hd__and2_2 _33585_ (.A(_11545_),
    .B(_11546_),
    .X(_11548_));
 sky130_fd_sc_hd__nand2_2 _33586_ (.A(_10862_),
    .B(_05733_),
    .Y(_11549_));
 sky130_fd_sc_hd__o21ai_2 _33587_ (.A1(_11547_),
    .A2(_11548_),
    .B1(_11549_),
    .Y(_11550_));
 sky130_fd_sc_hd__nand2_2 _33588_ (.A(_11545_),
    .B(_11546_),
    .Y(_11551_));
 sky130_fd_sc_hd__inv_2 _33589_ (.A(_11549_),
    .Y(_11552_));
 sky130_fd_sc_hd__nand3b_2 _33590_ (.A_N(_11547_),
    .B(_11551_),
    .C(_11552_),
    .Y(_11553_));
 sky130_fd_sc_hd__nand3_2 _33591_ (.A(_11544_),
    .B(_11550_),
    .C(_11553_),
    .Y(_11554_));
 sky130_fd_sc_hd__nor2_2 _33592_ (.A(_11203_),
    .B(_11201_),
    .Y(_11555_));
 sky130_fd_sc_hd__nor2_2 _33593_ (.A(_11202_),
    .B(_11555_),
    .Y(_11556_));
 sky130_fd_sc_hd__inv_2 _33594_ (.A(_11556_),
    .Y(_11557_));
 sky130_fd_sc_hd__o21ai_2 _33595_ (.A1(_11547_),
    .A2(_11548_),
    .B1(_11552_),
    .Y(_11558_));
 sky130_fd_sc_hd__nand3b_2 _33596_ (.A_N(_11547_),
    .B(_11551_),
    .C(_11549_),
    .Y(_11559_));
 sky130_fd_sc_hd__a21oi_2 _33597_ (.A1(_11181_),
    .A2(_11179_),
    .B1(_11543_),
    .Y(_11560_));
 sky130_fd_sc_hd__nand3_2 _33598_ (.A(_11558_),
    .B(_11559_),
    .C(_11560_),
    .Y(_11561_));
 sky130_fd_sc_hd__and3_2 _33599_ (.A(_11554_),
    .B(_11557_),
    .C(_11561_),
    .X(_11562_));
 sky130_fd_sc_hd__a21oi_2 _33600_ (.A1(_11554_),
    .A2(_11561_),
    .B1(_11557_),
    .Y(_11563_));
 sky130_fd_sc_hd__o2bb2ai_2 _33601_ (.A1_N(_11536_),
    .A2_N(_11542_),
    .B1(_11562_),
    .B2(_11563_),
    .Y(_11564_));
 sky130_fd_sc_hd__nand2_2 _33602_ (.A(_11193_),
    .B(_11221_),
    .Y(_11565_));
 sky130_fd_sc_hd__nand2_2 _33603_ (.A(_11565_),
    .B(_11199_),
    .Y(_11566_));
 sky130_fd_sc_hd__nor2_2 _33604_ (.A(_11563_),
    .B(_11562_),
    .Y(_11567_));
 sky130_fd_sc_hd__nand3_2 _33605_ (.A(_11542_),
    .B(_11536_),
    .C(_11567_),
    .Y(_11568_));
 sky130_fd_sc_hd__nand3_2 _33606_ (.A(_11564_),
    .B(_11566_),
    .C(_11568_),
    .Y(_11569_));
 sky130_fd_sc_hd__nand2_2 _33607_ (.A(_11542_),
    .B(_11536_),
    .Y(_11570_));
 sky130_fd_sc_hd__nand2_2 _33608_ (.A(_11570_),
    .B(_11567_),
    .Y(_11571_));
 sky130_fd_sc_hd__a21boi_2 _33609_ (.A1(_11221_),
    .A2(_11193_),
    .B1_N(_11199_),
    .Y(_11572_));
 sky130_fd_sc_hd__nand3b_2 _33610_ (.A_N(_11567_),
    .B(_11536_),
    .C(_11542_),
    .Y(_11573_));
 sky130_fd_sc_hd__nand3_2 _33611_ (.A(_11571_),
    .B(_11572_),
    .C(_11573_),
    .Y(_11574_));
 sky130_fd_sc_hd__nand2_2 _33612_ (.A(_09094_),
    .B(_05910_),
    .Y(_11575_));
 sky130_fd_sc_hd__nand2_2 _33613_ (.A(_09614_),
    .B(_07109_),
    .Y(_11576_));
 sky130_fd_sc_hd__nor2_2 _33614_ (.A(_11575_),
    .B(_11576_),
    .Y(_11577_));
 sky130_fd_sc_hd__and2_2 _33615_ (.A(_11575_),
    .B(_11576_),
    .X(_11578_));
 sky130_fd_sc_hd__nand2_2 _33616_ (.A(_08388_),
    .B(_08218_),
    .Y(_11579_));
 sky130_fd_sc_hd__o21ai_2 _33617_ (.A1(_11577_),
    .A2(_11578_),
    .B1(_11579_),
    .Y(_11580_));
 sky130_fd_sc_hd__or2_2 _33618_ (.A(_11575_),
    .B(_11576_),
    .X(_11581_));
 sky130_fd_sc_hd__nand2_2 _33619_ (.A(_11575_),
    .B(_11576_),
    .Y(_11582_));
 sky130_fd_sc_hd__inv_2 _33620_ (.A(_11579_),
    .Y(_11583_));
 sky130_fd_sc_hd__nand3_2 _33621_ (.A(_11581_),
    .B(_11582_),
    .C(_11583_),
    .Y(_11584_));
 sky130_fd_sc_hd__o21ai_2 _33622_ (.A1(_11231_),
    .A2(_11232_),
    .B1(_11237_),
    .Y(_11585_));
 sky130_fd_sc_hd__nand3_2 _33623_ (.A(_11580_),
    .B(_11584_),
    .C(_11585_),
    .Y(_11586_));
 sky130_fd_sc_hd__o21ai_2 _33624_ (.A1(_11577_),
    .A2(_11578_),
    .B1(_11583_),
    .Y(_11587_));
 sky130_fd_sc_hd__nand3_2 _33625_ (.A(_11581_),
    .B(_11582_),
    .C(_11579_),
    .Y(_11588_));
 sky130_fd_sc_hd__a21oi_2 _33626_ (.A1(_11235_),
    .A2(_11236_),
    .B1(_11233_),
    .Y(_11589_));
 sky130_fd_sc_hd__nand3_2 _33627_ (.A(_11587_),
    .B(_11588_),
    .C(_11589_),
    .Y(_11590_));
 sky130_fd_sc_hd__nand2_2 _33628_ (.A(_11586_),
    .B(_11590_),
    .Y(_11591_));
 sky130_fd_sc_hd__nand2_2 _33629_ (.A(_07894_),
    .B(_06206_),
    .Y(_11592_));
 sky130_fd_sc_hd__nand2_2 _33630_ (.A(_07895_),
    .B(_06560_),
    .Y(_11593_));
 sky130_fd_sc_hd__nor2_2 _33631_ (.A(_11592_),
    .B(_11593_),
    .Y(_11594_));
 sky130_fd_sc_hd__nor2_2 _33632_ (.A(_11251_),
    .B(_10268_),
    .Y(_11595_));
 sky130_fd_sc_hd__nand2_2 _33633_ (.A(_11592_),
    .B(_11593_),
    .Y(_11596_));
 sky130_fd_sc_hd__nand2_2 _33634_ (.A(_11595_),
    .B(_11596_),
    .Y(_11597_));
 sky130_fd_sc_hd__and2_2 _33635_ (.A(_11592_),
    .B(_11593_),
    .X(_11598_));
 sky130_fd_sc_hd__o21bai_2 _33636_ (.A1(_11594_),
    .A2(_11598_),
    .B1_N(_11595_),
    .Y(_11599_));
 sky130_fd_sc_hd__o21a_2 _33637_ (.A1(_11594_),
    .A2(_11597_),
    .B1(_11599_),
    .X(_11600_));
 sky130_fd_sc_hd__nand2_2 _33638_ (.A(_11591_),
    .B(_11600_),
    .Y(_11601_));
 sky130_fd_sc_hd__a21boi_2 _33639_ (.A1(_11214_),
    .A2(_11212_),
    .B1_N(_11209_),
    .Y(_11602_));
 sky130_fd_sc_hd__o21ai_2 _33640_ (.A1(_11594_),
    .A2(_11597_),
    .B1(_11599_),
    .Y(_11603_));
 sky130_fd_sc_hd__nand3_2 _33641_ (.A(_11586_),
    .B(_11590_),
    .C(_11603_),
    .Y(_11604_));
 sky130_fd_sc_hd__nand3_2 _33642_ (.A(_11601_),
    .B(_11602_),
    .C(_11604_),
    .Y(_11605_));
 sky130_fd_sc_hd__nand2_2 _33643_ (.A(_11591_),
    .B(_11603_),
    .Y(_11606_));
 sky130_fd_sc_hd__nand2_2 _33644_ (.A(_11212_),
    .B(_11214_),
    .Y(_11607_));
 sky130_fd_sc_hd__nand2_2 _33645_ (.A(_11607_),
    .B(_11209_),
    .Y(_11608_));
 sky130_fd_sc_hd__nand3_2 _33646_ (.A(_11600_),
    .B(_11586_),
    .C(_11590_),
    .Y(_11609_));
 sky130_fd_sc_hd__nand3_2 _33647_ (.A(_11606_),
    .B(_11608_),
    .C(_11609_),
    .Y(_11610_));
 sky130_fd_sc_hd__inv_2 _33648_ (.A(_11245_),
    .Y(_11611_));
 sky130_fd_sc_hd__and3_2 _33649_ (.A(_11241_),
    .B(_11255_),
    .C(_11254_),
    .X(_11612_));
 sky130_fd_sc_hd__o2bb2ai_2 _33650_ (.A1_N(_11605_),
    .A2_N(_11610_),
    .B1(_11611_),
    .B2(_11612_),
    .Y(_11613_));
 sky130_fd_sc_hd__inv_2 _33651_ (.A(_11613_),
    .Y(_11614_));
 sky130_fd_sc_hd__nand2_2 _33652_ (.A(_11256_),
    .B(_11245_),
    .Y(_11615_));
 sky130_fd_sc_hd__nand2_2 _33653_ (.A(_11615_),
    .B(_11241_),
    .Y(_11616_));
 sky130_fd_sc_hd__nand2_2 _33654_ (.A(_11605_),
    .B(_11616_),
    .Y(_11617_));
 sky130_fd_sc_hd__inv_2 _33655_ (.A(_11610_),
    .Y(_11618_));
 sky130_fd_sc_hd__nor2_2 _33656_ (.A(_11617_),
    .B(_11618_),
    .Y(_11619_));
 sky130_fd_sc_hd__o2bb2ai_2 _33657_ (.A1_N(_11569_),
    .A2_N(_11574_),
    .B1(_11614_),
    .B2(_11619_),
    .Y(_11620_));
 sky130_fd_sc_hd__o21a_2 _33658_ (.A1(_11618_),
    .A2(_11617_),
    .B1(_11613_),
    .X(_11621_));
 sky130_fd_sc_hd__nand3_2 _33659_ (.A(_11574_),
    .B(_11621_),
    .C(_11569_),
    .Y(_11622_));
 sky130_fd_sc_hd__a21oi_2 _33660_ (.A1(_11217_),
    .A2(_11222_),
    .B1(_11220_),
    .Y(_11623_));
 sky130_fd_sc_hd__o21ai_2 _33661_ (.A1(_11289_),
    .A2(_11623_),
    .B1(_11224_),
    .Y(_11624_));
 sky130_fd_sc_hd__a21oi_2 _33662_ (.A1(_11620_),
    .A2(_11622_),
    .B1(_11624_),
    .Y(_11625_));
 sky130_fd_sc_hd__nand2_2 _33663_ (.A(_11227_),
    .B(_11229_),
    .Y(_11626_));
 sky130_fd_sc_hd__nand2_2 _33664_ (.A(_11289_),
    .B(_11224_),
    .Y(_11627_));
 sky130_fd_sc_hd__o2111a_2 _33665_ (.A1(_11220_),
    .A2(_11626_),
    .B1(_11622_),
    .C1(_11627_),
    .D1(_11620_),
    .X(_11628_));
 sky130_fd_sc_hd__nand2_2 _33666_ (.A(_06822_),
    .B(_08447_),
    .Y(_11629_));
 sky130_fd_sc_hd__nand2_2 _33667_ (.A(_06828_),
    .B(_19585_),
    .Y(_11630_));
 sky130_fd_sc_hd__nor2_2 _33668_ (.A(_11629_),
    .B(_11630_),
    .Y(_11631_));
 sky130_fd_sc_hd__and2_2 _33669_ (.A(_11629_),
    .B(_11630_),
    .X(_11632_));
 sky130_fd_sc_hd__nand2_2 _33670_ (.A(_09386_),
    .B(_08490_),
    .Y(_11633_));
 sky130_fd_sc_hd__o21ai_2 _33671_ (.A1(_11631_),
    .A2(_11632_),
    .B1(_11633_),
    .Y(_11634_));
 sky130_fd_sc_hd__nand2_2 _33672_ (.A(_11246_),
    .B(_11247_),
    .Y(_11635_));
 sky130_fd_sc_hd__a31o_2 _33673_ (.A1(_11635_),
    .A2(_19353_),
    .A3(_19595_),
    .B1(_11248_),
    .X(_11636_));
 sky130_fd_sc_hd__nand2_2 _33674_ (.A(_11629_),
    .B(_11630_),
    .Y(_11637_));
 sky130_fd_sc_hd__inv_2 _33675_ (.A(_11633_),
    .Y(_11638_));
 sky130_fd_sc_hd__nand3b_2 _33676_ (.A_N(_11631_),
    .B(_11637_),
    .C(_11638_),
    .Y(_11639_));
 sky130_fd_sc_hd__nand3_2 _33677_ (.A(_11634_),
    .B(_11636_),
    .C(_11639_),
    .Y(_11640_));
 sky130_fd_sc_hd__o21ai_2 _33678_ (.A1(_11631_),
    .A2(_11632_),
    .B1(_11638_),
    .Y(_11641_));
 sky130_fd_sc_hd__nand3b_2 _33679_ (.A_N(_11631_),
    .B(_11637_),
    .C(_11633_),
    .Y(_11642_));
 sky130_fd_sc_hd__a21oi_2 _33680_ (.A1(_11252_),
    .A2(_11635_),
    .B1(_11248_),
    .Y(_11643_));
 sky130_fd_sc_hd__nand3_2 _33681_ (.A(_11641_),
    .B(_11642_),
    .C(_11643_),
    .Y(_11644_));
 sky130_fd_sc_hd__a21oi_2 _33682_ (.A1(_11297_),
    .A2(_11298_),
    .B1(_11296_),
    .Y(_11645_));
 sky130_fd_sc_hd__inv_2 _33683_ (.A(_11645_),
    .Y(_11646_));
 sky130_fd_sc_hd__a21o_2 _33684_ (.A1(_11640_),
    .A2(_11644_),
    .B1(_11646_),
    .X(_11647_));
 sky130_fd_sc_hd__nand3_2 _33685_ (.A(_11640_),
    .B(_11644_),
    .C(_11646_),
    .Y(_11648_));
 sky130_fd_sc_hd__o21ai_2 _33686_ (.A1(_11307_),
    .A2(_11305_),
    .B1(_11306_),
    .Y(_11649_));
 sky130_fd_sc_hd__a21oi_2 _33687_ (.A1(_11647_),
    .A2(_11648_),
    .B1(_11649_),
    .Y(_11650_));
 sky130_fd_sc_hd__and3_2 _33688_ (.A(_11647_),
    .B(_11649_),
    .C(_11648_),
    .X(_11651_));
 sky130_fd_sc_hd__a21o_2 _33689_ (.A1(_11331_),
    .A2(_11333_),
    .B1(_11330_),
    .X(_11652_));
 sky130_fd_sc_hd__nand2_2 _33690_ (.A(_06790_),
    .B(_08650_),
    .Y(_11653_));
 sky130_fd_sc_hd__nand2_2 _33691_ (.A(_08320_),
    .B(_07849_),
    .Y(_11654_));
 sky130_fd_sc_hd__nor2_2 _33692_ (.A(_11653_),
    .B(_11654_),
    .Y(_11655_));
 sky130_fd_sc_hd__nand2_2 _33693_ (.A(_11653_),
    .B(_11654_),
    .Y(_11656_));
 sky130_fd_sc_hd__nand2_2 _33694_ (.A(_19368_),
    .B(_19574_),
    .Y(_11657_));
 sky130_fd_sc_hd__inv_2 _33695_ (.A(_11657_),
    .Y(_11658_));
 sky130_fd_sc_hd__nand3b_2 _33696_ (.A_N(_11655_),
    .B(_11656_),
    .C(_11658_),
    .Y(_11659_));
 sky130_fd_sc_hd__buf_1 _33697_ (.A(_09677_),
    .X(_11660_));
 sky130_fd_sc_hd__nand3_2 _33698_ (.A(_19364_),
    .B(_19366_),
    .C(_19581_),
    .Y(_11661_));
 sky130_fd_sc_hd__o21ai_2 _33699_ (.A1(_11660_),
    .A2(_11661_),
    .B1(_11656_),
    .Y(_11662_));
 sky130_fd_sc_hd__nand2_2 _33700_ (.A(_11662_),
    .B(_11657_),
    .Y(_11663_));
 sky130_fd_sc_hd__nand3_2 _33701_ (.A(_11652_),
    .B(_11659_),
    .C(_11663_),
    .Y(_11664_));
 sky130_fd_sc_hd__inv_2 _33702_ (.A(_11664_),
    .Y(_11665_));
 sky130_fd_sc_hd__nand2_2 _33703_ (.A(_06256_),
    .B(_19570_),
    .Y(_11666_));
 sky130_fd_sc_hd__nand2_2 _33704_ (.A(_05670_),
    .B(_19567_),
    .Y(_11667_));
 sky130_fd_sc_hd__nor2_2 _33705_ (.A(_11666_),
    .B(_11667_),
    .Y(_11668_));
 sky130_fd_sc_hd__and2_2 _33706_ (.A(_11666_),
    .B(_11667_),
    .X(_11669_));
 sky130_fd_sc_hd__a211o_2 _33707_ (.A1(_19377_),
    .A2(_19566_),
    .B1(_11668_),
    .C1(_11669_),
    .X(_11670_));
 sky130_fd_sc_hd__inv_2 _33708_ (.A(_08645_),
    .Y(_11671_));
 sky130_fd_sc_hd__nor2_2 _33709_ (.A(_05497_),
    .B(_11671_),
    .Y(_11672_));
 sky130_fd_sc_hd__o21ai_2 _33710_ (.A1(_11668_),
    .A2(_11669_),
    .B1(_11672_),
    .Y(_11673_));
 sky130_fd_sc_hd__nand2_2 _33711_ (.A(_11670_),
    .B(_11673_),
    .Y(_11674_));
 sky130_fd_sc_hd__nand3b_2 _33712_ (.A_N(_11655_),
    .B(_11656_),
    .C(_11657_),
    .Y(_11675_));
 sky130_fd_sc_hd__a21oi_2 _33713_ (.A1(_11331_),
    .A2(_11333_),
    .B1(_11330_),
    .Y(_11676_));
 sky130_fd_sc_hd__nand2_2 _33714_ (.A(_11662_),
    .B(_11658_),
    .Y(_11677_));
 sky130_fd_sc_hd__nand3_2 _33715_ (.A(_11675_),
    .B(_11676_),
    .C(_11677_),
    .Y(_11678_));
 sky130_fd_sc_hd__nand2_2 _33716_ (.A(_11674_),
    .B(_11678_),
    .Y(_11679_));
 sky130_fd_sc_hd__inv_2 _33717_ (.A(_11674_),
    .Y(_11680_));
 sky130_fd_sc_hd__nand2_2 _33718_ (.A(_11664_),
    .B(_11678_),
    .Y(_11681_));
 sky130_fd_sc_hd__nand2_2 _33719_ (.A(_11680_),
    .B(_11681_),
    .Y(_11682_));
 sky130_fd_sc_hd__o21ai_2 _33720_ (.A1(_11665_),
    .A2(_11679_),
    .B1(_11682_),
    .Y(_11683_));
 sky130_fd_sc_hd__o21ai_2 _33721_ (.A1(_11650_),
    .A2(_11651_),
    .B1(_11683_),
    .Y(_11684_));
 sky130_fd_sc_hd__o21ai_2 _33722_ (.A1(_11277_),
    .A2(_11278_),
    .B1(_11263_),
    .Y(_11685_));
 sky130_fd_sc_hd__o21a_2 _33723_ (.A1(_11665_),
    .A2(_11679_),
    .B1(_11682_),
    .X(_11686_));
 sky130_fd_sc_hd__a21o_2 _33724_ (.A1(_11647_),
    .A2(_11648_),
    .B1(_11649_),
    .X(_11687_));
 sky130_fd_sc_hd__nand3_2 _33725_ (.A(_11647_),
    .B(_11649_),
    .C(_11648_),
    .Y(_11688_));
 sky130_fd_sc_hd__nand3_2 _33726_ (.A(_11686_),
    .B(_11687_),
    .C(_11688_),
    .Y(_11689_));
 sky130_fd_sc_hd__nand3_2 _33727_ (.A(_11684_),
    .B(_11685_),
    .C(_11689_),
    .Y(_11690_));
 sky130_fd_sc_hd__a21boi_2 _33728_ (.A1(_11261_),
    .A2(_11265_),
    .B1_N(_11263_),
    .Y(_11691_));
 sky130_fd_sc_hd__o21ai_2 _33729_ (.A1(_11650_),
    .A2(_11651_),
    .B1(_11686_),
    .Y(_11692_));
 sky130_fd_sc_hd__nand3_2 _33730_ (.A(_11687_),
    .B(_11688_),
    .C(_11683_),
    .Y(_11693_));
 sky130_fd_sc_hd__inv_2 _33731_ (.A(_11317_),
    .Y(_11694_));
 sky130_fd_sc_hd__a21oi_2 _33732_ (.A1(_11344_),
    .A2(_11313_),
    .B1(_11694_),
    .Y(_11695_));
 sky130_fd_sc_hd__a31oi_2 _33733_ (.A1(_11691_),
    .A2(_11692_),
    .A3(_11693_),
    .B1(_11695_),
    .Y(_11696_));
 sky130_fd_sc_hd__nand3_2 _33734_ (.A(_11691_),
    .B(_11692_),
    .C(_11693_),
    .Y(_11697_));
 sky130_fd_sc_hd__a21o_2 _33735_ (.A1(_11344_),
    .A2(_11313_),
    .B1(_11694_),
    .X(_11698_));
 sky130_fd_sc_hd__a21oi_2 _33736_ (.A1(_11697_),
    .A2(_11690_),
    .B1(_11698_),
    .Y(_11699_));
 sky130_fd_sc_hd__a21oi_2 _33737_ (.A1(_11690_),
    .A2(_11696_),
    .B1(_11699_),
    .Y(_11700_));
 sky130_fd_sc_hd__o21ai_2 _33738_ (.A1(_11625_),
    .A2(_11628_),
    .B1(_11700_),
    .Y(_11701_));
 sky130_fd_sc_hd__a21boi_2 _33739_ (.A1(_11360_),
    .A2(_11291_),
    .B1_N(_11282_),
    .Y(_11702_));
 sky130_fd_sc_hd__o21a_2 _33740_ (.A1(_11268_),
    .A2(_11267_),
    .B1(_11224_),
    .X(_11703_));
 sky130_fd_sc_hd__o2bb2ai_2 _33741_ (.A1_N(_11622_),
    .A2_N(_11620_),
    .B1(_11623_),
    .B2(_11703_),
    .Y(_11704_));
 sky130_fd_sc_hd__nand3_2 _33742_ (.A(_11624_),
    .B(_11620_),
    .C(_11622_),
    .Y(_11705_));
 sky130_fd_sc_hd__a21o_2 _33743_ (.A1(_11697_),
    .A2(_11690_),
    .B1(_11698_),
    .X(_11706_));
 sky130_fd_sc_hd__nand2_2 _33744_ (.A(_11696_),
    .B(_11690_),
    .Y(_11707_));
 sky130_fd_sc_hd__nand2_2 _33745_ (.A(_11706_),
    .B(_11707_),
    .Y(_11708_));
 sky130_fd_sc_hd__nand3_2 _33746_ (.A(_11704_),
    .B(_11705_),
    .C(_11708_),
    .Y(_11709_));
 sky130_fd_sc_hd__nand3_2 _33747_ (.A(_11701_),
    .B(_11702_),
    .C(_11709_),
    .Y(_11710_));
 sky130_fd_sc_hd__inv_2 _33748_ (.A(_11707_),
    .Y(_11711_));
 sky130_fd_sc_hd__o22ai_2 _33749_ (.A1(_11699_),
    .A2(_11711_),
    .B1(_11625_),
    .B2(_11628_),
    .Y(_11712_));
 sky130_fd_sc_hd__nand3_2 _33750_ (.A(_11704_),
    .B(_11700_),
    .C(_11705_),
    .Y(_11713_));
 sky130_fd_sc_hd__a21oi_2 _33751_ (.A1(_11269_),
    .A2(_11281_),
    .B1(_11276_),
    .Y(_11714_));
 sky130_fd_sc_hd__o21ai_2 _33752_ (.A1(_11367_),
    .A2(_11714_),
    .B1(_11282_),
    .Y(_11715_));
 sky130_fd_sc_hd__nand3_2 _33753_ (.A(_11712_),
    .B(_11713_),
    .C(_11715_),
    .Y(_11716_));
 sky130_fd_sc_hd__nand2_2 _33754_ (.A(_11710_),
    .B(_11716_),
    .Y(_11717_));
 sky130_fd_sc_hd__nand2_2 _33755_ (.A(_11450_),
    .B(_11404_),
    .Y(_11718_));
 sky130_fd_sc_hd__nand2_2 _33756_ (.A(_11718_),
    .B(_11408_),
    .Y(_11719_));
 sky130_fd_sc_hd__inv_2 _33757_ (.A(_11719_),
    .Y(_11720_));
 sky130_fd_sc_hd__a21oi_2 _33758_ (.A1(_11324_),
    .A2(_11326_),
    .B1(_11321_),
    .Y(_11721_));
 sky130_fd_sc_hd__nand2_2 _33759_ (.A(_05857_),
    .B(_19561_),
    .Y(_11722_));
 sky130_fd_sc_hd__nand2_2 _33760_ (.A(_09247_),
    .B(_09203_),
    .Y(_11723_));
 sky130_fd_sc_hd__nor2_2 _33761_ (.A(_11722_),
    .B(_11723_),
    .Y(_11724_));
 sky130_fd_sc_hd__and2_2 _33762_ (.A(_11722_),
    .B(_11723_),
    .X(_11725_));
 sky130_fd_sc_hd__nand2_2 _33763_ (.A(_08953_),
    .B(_09722_),
    .Y(_11726_));
 sky130_fd_sc_hd__o21ai_2 _33764_ (.A1(_11724_),
    .A2(_11725_),
    .B1(_11726_),
    .Y(_11727_));
 sky130_fd_sc_hd__nand2_2 _33765_ (.A(_11722_),
    .B(_11723_),
    .Y(_11728_));
 sky130_fd_sc_hd__inv_2 _33766_ (.A(_11726_),
    .Y(_11729_));
 sky130_fd_sc_hd__nand3b_2 _33767_ (.A_N(_11724_),
    .B(_11728_),
    .C(_11729_),
    .Y(_11730_));
 sky130_fd_sc_hd__nand3b_2 _33768_ (.A_N(_11721_),
    .B(_11727_),
    .C(_11730_),
    .Y(_11731_));
 sky130_fd_sc_hd__o21ai_2 _33769_ (.A1(_11724_),
    .A2(_11725_),
    .B1(_11729_),
    .Y(_11732_));
 sky130_fd_sc_hd__nand3b_2 _33770_ (.A_N(_11724_),
    .B(_11728_),
    .C(_11726_),
    .Y(_11733_));
 sky130_fd_sc_hd__nand3_2 _33771_ (.A(_11732_),
    .B(_11733_),
    .C(_11721_),
    .Y(_11734_));
 sky130_fd_sc_hd__nand2_2 _33772_ (.A(_11379_),
    .B(_11377_),
    .Y(_11735_));
 sky130_fd_sc_hd__a21o_2 _33773_ (.A1(_11731_),
    .A2(_11734_),
    .B1(_11735_),
    .X(_11736_));
 sky130_fd_sc_hd__nand2_2 _33774_ (.A(_11342_),
    .B(_11328_),
    .Y(_11737_));
 sky130_fd_sc_hd__nand2_2 _33775_ (.A(_11737_),
    .B(_11338_),
    .Y(_11738_));
 sky130_fd_sc_hd__nand3_2 _33776_ (.A(_11731_),
    .B(_11734_),
    .C(_11735_),
    .Y(_11739_));
 sky130_fd_sc_hd__nand3_2 _33777_ (.A(_11736_),
    .B(_11738_),
    .C(_11739_),
    .Y(_11740_));
 sky130_fd_sc_hd__a21oi_2 _33778_ (.A1(_11731_),
    .A2(_11734_),
    .B1(_11735_),
    .Y(_11741_));
 sky130_fd_sc_hd__and3_2 _33779_ (.A(_11731_),
    .B(_11734_),
    .C(_11735_),
    .X(_11742_));
 sky130_fd_sc_hd__o21bai_2 _33780_ (.A1(_11741_),
    .A2(_11742_),
    .B1_N(_11738_),
    .Y(_11743_));
 sky130_fd_sc_hd__nor2_2 _33781_ (.A(_11385_),
    .B(_11383_),
    .Y(_11744_));
 sky130_fd_sc_hd__o2bb2ai_2 _33782_ (.A1_N(_11740_),
    .A2_N(_11743_),
    .B1(_11381_),
    .B2(_11744_),
    .Y(_11745_));
 sky130_fd_sc_hd__nor2_2 _33783_ (.A(_11381_),
    .B(_11744_),
    .Y(_11746_));
 sky130_fd_sc_hd__nand3_2 _33784_ (.A(_11743_),
    .B(_11740_),
    .C(_11746_),
    .Y(_11747_));
 sky130_fd_sc_hd__nand2_2 _33785_ (.A(_11391_),
    .B(_11398_),
    .Y(_11748_));
 sky130_fd_sc_hd__nand2_2 _33786_ (.A(_11748_),
    .B(_11396_),
    .Y(_11749_));
 sky130_fd_sc_hd__a21oi_2 _33787_ (.A1(_11745_),
    .A2(_11747_),
    .B1(_11749_),
    .Y(_11750_));
 sky130_fd_sc_hd__a21oi_2 _33788_ (.A1(_11743_),
    .A2(_11740_),
    .B1(_11746_),
    .Y(_11751_));
 sky130_fd_sc_hd__a21oi_2 _33789_ (.A1(_11386_),
    .A2(_11390_),
    .B1(_11387_),
    .Y(_11752_));
 sky130_fd_sc_hd__a31oi_2 _33790_ (.A1(_11386_),
    .A2(_11387_),
    .A3(_11390_),
    .B1(_11402_),
    .Y(_11753_));
 sky130_fd_sc_hd__o21ai_2 _33791_ (.A1(_11752_),
    .A2(_11753_),
    .B1(_11747_),
    .Y(_11754_));
 sky130_fd_sc_hd__nor2_2 _33792_ (.A(_11751_),
    .B(_11754_),
    .Y(_11755_));
 sky130_fd_sc_hd__nand2_2 _33793_ (.A(_11422_),
    .B(_11423_),
    .Y(_11756_));
 sky130_fd_sc_hd__nand2_2 _33794_ (.A(_11421_),
    .B(_11438_),
    .Y(_11757_));
 sky130_fd_sc_hd__nand2_2 _33795_ (.A(_19395_),
    .B(_19542_),
    .Y(_11758_));
 sky130_fd_sc_hd__buf_1 _33796_ (.A(\pcpi_mul.rs1[32] ),
    .X(_11759_));
 sky130_fd_sc_hd__o21ai_2 _33797_ (.A1(_19397_),
    .A2(_05142_),
    .B1(_11759_),
    .Y(_11760_));
 sky130_fd_sc_hd__and3_2 _33798_ (.A(\pcpi_mul.rs1[32] ),
    .B(_19397_),
    .C(_05142_),
    .X(_11761_));
 sky130_fd_sc_hd__nor2_2 _33799_ (.A(_11760_),
    .B(_11761_),
    .Y(_11762_));
 sky130_fd_sc_hd__xnor2_2 _33800_ (.A(_11758_),
    .B(_11762_),
    .Y(_11763_));
 sky130_fd_sc_hd__buf_1 _33801_ (.A(_10535_),
    .X(_11764_));
 sky130_fd_sc_hd__buf_1 _33802_ (.A(\pcpi_mul.rs1[29] ),
    .X(_11765_));
 sky130_fd_sc_hd__nand3_2 _33803_ (.A(_06735_),
    .B(_05721_),
    .C(_11765_),
    .Y(_11766_));
 sky130_fd_sc_hd__a22o_2 _33804_ (.A1(_05712_),
    .A2(_19549_),
    .B1(_05892_),
    .B2(_19545_),
    .X(_11767_));
 sky130_fd_sc_hd__o21ai_2 _33805_ (.A1(_11764_),
    .A2(_11766_),
    .B1(_11767_),
    .Y(_11768_));
 sky130_fd_sc_hd__nand2_2 _33806_ (.A(_11768_),
    .B(_11418_),
    .Y(_11769_));
 sky130_fd_sc_hd__nor2_2 _33807_ (.A(_10535_),
    .B(_11766_),
    .Y(_11770_));
 sky130_fd_sc_hd__nand3b_2 _33808_ (.A_N(_11770_),
    .B(_11029_),
    .C(_11767_),
    .Y(_11771_));
 sky130_fd_sc_hd__a21oi_2 _33809_ (.A1(_11418_),
    .A2(_11414_),
    .B1(_11413_),
    .Y(_11772_));
 sky130_fd_sc_hd__nand3_2 _33810_ (.A(_11769_),
    .B(_11771_),
    .C(_11772_),
    .Y(_11773_));
 sky130_fd_sc_hd__nand2_2 _33811_ (.A(_11767_),
    .B(_11418_),
    .Y(_11774_));
 sky130_fd_sc_hd__a21o_2 _33812_ (.A1(_11025_),
    .A2(_11414_),
    .B1(_11413_),
    .X(_11775_));
 sky130_fd_sc_hd__nand2_2 _33813_ (.A(_11768_),
    .B(_11029_),
    .Y(_11776_));
 sky130_fd_sc_hd__o211ai_2 _33814_ (.A1(_11770_),
    .A2(_11774_),
    .B1(_11775_),
    .C1(_11776_),
    .Y(_11777_));
 sky130_fd_sc_hd__nand3_2 _33815_ (.A(_11763_),
    .B(_11773_),
    .C(_11777_),
    .Y(_11778_));
 sky130_fd_sc_hd__nand2_2 _33816_ (.A(_11777_),
    .B(_11773_),
    .Y(_11779_));
 sky130_fd_sc_hd__xor2_2 _33817_ (.A(_11758_),
    .B(_11762_),
    .X(_11780_));
 sky130_fd_sc_hd__nand2_2 _33818_ (.A(_11779_),
    .B(_11780_),
    .Y(_11781_));
 sky130_fd_sc_hd__o2111ai_2 _33819_ (.A1(_11420_),
    .A2(_11756_),
    .B1(_11757_),
    .C1(_11778_),
    .D1(_11781_),
    .Y(_11782_));
 sky130_fd_sc_hd__nand2_2 _33820_ (.A(_11757_),
    .B(_11425_),
    .Y(_11783_));
 sky130_fd_sc_hd__nand2_2 _33821_ (.A(_11779_),
    .B(_11763_),
    .Y(_11784_));
 sky130_fd_sc_hd__nand3_2 _33822_ (.A(_11780_),
    .B(_11773_),
    .C(_11777_),
    .Y(_11785_));
 sky130_fd_sc_hd__nand3_2 _33823_ (.A(_11783_),
    .B(_11784_),
    .C(_11785_),
    .Y(_11786_));
 sky130_fd_sc_hd__inv_2 _33824_ (.A(_11437_),
    .Y(_11787_));
 sky130_fd_sc_hd__nor2_2 _33825_ (.A(_11431_),
    .B(_11787_),
    .Y(_11788_));
 sky130_fd_sc_hd__inv_2 _33826_ (.A(_11788_),
    .Y(_11789_));
 sky130_fd_sc_hd__a21oi_2 _33827_ (.A1(_11782_),
    .A2(_11786_),
    .B1(_11789_),
    .Y(_11790_));
 sky130_fd_sc_hd__and3_2 _33828_ (.A(_11782_),
    .B(_11786_),
    .C(_11789_),
    .X(_11791_));
 sky130_fd_sc_hd__nor2_2 _33829_ (.A(_11790_),
    .B(_11791_),
    .Y(_11792_));
 sky130_fd_sc_hd__o21bai_2 _33830_ (.A1(_11750_),
    .A2(_11755_),
    .B1_N(_11792_),
    .Y(_11793_));
 sky130_fd_sc_hd__and3_2 _33831_ (.A(_11743_),
    .B(_11740_),
    .C(_11746_),
    .X(_11794_));
 sky130_fd_sc_hd__o21bai_2 _33832_ (.A1(_11751_),
    .A2(_11794_),
    .B1_N(_11749_),
    .Y(_11795_));
 sky130_fd_sc_hd__nand3_2 _33833_ (.A(_11749_),
    .B(_11745_),
    .C(_11747_),
    .Y(_11796_));
 sky130_fd_sc_hd__nand3_2 _33834_ (.A(_11795_),
    .B(_11796_),
    .C(_11792_),
    .Y(_11797_));
 sky130_fd_sc_hd__nand2_2 _33835_ (.A(_11350_),
    .B(_11354_),
    .Y(_11798_));
 sky130_fd_sc_hd__a21oi_2 _33836_ (.A1(_11793_),
    .A2(_11797_),
    .B1(_11798_),
    .Y(_11799_));
 sky130_fd_sc_hd__nor2_2 _33837_ (.A(_11720_),
    .B(_11799_),
    .Y(_11800_));
 sky130_fd_sc_hd__nand3_2 _33838_ (.A(_11798_),
    .B(_11793_),
    .C(_11797_),
    .Y(_11801_));
 sky130_fd_sc_hd__a21oi_2 _33839_ (.A1(_11782_),
    .A2(_11786_),
    .B1(_11788_),
    .Y(_11802_));
 sky130_fd_sc_hd__and3_2 _33840_ (.A(_11782_),
    .B(_11786_),
    .C(_11788_),
    .X(_11803_));
 sky130_fd_sc_hd__o22ai_2 _33841_ (.A1(_11802_),
    .A2(_11803_),
    .B1(_11751_),
    .B2(_11754_),
    .Y(_11804_));
 sky130_fd_sc_hd__nor2_2 _33842_ (.A(_11750_),
    .B(_11804_),
    .Y(_11805_));
 sky130_fd_sc_hd__a21oi_2 _33843_ (.A1(_11795_),
    .A2(_11796_),
    .B1(_11792_),
    .Y(_11806_));
 sky130_fd_sc_hd__nor2_2 _33844_ (.A(_11355_),
    .B(_11359_),
    .Y(_11807_));
 sky130_fd_sc_hd__o21ai_2 _33845_ (.A1(_11805_),
    .A2(_11806_),
    .B1(_11807_),
    .Y(_11808_));
 sky130_fd_sc_hd__a21oi_2 _33846_ (.A1(_11808_),
    .A2(_11801_),
    .B1(_11719_),
    .Y(_11809_));
 sky130_fd_sc_hd__a21oi_2 _33847_ (.A1(_11800_),
    .A2(_11801_),
    .B1(_11809_),
    .Y(_11810_));
 sky130_fd_sc_hd__nand2_2 _33848_ (.A(_11717_),
    .B(_11810_),
    .Y(_11811_));
 sky130_fd_sc_hd__a21boi_2 _33849_ (.A1(_11466_),
    .A2(_11369_),
    .B1_N(_11362_),
    .Y(_11812_));
 sky130_fd_sc_hd__o211a_2 _33850_ (.A1(_11359_),
    .A2(_11355_),
    .B1(_11797_),
    .C1(_11793_),
    .X(_11813_));
 sky130_fd_sc_hd__nand2_2 _33851_ (.A(_11808_),
    .B(_11719_),
    .Y(_11814_));
 sky130_fd_sc_hd__o21ai_2 _33852_ (.A1(_11799_),
    .A2(_11813_),
    .B1(_11720_),
    .Y(_11815_));
 sky130_fd_sc_hd__o21ai_2 _33853_ (.A1(_11813_),
    .A2(_11814_),
    .B1(_11815_),
    .Y(_11816_));
 sky130_fd_sc_hd__nand3_2 _33854_ (.A(_11816_),
    .B(_11716_),
    .C(_11710_),
    .Y(_11817_));
 sky130_fd_sc_hd__nand3_2 _33855_ (.A(_11811_),
    .B(_11812_),
    .C(_11817_),
    .Y(_11818_));
 sky130_fd_sc_hd__nor2_2 _33856_ (.A(_11813_),
    .B(_11814_),
    .Y(_11819_));
 sky130_fd_sc_hd__o2bb2ai_2 _33857_ (.A1_N(_11716_),
    .A2_N(_11710_),
    .B1(_11819_),
    .B2(_11809_),
    .Y(_11820_));
 sky130_fd_sc_hd__a21oi_2 _33858_ (.A1(_11358_),
    .A2(_11361_),
    .B1(_11162_),
    .Y(_11821_));
 sky130_fd_sc_hd__o21ai_2 _33859_ (.A1(_11474_),
    .A2(_11821_),
    .B1(_11362_),
    .Y(_11822_));
 sky130_fd_sc_hd__nand3_2 _33860_ (.A(_11810_),
    .B(_11716_),
    .C(_11710_),
    .Y(_11823_));
 sky130_fd_sc_hd__nand3_2 _33861_ (.A(_11820_),
    .B(_11822_),
    .C(_11823_),
    .Y(_11824_));
 sky130_fd_sc_hd__nand2_2 _33862_ (.A(_11448_),
    .B(_11445_),
    .Y(_11825_));
 sky130_fd_sc_hd__and2_2 _33863_ (.A(_11825_),
    .B(_11444_),
    .X(_11826_));
 sky130_fd_sc_hd__and3_2 _33864_ (.A(_11461_),
    .B(_11458_),
    .C(_11826_),
    .X(_11827_));
 sky130_fd_sc_hd__nor2_2 _33865_ (.A(_11462_),
    .B(_11465_),
    .Y(_11828_));
 sky130_fd_sc_hd__nor2_2 _33866_ (.A(_11826_),
    .B(_11828_),
    .Y(_11829_));
 sky130_fd_sc_hd__nor2_2 _33867_ (.A(_11827_),
    .B(_11829_),
    .Y(_11830_));
 sky130_fd_sc_hd__a21oi_2 _33868_ (.A1(_11818_),
    .A2(_11824_),
    .B1(_11830_),
    .Y(_11831_));
 sky130_fd_sc_hd__a21boi_2 _33869_ (.A1(_11484_),
    .A2(_11476_),
    .B1_N(_11468_),
    .Y(_11832_));
 sky130_fd_sc_hd__and3_2 _33870_ (.A(_11818_),
    .B(_11824_),
    .C(_11830_),
    .X(_11833_));
 sky130_fd_sc_hd__nor3_2 _33871_ (.A(_11831_),
    .B(_11832_),
    .C(_11833_),
    .Y(_11834_));
 sky130_fd_sc_hd__o21ai_2 _33872_ (.A1(_11831_),
    .A2(_11833_),
    .B1(_11832_),
    .Y(_11835_));
 sky130_fd_sc_hd__nand2_2 _33873_ (.A(_11835_),
    .B(_11481_),
    .Y(_11836_));
 sky130_fd_sc_hd__nor2_2 _33874_ (.A(_11834_),
    .B(_11836_),
    .Y(_11837_));
 sky130_fd_sc_hd__inv_2 _33875_ (.A(_11479_),
    .Y(_11838_));
 sky130_fd_sc_hd__and2_2 _33876_ (.A(_11110_),
    .B(_11102_),
    .X(_11839_));
 sky130_fd_sc_hd__a21o_2 _33877_ (.A1(_11818_),
    .A2(_11824_),
    .B1(_11830_),
    .X(_11840_));
 sky130_fd_sc_hd__nand3_2 _33878_ (.A(_11818_),
    .B(_11824_),
    .C(_11830_),
    .Y(_11841_));
 sky130_fd_sc_hd__nand2_2 _33879_ (.A(_11484_),
    .B(_11476_),
    .Y(_11842_));
 sky130_fd_sc_hd__nand2_2 _33880_ (.A(_11842_),
    .B(_11468_),
    .Y(_11843_));
 sky130_fd_sc_hd__a21oi_2 _33881_ (.A1(_11840_),
    .A2(_11841_),
    .B1(_11843_),
    .Y(_11844_));
 sky130_fd_sc_hd__o22ai_2 _33882_ (.A1(_11838_),
    .A2(_11839_),
    .B1(_11844_),
    .B2(_11834_),
    .Y(_11845_));
 sky130_fd_sc_hd__inv_2 _33883_ (.A(_11497_),
    .Y(_11846_));
 sky130_fd_sc_hd__o21ai_2 _33884_ (.A1(_11846_),
    .A2(_11488_),
    .B1(_11496_),
    .Y(_11847_));
 sky130_fd_sc_hd__nand2_2 _33885_ (.A(_11845_),
    .B(_11847_),
    .Y(_11848_));
 sky130_fd_sc_hd__o21ai_2 _33886_ (.A1(_11844_),
    .A2(_11834_),
    .B1(_11481_),
    .Y(_11849_));
 sky130_fd_sc_hd__nand3_2 _33887_ (.A(_11840_),
    .B(_11843_),
    .C(_11841_),
    .Y(_11850_));
 sky130_fd_sc_hd__nand3_2 _33888_ (.A(_11835_),
    .B(_11480_),
    .C(_11850_),
    .Y(_11851_));
 sky130_fd_sc_hd__nand3b_2 _33889_ (.A_N(_11847_),
    .B(_11849_),
    .C(_11851_),
    .Y(_11852_));
 sky130_fd_sc_hd__o21a_2 _33890_ (.A1(_11837_),
    .A2(_11848_),
    .B1(_11852_),
    .X(_11853_));
 sky130_fd_sc_hd__a21oi_2 _33891_ (.A1(_11141_),
    .A2(_11502_),
    .B1(_11501_),
    .Y(_11854_));
 sky130_fd_sc_hd__nor3_2 _33892_ (.A(_11501_),
    .B(_11503_),
    .C(_11142_),
    .Y(_11855_));
 sky130_fd_sc_hd__and2_2 _33893_ (.A(_11157_),
    .B(_11855_),
    .X(_11856_));
 sky130_fd_sc_hd__nor2_2 _33894_ (.A(_11854_),
    .B(_11856_),
    .Y(_11857_));
 sky130_fd_sc_hd__xnor2_2 _33895_ (.A(_11853_),
    .B(_11857_),
    .Y(_02653_));
 sky130_fd_sc_hd__inv_2 _33896_ (.A(_11713_),
    .Y(_11858_));
 sky130_fd_sc_hd__nand2_2 _33897_ (.A(_11712_),
    .B(_11715_),
    .Y(_11859_));
 sky130_fd_sc_hd__a21oi_2 _33898_ (.A1(_11712_),
    .A2(_11713_),
    .B1(_11715_),
    .Y(_11860_));
 sky130_fd_sc_hd__o22ai_2 _33899_ (.A1(_11858_),
    .A2(_11859_),
    .B1(_11816_),
    .B2(_11860_),
    .Y(_11861_));
 sky130_fd_sc_hd__nand2_2 _33900_ (.A(_11666_),
    .B(_11667_),
    .Y(_11862_));
 sky130_fd_sc_hd__a21oi_2 _33901_ (.A1(_11672_),
    .A2(_11862_),
    .B1(_11668_),
    .Y(_11863_));
 sky130_fd_sc_hd__nand2_2 _33902_ (.A(_05448_),
    .B(_19557_),
    .Y(_11864_));
 sky130_fd_sc_hd__nand2_2 _33903_ (.A(_05445_),
    .B(_19552_),
    .Y(_11865_));
 sky130_fd_sc_hd__nor2_2 _33904_ (.A(_11864_),
    .B(_11865_),
    .Y(_11866_));
 sky130_fd_sc_hd__nand2_2 _33905_ (.A(_11864_),
    .B(_11865_),
    .Y(_11867_));
 sky130_fd_sc_hd__nand2_2 _33906_ (.A(_05764_),
    .B(_19548_),
    .Y(_11868_));
 sky130_fd_sc_hd__inv_2 _33907_ (.A(_11868_),
    .Y(_11869_));
 sky130_fd_sc_hd__nand3b_2 _33908_ (.A_N(_11866_),
    .B(_11867_),
    .C(_11869_),
    .Y(_11870_));
 sky130_fd_sc_hd__and2_2 _33909_ (.A(_11864_),
    .B(_11865_),
    .X(_11871_));
 sky130_fd_sc_hd__o21ai_2 _33910_ (.A1(_11866_),
    .A2(_11871_),
    .B1(_11868_),
    .Y(_11872_));
 sky130_fd_sc_hd__nand3b_2 _33911_ (.A_N(_11863_),
    .B(_11870_),
    .C(_11872_),
    .Y(_11873_));
 sky130_fd_sc_hd__o21ai_2 _33912_ (.A1(_11866_),
    .A2(_11871_),
    .B1(_11869_),
    .Y(_11874_));
 sky130_fd_sc_hd__nand3b_2 _33913_ (.A_N(_11866_),
    .B(_11867_),
    .C(_11868_),
    .Y(_11875_));
 sky130_fd_sc_hd__nand3_2 _33914_ (.A(_11874_),
    .B(_11875_),
    .C(_11863_),
    .Y(_11876_));
 sky130_fd_sc_hd__nand2_2 _33915_ (.A(_11873_),
    .B(_11876_),
    .Y(_11877_));
 sky130_fd_sc_hd__a21oi_2 _33916_ (.A1(_11729_),
    .A2(_11728_),
    .B1(_11724_),
    .Y(_11878_));
 sky130_fd_sc_hd__nand2_2 _33917_ (.A(_11877_),
    .B(_11878_),
    .Y(_11879_));
 sky130_fd_sc_hd__nand3b_2 _33918_ (.A_N(_11878_),
    .B(_11873_),
    .C(_11876_),
    .Y(_11880_));
 sky130_fd_sc_hd__nand2_2 _33919_ (.A(_11679_),
    .B(_11664_),
    .Y(_11881_));
 sky130_fd_sc_hd__a21oi_2 _33920_ (.A1(_11879_),
    .A2(_11880_),
    .B1(_11881_),
    .Y(_11882_));
 sky130_fd_sc_hd__a21boi_2 _33921_ (.A1(_11673_),
    .A2(_11670_),
    .B1_N(_11678_),
    .Y(_11883_));
 sky130_fd_sc_hd__o211a_2 _33922_ (.A1(_11665_),
    .A2(_11883_),
    .B1(_11880_),
    .C1(_11879_),
    .X(_11884_));
 sky130_fd_sc_hd__nand2_2 _33923_ (.A(_11739_),
    .B(_11731_),
    .Y(_11885_));
 sky130_fd_sc_hd__o21ai_2 _33924_ (.A1(_11882_),
    .A2(_11884_),
    .B1(_11885_),
    .Y(_11886_));
 sky130_fd_sc_hd__a21boi_2 _33925_ (.A1(_11743_),
    .A2(_11746_),
    .B1_N(_11740_),
    .Y(_11887_));
 sky130_fd_sc_hd__a21o_2 _33926_ (.A1(_11879_),
    .A2(_11880_),
    .B1(_11881_),
    .X(_11888_));
 sky130_fd_sc_hd__inv_2 _33927_ (.A(_11885_),
    .Y(_11889_));
 sky130_fd_sc_hd__nand3_2 _33928_ (.A(_11881_),
    .B(_11879_),
    .C(_11880_),
    .Y(_11890_));
 sky130_fd_sc_hd__nand3_2 _33929_ (.A(_11888_),
    .B(_11889_),
    .C(_11890_),
    .Y(_11891_));
 sky130_fd_sc_hd__nand3_2 _33930_ (.A(_11886_),
    .B(_11887_),
    .C(_11891_),
    .Y(_11892_));
 sky130_fd_sc_hd__o21ai_2 _33931_ (.A1(_11882_),
    .A2(_11884_),
    .B1(_11889_),
    .Y(_11893_));
 sky130_fd_sc_hd__nand2_2 _33932_ (.A(_11736_),
    .B(_11738_),
    .Y(_11894_));
 sky130_fd_sc_hd__o2bb2ai_2 _33933_ (.A1_N(_11743_),
    .A2_N(_11746_),
    .B1(_11742_),
    .B2(_11894_),
    .Y(_11895_));
 sky130_fd_sc_hd__nand3_2 _33934_ (.A(_11888_),
    .B(_11885_),
    .C(_11890_),
    .Y(_11896_));
 sky130_fd_sc_hd__nand3_2 _33935_ (.A(_11893_),
    .B(_11895_),
    .C(_11896_),
    .Y(_11897_));
 sky130_fd_sc_hd__nand2_2 _33936_ (.A(_11892_),
    .B(_11897_),
    .Y(_11898_));
 sky130_fd_sc_hd__a21oi_2 _33937_ (.A1(_11767_),
    .A2(_11418_),
    .B1(_11770_),
    .Y(_11899_));
 sky130_fd_sc_hd__nand2_2 _33938_ (.A(_06051_),
    .B(_11037_),
    .Y(_11900_));
 sky130_fd_sc_hd__buf_1 _33939_ (.A(\pcpi_mul.rs1[31] ),
    .X(_11901_));
 sky130_fd_sc_hd__nand2_2 _33940_ (.A(_06054_),
    .B(_11901_),
    .Y(_11902_));
 sky130_fd_sc_hd__nor2_2 _33941_ (.A(_11900_),
    .B(_11902_),
    .Y(_11903_));
 sky130_fd_sc_hd__nand2_2 _33942_ (.A(_11900_),
    .B(_11902_),
    .Y(_11904_));
 sky130_fd_sc_hd__inv_2 _33943_ (.A(_11904_),
    .Y(_11905_));
 sky130_fd_sc_hd__o21ai_2 _33944_ (.A1(_11903_),
    .A2(_11905_),
    .B1(_11030_),
    .Y(_11906_));
 sky130_fd_sc_hd__inv_2 _33945_ (.A(_11903_),
    .Y(_11907_));
 sky130_fd_sc_hd__nand3_2 _33946_ (.A(_11907_),
    .B(_11026_),
    .C(_11904_),
    .Y(_11908_));
 sky130_fd_sc_hd__nand3b_2 _33947_ (.A_N(_11899_),
    .B(_11906_),
    .C(_11908_),
    .Y(_11909_));
 sky130_fd_sc_hd__o21ai_2 _33948_ (.A1(_11903_),
    .A2(_11905_),
    .B1(_11026_),
    .Y(_11910_));
 sky130_fd_sc_hd__nand3_2 _33949_ (.A(_11907_),
    .B(_11030_),
    .C(_11904_),
    .Y(_11911_));
 sky130_fd_sc_hd__nand3_2 _33950_ (.A(_11910_),
    .B(_11911_),
    .C(_11899_),
    .Y(_11912_));
 sky130_fd_sc_hd__inv_2 _33951_ (.A(_18156_),
    .Y(_11913_));
 sky130_fd_sc_hd__nor2_2 _33952_ (.A(_11913_),
    .B(_05150_),
    .Y(_11914_));
 sky130_fd_sc_hd__inv_2 _33953_ (.A(_11761_),
    .Y(_11915_));
 sky130_fd_sc_hd__nor2_2 _33954_ (.A(_05149_),
    .B(_11760_),
    .Y(_11916_));
 sky130_fd_sc_hd__nand2_2 _33955_ (.A(_11915_),
    .B(_11916_),
    .Y(_11917_));
 sky130_fd_sc_hd__o21a_2 _33956_ (.A1(_11762_),
    .A2(_11914_),
    .B1(_11917_),
    .X(_11918_));
 sky130_fd_sc_hd__buf_1 _33957_ (.A(_11918_),
    .X(_11919_));
 sky130_fd_sc_hd__a21o_2 _33958_ (.A1(_11909_),
    .A2(_11912_),
    .B1(_11919_),
    .X(_11920_));
 sky130_fd_sc_hd__nand3_2 _33959_ (.A(_11909_),
    .B(_11912_),
    .C(_11919_),
    .Y(_11921_));
 sky130_fd_sc_hd__a21bo_2 _33960_ (.A1(_11763_),
    .A2(_11773_),
    .B1_N(_11777_),
    .X(_11922_));
 sky130_fd_sc_hd__a21o_2 _33961_ (.A1(_11920_),
    .A2(_11921_),
    .B1(_11922_),
    .X(_11923_));
 sky130_fd_sc_hd__nand3_2 _33962_ (.A(_11922_),
    .B(_11920_),
    .C(_11921_),
    .Y(_11924_));
 sky130_fd_sc_hd__o21a_2 _33963_ (.A1(_11758_),
    .A2(_11760_),
    .B1(_11915_),
    .X(_11925_));
 sky130_fd_sc_hd__inv_2 _33964_ (.A(_11925_),
    .Y(_11926_));
 sky130_fd_sc_hd__a21o_2 _33965_ (.A1(_11923_),
    .A2(_11924_),
    .B1(_11926_),
    .X(_11927_));
 sky130_fd_sc_hd__a21oi_2 _33966_ (.A1(_11920_),
    .A2(_11921_),
    .B1(_11922_),
    .Y(_11928_));
 sky130_fd_sc_hd__nor2_2 _33967_ (.A(_11925_),
    .B(_11928_),
    .Y(_11929_));
 sky130_fd_sc_hd__nand2_2 _33968_ (.A(_11929_),
    .B(_11924_),
    .Y(_11930_));
 sky130_fd_sc_hd__nand2_2 _33969_ (.A(_11927_),
    .B(_11930_),
    .Y(_11931_));
 sky130_fd_sc_hd__nand2_2 _33970_ (.A(_11898_),
    .B(_11931_),
    .Y(_11932_));
 sky130_fd_sc_hd__nand2_2 _33971_ (.A(_11697_),
    .B(_11698_),
    .Y(_11933_));
 sky130_fd_sc_hd__nand2_2 _33972_ (.A(_11933_),
    .B(_11690_),
    .Y(_11934_));
 sky130_fd_sc_hd__a21oi_2 _33973_ (.A1(_11923_),
    .A2(_11924_),
    .B1(_11926_),
    .Y(_11935_));
 sky130_fd_sc_hd__a21oi_2 _33974_ (.A1(_11924_),
    .A2(_11929_),
    .B1(_11935_),
    .Y(_11936_));
 sky130_fd_sc_hd__nand3_2 _33975_ (.A(_11936_),
    .B(_11892_),
    .C(_11897_),
    .Y(_11937_));
 sky130_fd_sc_hd__nand3_2 _33976_ (.A(_11932_),
    .B(_11934_),
    .C(_11937_),
    .Y(_11938_));
 sky130_fd_sc_hd__nand2_2 _33977_ (.A(_11898_),
    .B(_11936_),
    .Y(_11939_));
 sky130_fd_sc_hd__a21boi_2 _33978_ (.A1(_11697_),
    .A2(_11698_),
    .B1_N(_11690_),
    .Y(_11940_));
 sky130_fd_sc_hd__nand3_2 _33979_ (.A(_11931_),
    .B(_11892_),
    .C(_11897_),
    .Y(_11941_));
 sky130_fd_sc_hd__nand3_2 _33980_ (.A(_11939_),
    .B(_11940_),
    .C(_11941_),
    .Y(_11942_));
 sky130_fd_sc_hd__a21oi_2 _33981_ (.A1(_11795_),
    .A2(_11792_),
    .B1(_11755_),
    .Y(_11943_));
 sky130_fd_sc_hd__inv_2 _33982_ (.A(_11943_),
    .Y(_11944_));
 sky130_fd_sc_hd__a21oi_2 _33983_ (.A1(_11938_),
    .A2(_11942_),
    .B1(_11944_),
    .Y(_11945_));
 sky130_fd_sc_hd__nand2_2 _33984_ (.A(_11938_),
    .B(_11942_),
    .Y(_11946_));
 sky130_fd_sc_hd__nor2_2 _33985_ (.A(_11943_),
    .B(_11946_),
    .Y(_11947_));
 sky130_fd_sc_hd__nor2_2 _33986_ (.A(_11945_),
    .B(_11947_),
    .Y(_11948_));
 sky130_fd_sc_hd__nand3_2 _33987_ (.A(\pcpi_mul.rs2[32] ),
    .B(\pcpi_mul.rs2[31] ),
    .C(_05211_),
    .Y(_11949_));
 sky130_fd_sc_hd__nor2_2 _33988_ (.A(_05213_),
    .B(_11949_),
    .Y(_11950_));
 sky130_fd_sc_hd__o22a_2 _33989_ (.A1(_05213_),
    .A2(_18181_),
    .B1(_11164_),
    .B2(_06105_),
    .X(_11951_));
 sky130_fd_sc_hd__nand2_2 _33990_ (.A(\pcpi_mul.rs2[30] ),
    .B(_05340_),
    .Y(_11952_));
 sky130_fd_sc_hd__o21ai_2 _33991_ (.A1(_11950_),
    .A2(_11951_),
    .B1(_11952_),
    .Y(_11953_));
 sky130_fd_sc_hd__o21bai_2 _33992_ (.A1(_11511_),
    .A2(_11510_),
    .B1_N(_11508_),
    .Y(_11954_));
 sky130_fd_sc_hd__a22o_2 _33993_ (.A1(_10699_),
    .A2(_05222_),
    .B1(_05320_),
    .B2(_10818_),
    .X(_11955_));
 sky130_fd_sc_hd__inv_2 _33994_ (.A(_11952_),
    .Y(_11956_));
 sky130_fd_sc_hd__nand3b_2 _33995_ (.A_N(_11950_),
    .B(_11955_),
    .C(_11956_),
    .Y(_11957_));
 sky130_fd_sc_hd__nand3_2 _33996_ (.A(_11953_),
    .B(_11954_),
    .C(_11957_),
    .Y(_11958_));
 sky130_fd_sc_hd__o21ai_2 _33997_ (.A1(_11950_),
    .A2(_11951_),
    .B1(_11956_),
    .Y(_11959_));
 sky130_fd_sc_hd__a21oi_2 _33998_ (.A1(_11515_),
    .A2(_11512_),
    .B1(_11508_),
    .Y(_11960_));
 sky130_fd_sc_hd__nand3b_2 _33999_ (.A_N(_11950_),
    .B(_11955_),
    .C(_11952_),
    .Y(_11961_));
 sky130_fd_sc_hd__nand3_2 _34000_ (.A(_11959_),
    .B(_11960_),
    .C(_11961_),
    .Y(_11962_));
 sky130_fd_sc_hd__nand2_2 _34001_ (.A(_11958_),
    .B(_11962_),
    .Y(_11963_));
 sky130_fd_sc_hd__nor2_2 _34002_ (.A(_06809_),
    .B(_10704_),
    .Y(_11964_));
 sky130_fd_sc_hd__inv_2 _34003_ (.A(_11964_),
    .Y(_11965_));
 sky130_fd_sc_hd__nand2_2 _34004_ (.A(_19322_),
    .B(_19615_),
    .Y(_11966_));
 sky130_fd_sc_hd__a22oi_2 _34005_ (.A1(_10138_),
    .A2(_05422_),
    .B1(_10141_),
    .B2(_19619_),
    .Y(_11967_));
 sky130_fd_sc_hd__nor2_2 _34006_ (.A(_11966_),
    .B(_11967_),
    .Y(_11968_));
 sky130_fd_sc_hd__inv_2 _34007_ (.A(_11966_),
    .Y(_11969_));
 sky130_fd_sc_hd__nor2_2 _34008_ (.A(_11967_),
    .B(_11964_),
    .Y(_11970_));
 sky130_fd_sc_hd__nor2_2 _34009_ (.A(_11969_),
    .B(_11970_),
    .Y(_11971_));
 sky130_fd_sc_hd__a21oi_2 _34010_ (.A1(_11965_),
    .A2(_11968_),
    .B1(_11971_),
    .Y(_11972_));
 sky130_fd_sc_hd__nand2_2 _34011_ (.A(_11963_),
    .B(_11972_),
    .Y(_11973_));
 sky130_fd_sc_hd__a21boi_2 _34012_ (.A1(_11518_),
    .A2(_11534_),
    .B1_N(_11522_),
    .Y(_11974_));
 sky130_fd_sc_hd__a22o_2 _34013_ (.A1(_19315_),
    .A2(_19622_),
    .B1(_09602_),
    .B2(_05426_),
    .X(_11975_));
 sky130_fd_sc_hd__nand2_2 _34014_ (.A(_11965_),
    .B(_11975_),
    .Y(_11976_));
 sky130_fd_sc_hd__nor2_2 _34015_ (.A(_11966_),
    .B(_11976_),
    .Y(_11977_));
 sky130_fd_sc_hd__o211ai_2 _34016_ (.A1(_11971_),
    .A2(_11977_),
    .B1(_11962_),
    .C1(_11958_),
    .Y(_11978_));
 sky130_fd_sc_hd__nand3_2 _34017_ (.A(_11973_),
    .B(_11974_),
    .C(_11978_),
    .Y(_11979_));
 sky130_fd_sc_hd__nand2_2 _34018_ (.A(_11518_),
    .B(_11534_),
    .Y(_11980_));
 sky130_fd_sc_hd__nand2_2 _34019_ (.A(_11980_),
    .B(_11522_),
    .Y(_11981_));
 sky130_fd_sc_hd__o2bb2ai_2 _34020_ (.A1_N(_11962_),
    .A2_N(_11958_),
    .B1(_11971_),
    .B2(_11977_),
    .Y(_11982_));
 sky130_fd_sc_hd__nand3_2 _34021_ (.A(_11972_),
    .B(_11958_),
    .C(_11962_),
    .Y(_11983_));
 sky130_fd_sc_hd__nand3_2 _34022_ (.A(_11981_),
    .B(_11982_),
    .C(_11983_),
    .Y(_11984_));
 sky130_fd_sc_hd__nand2_2 _34023_ (.A(_11979_),
    .B(_11984_),
    .Y(_11985_));
 sky130_fd_sc_hd__nand2_2 _34024_ (.A(\pcpi_mul.rs2[26] ),
    .B(_05516_),
    .Y(_11986_));
 sky130_fd_sc_hd__nand2_2 _34025_ (.A(_19330_),
    .B(_06497_),
    .Y(_11987_));
 sky130_fd_sc_hd__nor2_2 _34026_ (.A(_11986_),
    .B(_11987_),
    .Y(_11988_));
 sky130_fd_sc_hd__and2_2 _34027_ (.A(_11986_),
    .B(_11987_),
    .X(_11989_));
 sky130_fd_sc_hd__nand2_2 _34028_ (.A(_19333_),
    .B(_06369_),
    .Y(_11990_));
 sky130_fd_sc_hd__inv_2 _34029_ (.A(_11990_),
    .Y(_11991_));
 sky130_fd_sc_hd__o21ai_2 _34030_ (.A1(_11988_),
    .A2(_11989_),
    .B1(_11991_),
    .Y(_11992_));
 sky130_fd_sc_hd__nand2_2 _34031_ (.A(_11986_),
    .B(_11987_),
    .Y(_11993_));
 sky130_fd_sc_hd__nand3b_2 _34032_ (.A_N(_11988_),
    .B(_11993_),
    .C(_11990_),
    .Y(_11994_));
 sky130_fd_sc_hd__a22o_2 _34033_ (.A1(_09842_),
    .A2(_05269_),
    .B1(_10141_),
    .B2(_06606_),
    .X(_11995_));
 sky130_fd_sc_hd__a21oi_2 _34034_ (.A1(_11523_),
    .A2(_11995_),
    .B1(_11525_),
    .Y(_11996_));
 sky130_fd_sc_hd__nand3_2 _34035_ (.A(_11992_),
    .B(_11994_),
    .C(_11996_),
    .Y(_11997_));
 sky130_fd_sc_hd__a21o_2 _34036_ (.A1(_11552_),
    .A2(_11551_),
    .B1(_11547_),
    .X(_11998_));
 sky130_fd_sc_hd__and2_2 _34037_ (.A(_11997_),
    .B(_11998_),
    .X(_11999_));
 sky130_fd_sc_hd__nand3b_2 _34038_ (.A_N(_11988_),
    .B(_11993_),
    .C(_11991_),
    .Y(_12000_));
 sky130_fd_sc_hd__o21ai_2 _34039_ (.A1(_11988_),
    .A2(_11989_),
    .B1(_11990_),
    .Y(_12001_));
 sky130_fd_sc_hd__nand3b_2 _34040_ (.A_N(_11996_),
    .B(_12000_),
    .C(_12001_),
    .Y(_12002_));
 sky130_fd_sc_hd__a21oi_2 _34041_ (.A1(_12002_),
    .A2(_11997_),
    .B1(_11998_),
    .Y(_12003_));
 sky130_fd_sc_hd__a21oi_2 _34042_ (.A1(_11999_),
    .A2(_12002_),
    .B1(_12003_),
    .Y(_12004_));
 sky130_fd_sc_hd__nand2_2 _34043_ (.A(_11985_),
    .B(_12004_),
    .Y(_12005_));
 sky130_fd_sc_hd__a21boi_2 _34044_ (.A1(_11542_),
    .A2(_11567_),
    .B1_N(_11536_),
    .Y(_12006_));
 sky130_fd_sc_hd__nand3b_2 _34045_ (.A_N(_12004_),
    .B(_11984_),
    .C(_11979_),
    .Y(_12007_));
 sky130_fd_sc_hd__nand3_2 _34046_ (.A(_12005_),
    .B(_12006_),
    .C(_12007_),
    .Y(_12008_));
 sky130_fd_sc_hd__nand2_2 _34047_ (.A(_11542_),
    .B(_11567_),
    .Y(_12009_));
 sky130_fd_sc_hd__nand2_2 _34048_ (.A(_12009_),
    .B(_11536_),
    .Y(_12010_));
 sky130_fd_sc_hd__and3_2 _34049_ (.A(_12002_),
    .B(_11997_),
    .C(_11998_),
    .X(_12011_));
 sky130_fd_sc_hd__o2bb2ai_2 _34050_ (.A1_N(_11984_),
    .A2_N(_11979_),
    .B1(_12011_),
    .B2(_12003_),
    .Y(_12012_));
 sky130_fd_sc_hd__nand3_2 _34051_ (.A(_11979_),
    .B(_11984_),
    .C(_12004_),
    .Y(_12013_));
 sky130_fd_sc_hd__nand3_2 _34052_ (.A(_12010_),
    .B(_12012_),
    .C(_12013_),
    .Y(_12014_));
 sky130_fd_sc_hd__nand2_2 _34053_ (.A(_12008_),
    .B(_12014_),
    .Y(_12015_));
 sky130_fd_sc_hd__and3_2 _34054_ (.A(_11558_),
    .B(_11559_),
    .C(_11560_),
    .X(_12016_));
 sky130_fd_sc_hd__and2_2 _34055_ (.A(_11554_),
    .B(_11556_),
    .X(_12017_));
 sky130_fd_sc_hd__and4_2 _34056_ (.A(_19336_),
    .B(_19339_),
    .C(_08218_),
    .D(_07109_),
    .X(_12018_));
 sky130_fd_sc_hd__a22o_2 _34057_ (.A1(_08382_),
    .A2(_06538_),
    .B1(_08383_),
    .B2(_06724_),
    .X(_12019_));
 sky130_fd_sc_hd__nand2_2 _34058_ (.A(_19342_),
    .B(_06387_),
    .Y(_12020_));
 sky130_fd_sc_hd__inv_2 _34059_ (.A(_12020_),
    .Y(_12021_));
 sky130_fd_sc_hd__nand3b_2 _34060_ (.A_N(_12018_),
    .B(_12019_),
    .C(_12021_),
    .Y(_12022_));
 sky130_fd_sc_hd__a22oi_2 _34061_ (.A1(_19337_),
    .A2(_06726_),
    .B1(_19340_),
    .B2(_06059_),
    .Y(_12023_));
 sky130_fd_sc_hd__o21ai_2 _34062_ (.A1(_12023_),
    .A2(_12018_),
    .B1(_12020_),
    .Y(_12024_));
 sky130_fd_sc_hd__a21o_2 _34063_ (.A1(_11583_),
    .A2(_11582_),
    .B1(_11577_),
    .X(_12025_));
 sky130_fd_sc_hd__a21o_2 _34064_ (.A1(_12022_),
    .A2(_12024_),
    .B1(_12025_),
    .X(_12026_));
 sky130_fd_sc_hd__nand3_2 _34065_ (.A(_12022_),
    .B(_12025_),
    .C(_12024_),
    .Y(_12027_));
 sky130_fd_sc_hd__and4_2 _34066_ (.A(_07722_),
    .B(_07723_),
    .C(_06949_),
    .D(_06957_),
    .X(_12028_));
 sky130_fd_sc_hd__a22o_2 _34067_ (.A1(_07480_),
    .A2(_19593_),
    .B1(_19349_),
    .B2(_07360_),
    .X(_12029_));
 sky130_fd_sc_hd__inv_2 _34068_ (.A(_12029_),
    .Y(_12030_));
 sky130_fd_sc_hd__nor2_2 _34069_ (.A(_07052_),
    .B(_07832_),
    .Y(_12031_));
 sky130_fd_sc_hd__o21ai_2 _34070_ (.A1(_12028_),
    .A2(_12030_),
    .B1(_12031_),
    .Y(_12032_));
 sky130_fd_sc_hd__inv_2 _34071_ (.A(_12031_),
    .Y(_12033_));
 sky130_fd_sc_hd__nand3b_2 _34072_ (.A_N(_12028_),
    .B(_12033_),
    .C(_12029_),
    .Y(_12034_));
 sky130_fd_sc_hd__nand2_2 _34073_ (.A(_12032_),
    .B(_12034_),
    .Y(_12035_));
 sky130_fd_sc_hd__a21oi_2 _34074_ (.A1(_12026_),
    .A2(_12027_),
    .B1(_12035_),
    .Y(_12036_));
 sky130_fd_sc_hd__nor3_2 _34075_ (.A(_12031_),
    .B(_12028_),
    .C(_12030_),
    .Y(_12037_));
 sky130_fd_sc_hd__o21a_2 _34076_ (.A1(_12028_),
    .A2(_12030_),
    .B1(_12031_),
    .X(_12038_));
 sky130_fd_sc_hd__o211a_2 _34077_ (.A1(_12037_),
    .A2(_12038_),
    .B1(_12027_),
    .C1(_12026_),
    .X(_12039_));
 sky130_fd_sc_hd__o22ai_2 _34078_ (.A1(_12016_),
    .A2(_12017_),
    .B1(_12036_),
    .B2(_12039_),
    .Y(_12040_));
 sky130_fd_sc_hd__a21o_2 _34079_ (.A1(_12026_),
    .A2(_12027_),
    .B1(_12035_),
    .X(_12041_));
 sky130_fd_sc_hd__o21ai_2 _34080_ (.A1(_11556_),
    .A2(_12016_),
    .B1(_11554_),
    .Y(_12042_));
 sky130_fd_sc_hd__nand3_2 _34081_ (.A(_12026_),
    .B(_12035_),
    .C(_12027_),
    .Y(_12043_));
 sky130_fd_sc_hd__nand3_2 _34082_ (.A(_12041_),
    .B(_12042_),
    .C(_12043_),
    .Y(_12044_));
 sky130_fd_sc_hd__inv_2 _34083_ (.A(_11586_),
    .Y(_12045_));
 sky130_fd_sc_hd__a21o_2 _34084_ (.A1(_11590_),
    .A2(_11600_),
    .B1(_12045_),
    .X(_12046_));
 sky130_fd_sc_hd__a21oi_2 _34085_ (.A1(_12040_),
    .A2(_12044_),
    .B1(_12046_),
    .Y(_12047_));
 sky130_fd_sc_hd__and2_2 _34086_ (.A(_11600_),
    .B(_11590_),
    .X(_12048_));
 sky130_fd_sc_hd__o211a_2 _34087_ (.A1(_12045_),
    .A2(_12048_),
    .B1(_12044_),
    .C1(_12040_),
    .X(_12049_));
 sky130_fd_sc_hd__nor2_2 _34088_ (.A(_12047_),
    .B(_12049_),
    .Y(_12050_));
 sky130_fd_sc_hd__nand2_2 _34089_ (.A(_12015_),
    .B(_12050_),
    .Y(_12051_));
 sky130_fd_sc_hd__a21boi_2 _34090_ (.A1(_11574_),
    .A2(_11621_),
    .B1_N(_11569_),
    .Y(_12052_));
 sky130_fd_sc_hd__a21o_2 _34091_ (.A1(_12040_),
    .A2(_12044_),
    .B1(_12046_),
    .X(_12053_));
 sky130_fd_sc_hd__nand3_2 _34092_ (.A(_12040_),
    .B(_12044_),
    .C(_12046_),
    .Y(_12054_));
 sky130_fd_sc_hd__nand2_2 _34093_ (.A(_12053_),
    .B(_12054_),
    .Y(_12055_));
 sky130_fd_sc_hd__nand3_2 _34094_ (.A(_12055_),
    .B(_12014_),
    .C(_12008_),
    .Y(_12056_));
 sky130_fd_sc_hd__nand3_2 _34095_ (.A(_12051_),
    .B(_12052_),
    .C(_12056_),
    .Y(_12057_));
 sky130_fd_sc_hd__nand2_2 _34096_ (.A(_11574_),
    .B(_11621_),
    .Y(_12058_));
 sky130_fd_sc_hd__nand2_2 _34097_ (.A(_12058_),
    .B(_11569_),
    .Y(_12059_));
 sky130_fd_sc_hd__o2bb2ai_2 _34098_ (.A1_N(_12014_),
    .A2_N(_12008_),
    .B1(_12049_),
    .B2(_12047_),
    .Y(_12060_));
 sky130_fd_sc_hd__nand3_2 _34099_ (.A(_12050_),
    .B(_12014_),
    .C(_12008_),
    .Y(_12061_));
 sky130_fd_sc_hd__nand3_2 _34100_ (.A(_12059_),
    .B(_12060_),
    .C(_12061_),
    .Y(_12062_));
 sky130_fd_sc_hd__nand2_2 _34101_ (.A(_07898_),
    .B(_07156_),
    .Y(_12063_));
 sky130_fd_sc_hd__nand2_2 _34102_ (.A(_08345_),
    .B(_07593_),
    .Y(_12064_));
 sky130_fd_sc_hd__nor2_2 _34103_ (.A(_12063_),
    .B(_12064_),
    .Y(_12065_));
 sky130_fd_sc_hd__and2_2 _34104_ (.A(_12063_),
    .B(_12064_),
    .X(_12066_));
 sky130_fd_sc_hd__nand2_2 _34105_ (.A(_09386_),
    .B(_19580_),
    .Y(_12067_));
 sky130_fd_sc_hd__o21ai_2 _34106_ (.A1(_12065_),
    .A2(_12066_),
    .B1(_12067_),
    .Y(_12068_));
 sky130_fd_sc_hd__buf_1 _34107_ (.A(_19352_),
    .X(_12069_));
 sky130_fd_sc_hd__a31o_2 _34108_ (.A1(_11596_),
    .A2(_12069_),
    .A3(_19591_),
    .B1(_11594_),
    .X(_12070_));
 sky130_fd_sc_hd__nand2_2 _34109_ (.A(_12063_),
    .B(_12064_),
    .Y(_12071_));
 sky130_fd_sc_hd__inv_2 _34110_ (.A(_12067_),
    .Y(_12072_));
 sky130_fd_sc_hd__nand3b_2 _34111_ (.A_N(_12065_),
    .B(_12071_),
    .C(_12072_),
    .Y(_12073_));
 sky130_fd_sc_hd__nand3_2 _34112_ (.A(_12068_),
    .B(_12070_),
    .C(_12073_),
    .Y(_12074_));
 sky130_fd_sc_hd__o21ai_2 _34113_ (.A1(_12065_),
    .A2(_12066_),
    .B1(_12072_),
    .Y(_12075_));
 sky130_fd_sc_hd__nand3b_2 _34114_ (.A_N(_12065_),
    .B(_12071_),
    .C(_12067_),
    .Y(_12076_));
 sky130_fd_sc_hd__a21oi_2 _34115_ (.A1(_11595_),
    .A2(_11596_),
    .B1(_11594_),
    .Y(_12077_));
 sky130_fd_sc_hd__nand3_2 _34116_ (.A(_12075_),
    .B(_12076_),
    .C(_12077_),
    .Y(_12078_));
 sky130_fd_sc_hd__a21o_2 _34117_ (.A1(_11638_),
    .A2(_11637_),
    .B1(_11631_),
    .X(_12079_));
 sky130_fd_sc_hd__a21oi_2 _34118_ (.A1(_12074_),
    .A2(_12078_),
    .B1(_12079_),
    .Y(_12080_));
 sky130_fd_sc_hd__and3_2 _34119_ (.A(_12074_),
    .B(_12078_),
    .C(_12079_),
    .X(_12081_));
 sky130_fd_sc_hd__nand2_2 _34120_ (.A(_11644_),
    .B(_11646_),
    .Y(_12082_));
 sky130_fd_sc_hd__nand2_2 _34121_ (.A(_12082_),
    .B(_11640_),
    .Y(_12083_));
 sky130_fd_sc_hd__o21bai_2 _34122_ (.A1(_12080_),
    .A2(_12081_),
    .B1_N(_12083_),
    .Y(_12084_));
 sky130_fd_sc_hd__a21o_2 _34123_ (.A1(_12074_),
    .A2(_12078_),
    .B1(_12079_),
    .X(_12085_));
 sky130_fd_sc_hd__nand3_2 _34124_ (.A(_12074_),
    .B(_12078_),
    .C(_12079_),
    .Y(_12086_));
 sky130_fd_sc_hd__nand3_2 _34125_ (.A(_12085_),
    .B(_12083_),
    .C(_12086_),
    .Y(_12087_));
 sky130_fd_sc_hd__inv_2 _34126_ (.A(\pcpi_mul.rs1[23] ),
    .Y(_12088_));
 sky130_fd_sc_hd__buf_1 _34127_ (.A(_12088_),
    .X(_12089_));
 sky130_fd_sc_hd__buf_1 _34128_ (.A(_12089_),
    .X(_12090_));
 sky130_fd_sc_hd__nand3_2 _34129_ (.A(_06278_),
    .B(_07450_),
    .C(_08497_),
    .Y(_12091_));
 sky130_fd_sc_hd__a22o_2 _34130_ (.A1(_06271_),
    .A2(_19578_),
    .B1(_06273_),
    .B2(_09994_),
    .X(_12092_));
 sky130_fd_sc_hd__o21ai_2 _34131_ (.A1(_09679_),
    .A2(_12091_),
    .B1(_12092_),
    .Y(_12093_));
 sky130_fd_sc_hd__o21ai_2 _34132_ (.A1(_06121_),
    .A2(_12090_),
    .B1(_12093_),
    .Y(_12094_));
 sky130_fd_sc_hd__nor2_2 _34133_ (.A(_11660_),
    .B(_12091_),
    .Y(_12095_));
 sky130_fd_sc_hd__nor2_2 _34134_ (.A(_06119_),
    .B(_12089_),
    .Y(_12096_));
 sky130_fd_sc_hd__nand3b_2 _34135_ (.A_N(_12095_),
    .B(_12092_),
    .C(_12096_),
    .Y(_12097_));
 sky130_fd_sc_hd__a21o_2 _34136_ (.A1(_11658_),
    .A2(_11656_),
    .B1(_11655_),
    .X(_12098_));
 sky130_fd_sc_hd__a21o_2 _34137_ (.A1(_12094_),
    .A2(_12097_),
    .B1(_12098_),
    .X(_12099_));
 sky130_fd_sc_hd__nand3_2 _34138_ (.A(_12094_),
    .B(_12097_),
    .C(_12098_),
    .Y(_12100_));
 sky130_fd_sc_hd__a22oi_2 _34139_ (.A1(_05807_),
    .A2(_08664_),
    .B1(_08331_),
    .B2(_08920_),
    .Y(_12101_));
 sky130_fd_sc_hd__nand2_2 _34140_ (.A(_19376_),
    .B(_19562_),
    .Y(_12102_));
 sky130_fd_sc_hd__inv_2 _34141_ (.A(_12102_),
    .Y(_12103_));
 sky130_fd_sc_hd__nand2_2 _34142_ (.A(_10380_),
    .B(_08664_),
    .Y(_12104_));
 sky130_fd_sc_hd__nor2_2 _34143_ (.A(_06807_),
    .B(_12104_),
    .Y(_12105_));
 sky130_fd_sc_hd__nor3_2 _34144_ (.A(_12101_),
    .B(_12103_),
    .C(_12105_),
    .Y(_12106_));
 sky130_fd_sc_hd__o21a_2 _34145_ (.A1(_12101_),
    .A2(_12105_),
    .B1(_12103_),
    .X(_12107_));
 sky130_fd_sc_hd__nor2_2 _34146_ (.A(_12106_),
    .B(_12107_),
    .Y(_12108_));
 sky130_fd_sc_hd__a21o_2 _34147_ (.A1(_12099_),
    .A2(_12100_),
    .B1(_12108_),
    .X(_12109_));
 sky130_fd_sc_hd__nand3_2 _34148_ (.A(_12099_),
    .B(_12100_),
    .C(_12108_),
    .Y(_12110_));
 sky130_fd_sc_hd__nand2_2 _34149_ (.A(_12109_),
    .B(_12110_),
    .Y(_12111_));
 sky130_fd_sc_hd__a21oi_2 _34150_ (.A1(_12084_),
    .A2(_12087_),
    .B1(_12111_),
    .Y(_12112_));
 sky130_fd_sc_hd__nand2_2 _34151_ (.A(_12085_),
    .B(_12083_),
    .Y(_12113_));
 sky130_fd_sc_hd__o211a_2 _34152_ (.A1(_12081_),
    .A2(_12113_),
    .B1(_12084_),
    .C1(_12111_),
    .X(_12114_));
 sky130_fd_sc_hd__o21ai_2 _34153_ (.A1(_11611_),
    .A2(_11612_),
    .B1(_11610_),
    .Y(_12115_));
 sky130_fd_sc_hd__nand2_2 _34154_ (.A(_12115_),
    .B(_11605_),
    .Y(_12116_));
 sky130_fd_sc_hd__o21ai_2 _34155_ (.A1(_12112_),
    .A2(_12114_),
    .B1(_12116_),
    .Y(_12117_));
 sky130_fd_sc_hd__a21o_2 _34156_ (.A1(_12084_),
    .A2(_12087_),
    .B1(_12111_),
    .X(_12118_));
 sky130_fd_sc_hd__nand3_2 _34157_ (.A(_12111_),
    .B(_12084_),
    .C(_12087_),
    .Y(_12119_));
 sky130_fd_sc_hd__nand2_2 _34158_ (.A(_11617_),
    .B(_11610_),
    .Y(_12120_));
 sky130_fd_sc_hd__nand3_2 _34159_ (.A(_12118_),
    .B(_12119_),
    .C(_12120_),
    .Y(_12121_));
 sky130_fd_sc_hd__o21a_2 _34160_ (.A1(_11683_),
    .A2(_11650_),
    .B1(_11688_),
    .X(_12122_));
 sky130_fd_sc_hd__inv_2 _34161_ (.A(_12122_),
    .Y(_12123_));
 sky130_fd_sc_hd__a21o_2 _34162_ (.A1(_12117_),
    .A2(_12121_),
    .B1(_12123_),
    .X(_12124_));
 sky130_fd_sc_hd__nand3_2 _34163_ (.A(_12117_),
    .B(_12121_),
    .C(_12123_),
    .Y(_12125_));
 sky130_fd_sc_hd__nand2_2 _34164_ (.A(_12124_),
    .B(_12125_),
    .Y(_12126_));
 sky130_fd_sc_hd__a21o_2 _34165_ (.A1(_12057_),
    .A2(_12062_),
    .B1(_12126_),
    .X(_12127_));
 sky130_fd_sc_hd__a21oi_2 _34166_ (.A1(_11704_),
    .A2(_11700_),
    .B1(_11628_),
    .Y(_12128_));
 sky130_fd_sc_hd__nand3_2 _34167_ (.A(_12126_),
    .B(_12062_),
    .C(_12057_),
    .Y(_12129_));
 sky130_fd_sc_hd__nand3_2 _34168_ (.A(_12127_),
    .B(_12128_),
    .C(_12129_),
    .Y(_12130_));
 sky130_fd_sc_hd__o21ai_2 _34169_ (.A1(_11708_),
    .A2(_11625_),
    .B1(_11705_),
    .Y(_12131_));
 sky130_fd_sc_hd__inv_2 _34170_ (.A(_12125_),
    .Y(_12132_));
 sky130_fd_sc_hd__a21oi_2 _34171_ (.A1(_12117_),
    .A2(_12121_),
    .B1(_12123_),
    .Y(_12133_));
 sky130_fd_sc_hd__o2bb2ai_2 _34172_ (.A1_N(_12062_),
    .A2_N(_12057_),
    .B1(_12132_),
    .B2(_12133_),
    .Y(_12134_));
 sky130_fd_sc_hd__nand2_2 _34173_ (.A(_12118_),
    .B(_12119_),
    .Y(_12135_));
 sky130_fd_sc_hd__a21oi_2 _34174_ (.A1(_12135_),
    .A2(_12116_),
    .B1(_12122_),
    .Y(_12136_));
 sky130_fd_sc_hd__a21oi_2 _34175_ (.A1(_12121_),
    .A2(_12136_),
    .B1(_12133_),
    .Y(_12137_));
 sky130_fd_sc_hd__nand3_2 _34176_ (.A(_12137_),
    .B(_12062_),
    .C(_12057_),
    .Y(_12138_));
 sky130_fd_sc_hd__nand3_2 _34177_ (.A(_12131_),
    .B(_12134_),
    .C(_12138_),
    .Y(_12139_));
 sky130_fd_sc_hd__nand3_2 _34178_ (.A(_11948_),
    .B(_12130_),
    .C(_12139_),
    .Y(_12140_));
 sky130_fd_sc_hd__o2bb2ai_2 _34179_ (.A1_N(_12139_),
    .A2_N(_12130_),
    .B1(_11947_),
    .B2(_11945_),
    .Y(_12141_));
 sky130_fd_sc_hd__nand3_2 _34180_ (.A(_11861_),
    .B(_12140_),
    .C(_12141_),
    .Y(_12142_));
 sky130_fd_sc_hd__a21boi_2 _34181_ (.A1(_11810_),
    .A2(_11710_),
    .B1_N(_11716_),
    .Y(_12143_));
 sky130_fd_sc_hd__nand2_2 _34182_ (.A(_11944_),
    .B(_11942_),
    .Y(_12144_));
 sky130_fd_sc_hd__inv_2 _34183_ (.A(_11938_),
    .Y(_12145_));
 sky130_fd_sc_hd__nand2_2 _34184_ (.A(_11946_),
    .B(_11943_),
    .Y(_12146_));
 sky130_fd_sc_hd__o21ai_2 _34185_ (.A1(_12144_),
    .A2(_12145_),
    .B1(_12146_),
    .Y(_12147_));
 sky130_fd_sc_hd__a21o_2 _34186_ (.A1(_12130_),
    .A2(_12139_),
    .B1(_12147_),
    .X(_12148_));
 sky130_fd_sc_hd__nand3_2 _34187_ (.A(_12130_),
    .B(_12147_),
    .C(_12139_),
    .Y(_12149_));
 sky130_fd_sc_hd__nand3_2 _34188_ (.A(_12143_),
    .B(_12148_),
    .C(_12149_),
    .Y(_12150_));
 sky130_fd_sc_hd__and2_2 _34189_ (.A(_11786_),
    .B(_11789_),
    .X(_12151_));
 sky130_fd_sc_hd__inv_2 _34190_ (.A(_12151_),
    .Y(_12152_));
 sky130_fd_sc_hd__nand2_2 _34191_ (.A(_12152_),
    .B(_11782_),
    .Y(_12153_));
 sky130_fd_sc_hd__nand2_2 _34192_ (.A(_11814_),
    .B(_11801_),
    .Y(_12154_));
 sky130_fd_sc_hd__inv_2 _34193_ (.A(_12154_),
    .Y(_12155_));
 sky130_fd_sc_hd__nor2_2 _34194_ (.A(_12153_),
    .B(_12155_),
    .Y(_12156_));
 sky130_fd_sc_hd__inv_2 _34195_ (.A(_12153_),
    .Y(_12157_));
 sky130_fd_sc_hd__nor2_2 _34196_ (.A(_12157_),
    .B(_12154_),
    .Y(_12158_));
 sky130_fd_sc_hd__o2bb2ai_2 _34197_ (.A1_N(_12142_),
    .A2_N(_12150_),
    .B1(_12156_),
    .B2(_12158_),
    .Y(_12159_));
 sky130_fd_sc_hd__a21boi_2 _34198_ (.A1(_11818_),
    .A2(_11830_),
    .B1_N(_11824_),
    .Y(_12160_));
 sky130_fd_sc_hd__nor2_2 _34199_ (.A(_12158_),
    .B(_12156_),
    .Y(_12161_));
 sky130_fd_sc_hd__nand3_2 _34200_ (.A(_12150_),
    .B(_12142_),
    .C(_12161_),
    .Y(_12162_));
 sky130_fd_sc_hd__nand3_2 _34201_ (.A(_12159_),
    .B(_12160_),
    .C(_12162_),
    .Y(_12163_));
 sky130_fd_sc_hd__nor2_2 _34202_ (.A(_12157_),
    .B(_12155_),
    .Y(_12164_));
 sky130_fd_sc_hd__nor2_2 _34203_ (.A(_12153_),
    .B(_12154_),
    .Y(_12165_));
 sky130_fd_sc_hd__o2bb2ai_2 _34204_ (.A1_N(_12142_),
    .A2_N(_12150_),
    .B1(_12164_),
    .B2(_12165_),
    .Y(_12166_));
 sky130_fd_sc_hd__inv_2 _34205_ (.A(_11823_),
    .Y(_12167_));
 sky130_fd_sc_hd__nand2_2 _34206_ (.A(_11820_),
    .B(_11822_),
    .Y(_12168_));
 sky130_fd_sc_hd__o2bb2ai_2 _34207_ (.A1_N(_11830_),
    .A2_N(_11818_),
    .B1(_12167_),
    .B2(_12168_),
    .Y(_12169_));
 sky130_fd_sc_hd__nor2_2 _34208_ (.A(_12165_),
    .B(_12164_),
    .Y(_12170_));
 sky130_fd_sc_hd__nand3_2 _34209_ (.A(_12150_),
    .B(_12142_),
    .C(_12170_),
    .Y(_12171_));
 sky130_fd_sc_hd__nand3_2 _34210_ (.A(_12166_),
    .B(_12169_),
    .C(_12171_),
    .Y(_12172_));
 sky130_fd_sc_hd__nand2_2 _34211_ (.A(_12163_),
    .B(_12172_),
    .Y(_12173_));
 sky130_fd_sc_hd__inv_2 _34212_ (.A(_11829_),
    .Y(_12174_));
 sky130_fd_sc_hd__a22oi_2 _34213_ (.A1(_12173_),
    .A2(_12174_),
    .B1(_11836_),
    .B2(_11850_),
    .Y(_12175_));
 sky130_fd_sc_hd__nand3_2 _34214_ (.A(_12163_),
    .B(_12172_),
    .C(_11829_),
    .Y(_12176_));
 sky130_fd_sc_hd__o2bb2ai_2 _34215_ (.A1_N(_12172_),
    .A2_N(_12163_),
    .B1(_11828_),
    .B2(_11826_),
    .Y(_12177_));
 sky130_fd_sc_hd__nand2_2 _34216_ (.A(_11840_),
    .B(_11843_),
    .Y(_12178_));
 sky130_fd_sc_hd__o22ai_2 _34217_ (.A1(_11833_),
    .A2(_12178_),
    .B1(_11480_),
    .B2(_11844_),
    .Y(_12179_));
 sky130_fd_sc_hd__a21oi_2 _34218_ (.A1(_12177_),
    .A2(_12176_),
    .B1(_12179_),
    .Y(_12180_));
 sky130_fd_sc_hd__a21oi_2 _34219_ (.A1(_12175_),
    .A2(_12176_),
    .B1(_12180_),
    .Y(_12181_));
 sky130_fd_sc_hd__o211ai_2 _34220_ (.A1(_11834_),
    .A2(_11836_),
    .B1(_11847_),
    .C1(_11845_),
    .Y(_12182_));
 sky130_fd_sc_hd__nand2_2 _34221_ (.A(_11857_),
    .B(_12182_),
    .Y(_12183_));
 sky130_fd_sc_hd__nand2_2 _34222_ (.A(_12183_),
    .B(_11852_),
    .Y(_12184_));
 sky130_fd_sc_hd__xnor2_2 _34223_ (.A(_12181_),
    .B(_12184_),
    .Y(_02654_));
 sky130_fd_sc_hd__inv_2 _34224_ (.A(_12176_),
    .Y(_12185_));
 sky130_fd_sc_hd__nand2_2 _34225_ (.A(_12179_),
    .B(_12177_),
    .Y(_12186_));
 sky130_fd_sc_hd__a21o_2 _34226_ (.A1(_12177_),
    .A2(_12176_),
    .B1(_12179_),
    .X(_12187_));
 sky130_fd_sc_hd__o2111a_2 _34227_ (.A1(_12185_),
    .A2(_12186_),
    .B1(_12182_),
    .C1(_11852_),
    .D1(_12187_),
    .X(_12188_));
 sky130_fd_sc_hd__nand2_2 _34228_ (.A(_11856_),
    .B(_12188_),
    .Y(_12189_));
 sky130_fd_sc_hd__nand2_2 _34229_ (.A(_11930_),
    .B(_11924_),
    .Y(_12190_));
 sky130_fd_sc_hd__inv_2 _34230_ (.A(_12190_),
    .Y(_12191_));
 sky130_fd_sc_hd__nand2_2 _34231_ (.A(_12144_),
    .B(_11938_),
    .Y(_12192_));
 sky130_fd_sc_hd__inv_2 _34232_ (.A(_12192_),
    .Y(_12193_));
 sky130_fd_sc_hd__nor2_2 _34233_ (.A(_12191_),
    .B(_12193_),
    .Y(_12194_));
 sky130_fd_sc_hd__nor2_2 _34234_ (.A(_12190_),
    .B(_12192_),
    .Y(_12195_));
 sky130_fd_sc_hd__inv_2 _34235_ (.A(_12061_),
    .Y(_12196_));
 sky130_fd_sc_hd__nand2_2 _34236_ (.A(_12059_),
    .B(_12060_),
    .Y(_12197_));
 sky130_fd_sc_hd__a21oi_2 _34237_ (.A1(_12060_),
    .A2(_12061_),
    .B1(_12059_),
    .Y(_12198_));
 sky130_fd_sc_hd__o22ai_2 _34238_ (.A1(_12196_),
    .A2(_12197_),
    .B1(_12126_),
    .B2(_12198_),
    .Y(_12199_));
 sky130_fd_sc_hd__inv_2 _34239_ (.A(_12013_),
    .Y(_12200_));
 sky130_fd_sc_hd__nand2_2 _34240_ (.A(_12010_),
    .B(_12012_),
    .Y(_12201_));
 sky130_fd_sc_hd__a21oi_2 _34241_ (.A1(_12012_),
    .A2(_12013_),
    .B1(_12010_),
    .Y(_12202_));
 sky130_fd_sc_hd__o22ai_2 _34242_ (.A1(_12200_),
    .A2(_12201_),
    .B1(_12055_),
    .B2(_12202_),
    .Y(_12203_));
 sky130_fd_sc_hd__nand2_2 _34243_ (.A(_11979_),
    .B(_12004_),
    .Y(_12204_));
 sky130_fd_sc_hd__nand2_2 _34244_ (.A(_12204_),
    .B(_11984_),
    .Y(_12205_));
 sky130_fd_sc_hd__inv_2 _34245_ (.A(_11957_),
    .Y(_12206_));
 sky130_fd_sc_hd__nand2_2 _34246_ (.A(_11953_),
    .B(_11954_),
    .Y(_12207_));
 sky130_fd_sc_hd__o2bb2ai_2 _34247_ (.A1_N(_11962_),
    .A2_N(_11972_),
    .B1(_12206_),
    .B2(_12207_),
    .Y(_12208_));
 sky130_fd_sc_hd__nand3_2 _34248_ (.A(_10817_),
    .B(\pcpi_mul.rs2[31] ),
    .C(_05193_),
    .Y(_12209_));
 sky130_fd_sc_hd__nor2_2 _34249_ (.A(_05212_),
    .B(_12209_),
    .Y(_12210_));
 sky130_fd_sc_hd__o22a_2 _34250_ (.A1(_05222_),
    .A2(_18181_),
    .B1(_11164_),
    .B2(_05855_),
    .X(_12211_));
 sky130_fd_sc_hd__nand2_2 _34251_ (.A(\pcpi_mul.rs2[30] ),
    .B(_05342_),
    .Y(_12212_));
 sky130_fd_sc_hd__inv_2 _34252_ (.A(_12212_),
    .Y(_12213_));
 sky130_fd_sc_hd__o21ai_2 _34253_ (.A1(_12210_),
    .A2(_12211_),
    .B1(_12213_),
    .Y(_12214_));
 sky130_fd_sc_hd__a2bb2oi_2 _34254_ (.A1_N(_19631_),
    .A2_N(_11949_),
    .B1(_11956_),
    .B2(_11955_),
    .Y(_12215_));
 sky130_fd_sc_hd__a22o_2 _34255_ (.A1(_19307_),
    .A2(_19625_),
    .B1(_06105_),
    .B2(_11514_),
    .X(_12216_));
 sky130_fd_sc_hd__nand3b_2 _34256_ (.A_N(_12210_),
    .B(_12216_),
    .C(_12212_),
    .Y(_12217_));
 sky130_fd_sc_hd__nand3_2 _34257_ (.A(_12214_),
    .B(_12215_),
    .C(_12217_),
    .Y(_12218_));
 sky130_fd_sc_hd__o21ai_2 _34258_ (.A1(_12210_),
    .A2(_12211_),
    .B1(_12212_),
    .Y(_12219_));
 sky130_fd_sc_hd__o22ai_2 _34259_ (.A1(_06622_),
    .A2(_11949_),
    .B1(_11952_),
    .B2(_11951_),
    .Y(_12220_));
 sky130_fd_sc_hd__nand3b_2 _34260_ (.A_N(_12210_),
    .B(_12216_),
    .C(_12213_),
    .Y(_12221_));
 sky130_fd_sc_hd__nand3_2 _34261_ (.A(_12219_),
    .B(_12220_),
    .C(_12221_),
    .Y(_12222_));
 sky130_fd_sc_hd__nand2_2 _34262_ (.A(_09841_),
    .B(_19618_),
    .Y(_12223_));
 sky130_fd_sc_hd__nand2_2 _34263_ (.A(\pcpi_mul.rs2[28] ),
    .B(_19615_),
    .Y(_12224_));
 sky130_fd_sc_hd__nor2_2 _34264_ (.A(_12223_),
    .B(_12224_),
    .Y(_12225_));
 sky130_fd_sc_hd__and2_2 _34265_ (.A(_12223_),
    .B(_12224_),
    .X(_12226_));
 sky130_fd_sc_hd__nand2_2 _34266_ (.A(_19322_),
    .B(_19613_),
    .Y(_12227_));
 sky130_fd_sc_hd__o21ai_2 _34267_ (.A1(_12225_),
    .A2(_12226_),
    .B1(_12227_),
    .Y(_12228_));
 sky130_fd_sc_hd__inv_2 _34268_ (.A(_12228_),
    .Y(_12229_));
 sky130_fd_sc_hd__inv_2 _34269_ (.A(_12227_),
    .Y(_12230_));
 sky130_fd_sc_hd__nand2_2 _34270_ (.A(_12223_),
    .B(_12224_),
    .Y(_12231_));
 sky130_fd_sc_hd__nand2_2 _34271_ (.A(_12230_),
    .B(_12231_),
    .Y(_12232_));
 sky130_fd_sc_hd__nor2_2 _34272_ (.A(_12225_),
    .B(_12232_),
    .Y(_12233_));
 sky130_fd_sc_hd__o2bb2ai_2 _34273_ (.A1_N(_12218_),
    .A2_N(_12222_),
    .B1(_12229_),
    .B2(_12233_),
    .Y(_12234_));
 sky130_fd_sc_hd__o21a_2 _34274_ (.A1(_12225_),
    .A2(_12232_),
    .B1(_12228_),
    .X(_12235_));
 sky130_fd_sc_hd__nand3_2 _34275_ (.A(_12222_),
    .B(_12218_),
    .C(_12235_),
    .Y(_12236_));
 sky130_fd_sc_hd__nand3_2 _34276_ (.A(_12208_),
    .B(_12234_),
    .C(_12236_),
    .Y(_12237_));
 sky130_fd_sc_hd__nand2_2 _34277_ (.A(_12222_),
    .B(_12218_),
    .Y(_12238_));
 sky130_fd_sc_hd__nand2_2 _34278_ (.A(_12238_),
    .B(_12235_),
    .Y(_12239_));
 sky130_fd_sc_hd__a21boi_2 _34279_ (.A1(_11972_),
    .A2(_11962_),
    .B1_N(_11958_),
    .Y(_12240_));
 sky130_fd_sc_hd__nand3b_2 _34280_ (.A_N(_12235_),
    .B(_12218_),
    .C(_12222_),
    .Y(_12241_));
 sky130_fd_sc_hd__nand3_2 _34281_ (.A(_12239_),
    .B(_12240_),
    .C(_12241_),
    .Y(_12242_));
 sky130_fd_sc_hd__a21oi_2 _34282_ (.A1(_11975_),
    .A2(_11969_),
    .B1(_11964_),
    .Y(_12243_));
 sky130_fd_sc_hd__nand2_2 _34283_ (.A(_09339_),
    .B(_19608_),
    .Y(_12244_));
 sky130_fd_sc_hd__nand2_2 _34284_ (.A(_19330_),
    .B(_06539_),
    .Y(_12245_));
 sky130_fd_sc_hd__nor2_2 _34285_ (.A(_12244_),
    .B(_12245_),
    .Y(_12246_));
 sky130_fd_sc_hd__nand2_2 _34286_ (.A(_12244_),
    .B(_12245_),
    .Y(_12247_));
 sky130_fd_sc_hd__nand2_2 _34287_ (.A(_19333_),
    .B(_06732_),
    .Y(_12248_));
 sky130_fd_sc_hd__inv_2 _34288_ (.A(_12248_),
    .Y(_12249_));
 sky130_fd_sc_hd__nand3b_2 _34289_ (.A_N(_12246_),
    .B(_12247_),
    .C(_12249_),
    .Y(_12250_));
 sky130_fd_sc_hd__and2_2 _34290_ (.A(_12244_),
    .B(_12245_),
    .X(_12251_));
 sky130_fd_sc_hd__o21ai_2 _34291_ (.A1(_12246_),
    .A2(_12251_),
    .B1(_12248_),
    .Y(_12252_));
 sky130_fd_sc_hd__nand3b_2 _34292_ (.A_N(_12243_),
    .B(_12250_),
    .C(_12252_),
    .Y(_12253_));
 sky130_fd_sc_hd__o21ai_2 _34293_ (.A1(_12246_),
    .A2(_12251_),
    .B1(_12249_),
    .Y(_12254_));
 sky130_fd_sc_hd__nand3b_2 _34294_ (.A_N(_12246_),
    .B(_12247_),
    .C(_12248_),
    .Y(_12255_));
 sky130_fd_sc_hd__nand3_2 _34295_ (.A(_12254_),
    .B(_12255_),
    .C(_12243_),
    .Y(_12256_));
 sky130_fd_sc_hd__a21o_2 _34296_ (.A1(_11991_),
    .A2(_11993_),
    .B1(_11988_),
    .X(_12257_));
 sky130_fd_sc_hd__and3_2 _34297_ (.A(_12253_),
    .B(_12256_),
    .C(_12257_),
    .X(_12258_));
 sky130_fd_sc_hd__a21oi_2 _34298_ (.A1(_12253_),
    .A2(_12256_),
    .B1(_12257_),
    .Y(_12259_));
 sky130_fd_sc_hd__o2bb2ai_2 _34299_ (.A1_N(_12237_),
    .A2_N(_12242_),
    .B1(_12258_),
    .B2(_12259_),
    .Y(_12260_));
 sky130_fd_sc_hd__nor2_2 _34300_ (.A(_12259_),
    .B(_12258_),
    .Y(_12261_));
 sky130_fd_sc_hd__nand3_2 _34301_ (.A(_12242_),
    .B(_12237_),
    .C(_12261_),
    .Y(_12262_));
 sky130_fd_sc_hd__nand3_2 _34302_ (.A(_12205_),
    .B(_12260_),
    .C(_12262_),
    .Y(_12263_));
 sky130_fd_sc_hd__nand2_2 _34303_ (.A(_12242_),
    .B(_12237_),
    .Y(_12264_));
 sky130_fd_sc_hd__nand2_2 _34304_ (.A(_12264_),
    .B(_12261_),
    .Y(_12265_));
 sky130_fd_sc_hd__a21boi_2 _34305_ (.A1(_11979_),
    .A2(_12004_),
    .B1_N(_11984_),
    .Y(_12266_));
 sky130_fd_sc_hd__nand3b_2 _34306_ (.A_N(_12261_),
    .B(_12237_),
    .C(_12242_),
    .Y(_12267_));
 sky130_fd_sc_hd__nand3_2 _34307_ (.A(_12265_),
    .B(_12266_),
    .C(_12267_),
    .Y(_12268_));
 sky130_fd_sc_hd__nand2_2 _34308_ (.A(_08391_),
    .B(_07311_),
    .Y(_12269_));
 sky130_fd_sc_hd__nand2_2 _34309_ (.A(_09614_),
    .B(_06387_),
    .Y(_12270_));
 sky130_fd_sc_hd__nor2_2 _34310_ (.A(_12269_),
    .B(_12270_),
    .Y(_12271_));
 sky130_fd_sc_hd__nand2_2 _34311_ (.A(_08388_),
    .B(_06957_),
    .Y(_12272_));
 sky130_fd_sc_hd__inv_2 _34312_ (.A(_12272_),
    .Y(_12273_));
 sky130_fd_sc_hd__nand2_2 _34313_ (.A(_12269_),
    .B(_12270_),
    .Y(_12274_));
 sky130_fd_sc_hd__nand2_2 _34314_ (.A(_12273_),
    .B(_12274_),
    .Y(_12275_));
 sky130_fd_sc_hd__a21o_2 _34315_ (.A1(_12019_),
    .A2(_12021_),
    .B1(_12018_),
    .X(_12276_));
 sky130_fd_sc_hd__and2_2 _34316_ (.A(_12269_),
    .B(_12270_),
    .X(_12277_));
 sky130_fd_sc_hd__o21ai_2 _34317_ (.A1(_12271_),
    .A2(_12277_),
    .B1(_12272_),
    .Y(_12278_));
 sky130_fd_sc_hd__o211ai_2 _34318_ (.A1(_12271_),
    .A2(_12275_),
    .B1(_12276_),
    .C1(_12278_),
    .Y(_12279_));
 sky130_fd_sc_hd__o21ai_2 _34319_ (.A1(_12271_),
    .A2(_12277_),
    .B1(_12273_),
    .Y(_12280_));
 sky130_fd_sc_hd__or2_2 _34320_ (.A(_12269_),
    .B(_12270_),
    .X(_12281_));
 sky130_fd_sc_hd__nand3_2 _34321_ (.A(_12281_),
    .B(_12272_),
    .C(_12274_),
    .Y(_12282_));
 sky130_fd_sc_hd__a21oi_2 _34322_ (.A1(_12019_),
    .A2(_12021_),
    .B1(_12018_),
    .Y(_12283_));
 sky130_fd_sc_hd__nand3_2 _34323_ (.A(_12280_),
    .B(_12282_),
    .C(_12283_),
    .Y(_12284_));
 sky130_fd_sc_hd__nand2_2 _34324_ (.A(_12279_),
    .B(_12284_),
    .Y(_12285_));
 sky130_fd_sc_hd__nand2_2 _34325_ (.A(_07894_),
    .B(_06946_),
    .Y(_12286_));
 sky130_fd_sc_hd__nand2_2 _34326_ (.A(_07723_),
    .B(_19588_),
    .Y(_12287_));
 sky130_fd_sc_hd__nor2_2 _34327_ (.A(_12286_),
    .B(_12287_),
    .Y(_12288_));
 sky130_fd_sc_hd__nor2_2 _34328_ (.A(_11251_),
    .B(_08604_),
    .Y(_12289_));
 sky130_fd_sc_hd__and2_2 _34329_ (.A(_12286_),
    .B(_12287_),
    .X(_12290_));
 sky130_fd_sc_hd__nor3_2 _34330_ (.A(_12288_),
    .B(_12289_),
    .C(_12290_),
    .Y(_12291_));
 sky130_fd_sc_hd__o21ai_2 _34331_ (.A1(_12288_),
    .A2(_12290_),
    .B1(_12289_),
    .Y(_12292_));
 sky130_fd_sc_hd__and2b_2 _34332_ (.A_N(_12291_),
    .B(_12292_),
    .X(_12293_));
 sky130_fd_sc_hd__nand2_2 _34333_ (.A(_12285_),
    .B(_12293_),
    .Y(_12294_));
 sky130_fd_sc_hd__or2b_2 _34334_ (.A(_12291_),
    .B_N(_12292_),
    .X(_12295_));
 sky130_fd_sc_hd__nand3_2 _34335_ (.A(_12295_),
    .B(_12279_),
    .C(_12284_),
    .Y(_12296_));
 sky130_fd_sc_hd__nand2_2 _34336_ (.A(_11997_),
    .B(_11998_),
    .Y(_12297_));
 sky130_fd_sc_hd__nand2_2 _34337_ (.A(_12297_),
    .B(_12002_),
    .Y(_12298_));
 sky130_fd_sc_hd__a21o_2 _34338_ (.A1(_12294_),
    .A2(_12296_),
    .B1(_12298_),
    .X(_12299_));
 sky130_fd_sc_hd__nand3_2 _34339_ (.A(_12294_),
    .B(_12296_),
    .C(_12298_),
    .Y(_12300_));
 sky130_fd_sc_hd__nand2_2 _34340_ (.A(_12026_),
    .B(_12035_),
    .Y(_12301_));
 sky130_fd_sc_hd__nand2_2 _34341_ (.A(_12301_),
    .B(_12027_),
    .Y(_12302_));
 sky130_fd_sc_hd__a21oi_2 _34342_ (.A1(_12299_),
    .A2(_12300_),
    .B1(_12302_),
    .Y(_12303_));
 sky130_fd_sc_hd__and2_2 _34343_ (.A(_12301_),
    .B(_12027_),
    .X(_12304_));
 sky130_fd_sc_hd__buf_1 _34344_ (.A(_12304_),
    .X(_12305_));
 sky130_fd_sc_hd__nand2_2 _34345_ (.A(_12299_),
    .B(_12300_),
    .Y(_12306_));
 sky130_fd_sc_hd__nor2_2 _34346_ (.A(_12305_),
    .B(_12306_),
    .Y(_12307_));
 sky130_fd_sc_hd__o2bb2ai_2 _34347_ (.A1_N(_12263_),
    .A2_N(_12268_),
    .B1(_12303_),
    .B2(_12307_),
    .Y(_12308_));
 sky130_fd_sc_hd__nand2_2 _34348_ (.A(_12306_),
    .B(_12302_),
    .Y(_12309_));
 sky130_fd_sc_hd__nand3_2 _34349_ (.A(_12299_),
    .B(_12300_),
    .C(_12305_),
    .Y(_12310_));
 sky130_fd_sc_hd__nand2_2 _34350_ (.A(_12309_),
    .B(_12310_),
    .Y(_12311_));
 sky130_fd_sc_hd__nand3_2 _34351_ (.A(_12311_),
    .B(_12268_),
    .C(_12263_),
    .Y(_12312_));
 sky130_fd_sc_hd__nand3_2 _34352_ (.A(_12203_),
    .B(_12308_),
    .C(_12312_),
    .Y(_12313_));
 sky130_fd_sc_hd__and3_2 _34353_ (.A(_12294_),
    .B(_12296_),
    .C(_12298_),
    .X(_12314_));
 sky130_fd_sc_hd__nand2_2 _34354_ (.A(_12299_),
    .B(_12302_),
    .Y(_12315_));
 sky130_fd_sc_hd__a21oi_2 _34355_ (.A1(_12294_),
    .A2(_12296_),
    .B1(_12298_),
    .Y(_12316_));
 sky130_fd_sc_hd__o21ai_2 _34356_ (.A1(_12316_),
    .A2(_12314_),
    .B1(_12305_),
    .Y(_12317_));
 sky130_fd_sc_hd__o21ai_2 _34357_ (.A1(_12314_),
    .A2(_12315_),
    .B1(_12317_),
    .Y(_12318_));
 sky130_fd_sc_hd__nand3_2 _34358_ (.A(_12318_),
    .B(_12268_),
    .C(_12263_),
    .Y(_12319_));
 sky130_fd_sc_hd__inv_2 _34359_ (.A(_12310_),
    .Y(_12320_));
 sky130_fd_sc_hd__and2_2 _34360_ (.A(_12306_),
    .B(_12302_),
    .X(_12321_));
 sky130_fd_sc_hd__o2bb2ai_2 _34361_ (.A1_N(_12263_),
    .A2_N(_12268_),
    .B1(_12320_),
    .B2(_12321_),
    .Y(_12322_));
 sky130_fd_sc_hd__o2111ai_2 _34362_ (.A1(_12202_),
    .A2(_12055_),
    .B1(_12014_),
    .C1(_12319_),
    .D1(_12322_),
    .Y(_12323_));
 sky130_fd_sc_hd__nand2_2 _34363_ (.A(_12111_),
    .B(_12084_),
    .Y(_12324_));
 sky130_fd_sc_hd__and2_2 _34364_ (.A(_12324_),
    .B(_12087_),
    .X(_12325_));
 sky130_fd_sc_hd__a21o_2 _34365_ (.A1(_12031_),
    .A2(_12029_),
    .B1(_12028_),
    .X(_12326_));
 sky130_fd_sc_hd__nand2_2 _34366_ (.A(_09018_),
    .B(_09248_),
    .Y(_12327_));
 sky130_fd_sc_hd__nand2_2 _34367_ (.A(_06828_),
    .B(_07590_),
    .Y(_12328_));
 sky130_fd_sc_hd__nor2_2 _34368_ (.A(_12327_),
    .B(_12328_),
    .Y(_12329_));
 sky130_fd_sc_hd__and2_2 _34369_ (.A(_12327_),
    .B(_12328_),
    .X(_12330_));
 sky130_fd_sc_hd__nand2_2 _34370_ (.A(_09386_),
    .B(_08651_),
    .Y(_12331_));
 sky130_fd_sc_hd__o21ai_2 _34371_ (.A1(_12329_),
    .A2(_12330_),
    .B1(_12331_),
    .Y(_12332_));
 sky130_fd_sc_hd__or2_2 _34372_ (.A(_12327_),
    .B(_12328_),
    .X(_12333_));
 sky130_fd_sc_hd__inv_2 _34373_ (.A(_12331_),
    .Y(_12334_));
 sky130_fd_sc_hd__nand2_2 _34374_ (.A(_12327_),
    .B(_12328_),
    .Y(_12335_));
 sky130_fd_sc_hd__nand3_2 _34375_ (.A(_12333_),
    .B(_12334_),
    .C(_12335_),
    .Y(_12336_));
 sky130_fd_sc_hd__nand3_2 _34376_ (.A(_12326_),
    .B(_12332_),
    .C(_12336_),
    .Y(_12337_));
 sky130_fd_sc_hd__o21ai_2 _34377_ (.A1(_12329_),
    .A2(_12330_),
    .B1(_12334_),
    .Y(_12338_));
 sky130_fd_sc_hd__nand3_2 _34378_ (.A(_12333_),
    .B(_12331_),
    .C(_12335_),
    .Y(_12339_));
 sky130_fd_sc_hd__a21oi_2 _34379_ (.A1(_12031_),
    .A2(_12029_),
    .B1(_12028_),
    .Y(_12340_));
 sky130_fd_sc_hd__nand3_2 _34380_ (.A(_12338_),
    .B(_12339_),
    .C(_12340_),
    .Y(_12341_));
 sky130_fd_sc_hd__a21o_2 _34381_ (.A1(_12072_),
    .A2(_12071_),
    .B1(_12065_),
    .X(_12342_));
 sky130_fd_sc_hd__a21o_2 _34382_ (.A1(_12337_),
    .A2(_12341_),
    .B1(_12342_),
    .X(_12343_));
 sky130_fd_sc_hd__nand2_2 _34383_ (.A(_12078_),
    .B(_12079_),
    .Y(_12344_));
 sky130_fd_sc_hd__nand2_2 _34384_ (.A(_12344_),
    .B(_12074_),
    .Y(_12345_));
 sky130_fd_sc_hd__nand3_2 _34385_ (.A(_12337_),
    .B(_12341_),
    .C(_12342_),
    .Y(_12346_));
 sky130_fd_sc_hd__and3_2 _34386_ (.A(_12343_),
    .B(_12345_),
    .C(_12346_),
    .X(_12347_));
 sky130_fd_sc_hd__nor2_2 _34387_ (.A(_12089_),
    .B(_12091_),
    .Y(_12348_));
 sky130_fd_sc_hd__buf_1 _34388_ (.A(_08497_),
    .X(_12349_));
 sky130_fd_sc_hd__a22o_2 _34389_ (.A1(_19364_),
    .A2(_12349_),
    .B1(_19366_),
    .B2(_19571_),
    .X(_12350_));
 sky130_fd_sc_hd__nand2_2 _34390_ (.A(_19368_),
    .B(_08664_),
    .Y(_12351_));
 sky130_fd_sc_hd__nand3b_2 _34391_ (.A_N(_12348_),
    .B(_12350_),
    .C(_12351_),
    .Y(_12352_));
 sky130_fd_sc_hd__a22oi_2 _34392_ (.A1(_19364_),
    .A2(_12349_),
    .B1(_19366_),
    .B2(_19571_),
    .Y(_12353_));
 sky130_fd_sc_hd__inv_2 _34393_ (.A(_12351_),
    .Y(_12354_));
 sky130_fd_sc_hd__o21ai_2 _34394_ (.A1(_12353_),
    .A2(_12348_),
    .B1(_12354_),
    .Y(_12355_));
 sky130_fd_sc_hd__a21oi_2 _34395_ (.A1(_12096_),
    .A2(_12092_),
    .B1(_12095_),
    .Y(_12356_));
 sky130_fd_sc_hd__a21o_2 _34396_ (.A1(_12352_),
    .A2(_12355_),
    .B1(_12356_),
    .X(_12357_));
 sky130_fd_sc_hd__inv_2 _34397_ (.A(_12357_),
    .Y(_12358_));
 sky130_fd_sc_hd__nand2_2 _34398_ (.A(_06256_),
    .B(_08645_),
    .Y(_12359_));
 sky130_fd_sc_hd__nand2_2 _34399_ (.A(_19373_),
    .B(_19561_),
    .Y(_12360_));
 sky130_fd_sc_hd__nor2_2 _34400_ (.A(_12359_),
    .B(_12360_),
    .Y(_12361_));
 sky130_fd_sc_hd__nand2_2 _34401_ (.A(_12359_),
    .B(_12360_),
    .Y(_12362_));
 sky130_fd_sc_hd__inv_2 _34402_ (.A(_12362_),
    .Y(_12363_));
 sky130_fd_sc_hd__nand2_2 _34403_ (.A(_06616_),
    .B(_09736_),
    .Y(_12364_));
 sky130_fd_sc_hd__inv_2 _34404_ (.A(_12364_),
    .Y(_12365_));
 sky130_fd_sc_hd__o21ai_2 _34405_ (.A1(_12361_),
    .A2(_12363_),
    .B1(_12365_),
    .Y(_12366_));
 sky130_fd_sc_hd__nand3b_2 _34406_ (.A_N(_12361_),
    .B(_12364_),
    .C(_12362_),
    .Y(_12367_));
 sky130_fd_sc_hd__nand2_2 _34407_ (.A(_12366_),
    .B(_12367_),
    .Y(_12368_));
 sky130_fd_sc_hd__nand3_2 _34408_ (.A(_12352_),
    .B(_12356_),
    .C(_12355_),
    .Y(_12369_));
 sky130_fd_sc_hd__nand2_2 _34409_ (.A(_12368_),
    .B(_12369_),
    .Y(_12370_));
 sky130_fd_sc_hd__a21o_2 _34410_ (.A1(_12357_),
    .A2(_12369_),
    .B1(_12368_),
    .X(_12371_));
 sky130_fd_sc_hd__o21a_2 _34411_ (.A1(_12358_),
    .A2(_12370_),
    .B1(_12371_),
    .X(_12372_));
 sky130_fd_sc_hd__a21o_2 _34412_ (.A1(_12343_),
    .A2(_12346_),
    .B1(_12345_),
    .X(_12373_));
 sky130_fd_sc_hd__nand2_2 _34413_ (.A(_12372_),
    .B(_12373_),
    .Y(_12374_));
 sky130_fd_sc_hd__a21oi_2 _34414_ (.A1(_12343_),
    .A2(_12346_),
    .B1(_12345_),
    .Y(_12375_));
 sky130_fd_sc_hd__o21ai_2 _34415_ (.A1(_12370_),
    .A2(_12358_),
    .B1(_12371_),
    .Y(_12376_));
 sky130_fd_sc_hd__o21ai_2 _34416_ (.A1(_12375_),
    .A2(_12347_),
    .B1(_12376_),
    .Y(_12377_));
 sky130_fd_sc_hd__nand2_2 _34417_ (.A(_12040_),
    .B(_12046_),
    .Y(_12378_));
 sky130_fd_sc_hd__nand2_2 _34418_ (.A(_12378_),
    .B(_12044_),
    .Y(_12379_));
 sky130_fd_sc_hd__o211ai_2 _34419_ (.A1(_12347_),
    .A2(_12374_),
    .B1(_12377_),
    .C1(_12379_),
    .Y(_12380_));
 sky130_fd_sc_hd__o21ai_2 _34420_ (.A1(_12375_),
    .A2(_12347_),
    .B1(_12372_),
    .Y(_12381_));
 sky130_fd_sc_hd__a21boi_2 _34421_ (.A1(_12040_),
    .A2(_12046_),
    .B1_N(_12044_),
    .Y(_12382_));
 sky130_fd_sc_hd__nand3_2 _34422_ (.A(_12343_),
    .B(_12345_),
    .C(_12346_),
    .Y(_12383_));
 sky130_fd_sc_hd__nand3_2 _34423_ (.A(_12373_),
    .B(_12383_),
    .C(_12376_),
    .Y(_12384_));
 sky130_fd_sc_hd__nand3_2 _34424_ (.A(_12381_),
    .B(_12382_),
    .C(_12384_),
    .Y(_12385_));
 sky130_fd_sc_hd__nand2_2 _34425_ (.A(_12380_),
    .B(_12385_),
    .Y(_12386_));
 sky130_fd_sc_hd__nor2_2 _34426_ (.A(_12325_),
    .B(_12386_),
    .Y(_12387_));
 sky130_fd_sc_hd__nand2_2 _34427_ (.A(_12324_),
    .B(_12087_),
    .Y(_12388_));
 sky130_fd_sc_hd__a21oi_2 _34428_ (.A1(_12380_),
    .A2(_12385_),
    .B1(_12388_),
    .Y(_12389_));
 sky130_fd_sc_hd__o2bb2ai_2 _34429_ (.A1_N(_12313_),
    .A2_N(_12323_),
    .B1(_12387_),
    .B2(_12389_),
    .Y(_12390_));
 sky130_fd_sc_hd__a31oi_2 _34430_ (.A1(_12382_),
    .A2(_12381_),
    .A3(_12384_),
    .B1(_12325_),
    .Y(_12391_));
 sky130_fd_sc_hd__a21oi_2 _34431_ (.A1(_12380_),
    .A2(_12391_),
    .B1(_12389_),
    .Y(_12392_));
 sky130_fd_sc_hd__nand3_2 _34432_ (.A(_12392_),
    .B(_12313_),
    .C(_12323_),
    .Y(_12393_));
 sky130_fd_sc_hd__nand3_2 _34433_ (.A(_12199_),
    .B(_12390_),
    .C(_12393_),
    .Y(_12394_));
 sky130_fd_sc_hd__nand2_2 _34434_ (.A(_12386_),
    .B(_12325_),
    .Y(_12395_));
 sky130_fd_sc_hd__nand2_2 _34435_ (.A(_12391_),
    .B(_12380_),
    .Y(_12396_));
 sky130_fd_sc_hd__nand2_2 _34436_ (.A(_12395_),
    .B(_12396_),
    .Y(_12397_));
 sky130_fd_sc_hd__a21o_2 _34437_ (.A1(_12323_),
    .A2(_12313_),
    .B1(_12397_),
    .X(_12398_));
 sky130_fd_sc_hd__a21boi_2 _34438_ (.A1(_12137_),
    .A2(_12057_),
    .B1_N(_12062_),
    .Y(_12399_));
 sky130_fd_sc_hd__nand3_2 _34439_ (.A(_12397_),
    .B(_12323_),
    .C(_12313_),
    .Y(_12400_));
 sky130_fd_sc_hd__nand3_2 _34440_ (.A(_12398_),
    .B(_12399_),
    .C(_12400_),
    .Y(_12401_));
 sky130_fd_sc_hd__o22a_2 _34441_ (.A1(_06807_),
    .A2(_12104_),
    .B1(_12102_),
    .B2(_12101_),
    .X(_12402_));
 sky130_fd_sc_hd__nand2_2 _34442_ (.A(_05857_),
    .B(_11410_),
    .Y(_12403_));
 sky130_fd_sc_hd__nand2_2 _34443_ (.A(_09247_),
    .B(_19548_),
    .Y(_12404_));
 sky130_fd_sc_hd__nor2_2 _34444_ (.A(_12403_),
    .B(_12404_),
    .Y(_12405_));
 sky130_fd_sc_hd__and2_2 _34445_ (.A(_12403_),
    .B(_12404_),
    .X(_12406_));
 sky130_fd_sc_hd__nand2_2 _34446_ (.A(_08953_),
    .B(_11037_),
    .Y(_12407_));
 sky130_fd_sc_hd__o21ai_2 _34447_ (.A1(_12405_),
    .A2(_12406_),
    .B1(_12407_),
    .Y(_12408_));
 sky130_fd_sc_hd__nand2_2 _34448_ (.A(_12403_),
    .B(_12404_),
    .Y(_12409_));
 sky130_fd_sc_hd__inv_2 _34449_ (.A(_12407_),
    .Y(_12410_));
 sky130_fd_sc_hd__nand3b_2 _34450_ (.A_N(_12405_),
    .B(_12409_),
    .C(_12410_),
    .Y(_12411_));
 sky130_fd_sc_hd__nand3b_2 _34451_ (.A_N(_12402_),
    .B(_12408_),
    .C(_12411_),
    .Y(_12412_));
 sky130_fd_sc_hd__o21ai_2 _34452_ (.A1(_12405_),
    .A2(_12406_),
    .B1(_12410_),
    .Y(_12413_));
 sky130_fd_sc_hd__nand3b_2 _34453_ (.A_N(_12405_),
    .B(_12409_),
    .C(_12407_),
    .Y(_12414_));
 sky130_fd_sc_hd__nand3_2 _34454_ (.A(_12413_),
    .B(_12414_),
    .C(_12402_),
    .Y(_12415_));
 sky130_fd_sc_hd__a21oi_2 _34455_ (.A1(_11869_),
    .A2(_11867_),
    .B1(_11866_),
    .Y(_12416_));
 sky130_fd_sc_hd__inv_2 _34456_ (.A(_12416_),
    .Y(_12417_));
 sky130_fd_sc_hd__a21oi_2 _34457_ (.A1(_12412_),
    .A2(_12415_),
    .B1(_12417_),
    .Y(_12418_));
 sky130_fd_sc_hd__nand3_2 _34458_ (.A(_12412_),
    .B(_12415_),
    .C(_12417_),
    .Y(_12419_));
 sky130_fd_sc_hd__inv_2 _34459_ (.A(_12419_),
    .Y(_12420_));
 sky130_fd_sc_hd__a21oi_2 _34460_ (.A1(_12094_),
    .A2(_12097_),
    .B1(_12098_),
    .Y(_12421_));
 sky130_fd_sc_hd__o21ai_2 _34461_ (.A1(_12108_),
    .A2(_12421_),
    .B1(_12100_),
    .Y(_12422_));
 sky130_fd_sc_hd__o21bai_2 _34462_ (.A1(_12418_),
    .A2(_12420_),
    .B1_N(_12422_),
    .Y(_12423_));
 sky130_fd_sc_hd__a21o_2 _34463_ (.A1(_12412_),
    .A2(_12415_),
    .B1(_12417_),
    .X(_12424_));
 sky130_fd_sc_hd__nand3_2 _34464_ (.A(_12424_),
    .B(_12422_),
    .C(_12419_),
    .Y(_12425_));
 sky130_fd_sc_hd__nand2_2 _34465_ (.A(_11880_),
    .B(_11873_),
    .Y(_12426_));
 sky130_fd_sc_hd__a21o_2 _34466_ (.A1(_12423_),
    .A2(_12425_),
    .B1(_12426_),
    .X(_12427_));
 sky130_fd_sc_hd__o21ai_2 _34467_ (.A1(_11889_),
    .A2(_11882_),
    .B1(_11890_),
    .Y(_12428_));
 sky130_fd_sc_hd__nand3_2 _34468_ (.A(_12423_),
    .B(_12425_),
    .C(_12426_),
    .Y(_12429_));
 sky130_fd_sc_hd__nand3_2 _34469_ (.A(_12427_),
    .B(_12428_),
    .C(_12429_),
    .Y(_12430_));
 sky130_fd_sc_hd__a21oi_2 _34470_ (.A1(_12423_),
    .A2(_12425_),
    .B1(_12426_),
    .Y(_12431_));
 sky130_fd_sc_hd__inv_2 _34471_ (.A(_12426_),
    .Y(_12432_));
 sky130_fd_sc_hd__a21oi_2 _34472_ (.A1(_12424_),
    .A2(_12419_),
    .B1(_12422_),
    .Y(_12433_));
 sky130_fd_sc_hd__nor3b_2 _34473_ (.A(_12432_),
    .B(_12433_),
    .C_N(_12425_),
    .Y(_12434_));
 sky130_fd_sc_hd__o21bai_2 _34474_ (.A1(_12431_),
    .A2(_12434_),
    .B1_N(_12428_),
    .Y(_12435_));
 sky130_fd_sc_hd__nand2_2 _34475_ (.A(_06199_),
    .B(_19540_),
    .Y(_12436_));
 sky130_fd_sc_hd__nand2_2 _34476_ (.A(_18156_),
    .B(_19391_),
    .Y(_12437_));
 sky130_fd_sc_hd__o21ai_2 _34477_ (.A1(_12436_),
    .A2(_12437_),
    .B1(_11029_),
    .Y(_12438_));
 sky130_fd_sc_hd__a21o_2 _34478_ (.A1(_12436_),
    .A2(_12437_),
    .B1(_12438_),
    .X(_12439_));
 sky130_fd_sc_hd__nor2_2 _34479_ (.A(_12436_),
    .B(_12437_),
    .Y(_12440_));
 sky130_fd_sc_hd__and2_2 _34480_ (.A(_12436_),
    .B(_12437_),
    .X(_12441_));
 sky130_fd_sc_hd__o21ai_2 _34481_ (.A1(_12440_),
    .A2(_12441_),
    .B1(_11025_),
    .Y(_12442_));
 sky130_fd_sc_hd__a21oi_2 _34482_ (.A1(_11025_),
    .A2(_11904_),
    .B1(_11903_),
    .Y(_12443_));
 sky130_fd_sc_hd__a21oi_2 _34483_ (.A1(_12439_),
    .A2(_12442_),
    .B1(_12443_),
    .Y(_12444_));
 sky130_fd_sc_hd__nand3_2 _34484_ (.A(_12439_),
    .B(_12442_),
    .C(_12443_),
    .Y(_12445_));
 sky130_fd_sc_hd__nand2_2 _34485_ (.A(_11918_),
    .B(_12445_),
    .Y(_12446_));
 sky130_fd_sc_hd__nor2_2 _34486_ (.A(_12444_),
    .B(_12446_),
    .Y(_12447_));
 sky130_fd_sc_hd__a21o_2 _34487_ (.A1(_12439_),
    .A2(_12442_),
    .B1(_12443_),
    .X(_12448_));
 sky130_fd_sc_hd__a21oi_2 _34488_ (.A1(_12448_),
    .A2(_12445_),
    .B1(_11919_),
    .Y(_12449_));
 sky130_fd_sc_hd__nand2_2 _34489_ (.A(_11912_),
    .B(_11919_),
    .Y(_12450_));
 sky130_fd_sc_hd__nand2_2 _34490_ (.A(_12450_),
    .B(_11909_),
    .Y(_12451_));
 sky130_fd_sc_hd__o21bai_2 _34491_ (.A1(_12447_),
    .A2(_12449_),
    .B1_N(_12451_),
    .Y(_12452_));
 sky130_fd_sc_hd__a21o_2 _34492_ (.A1(_12448_),
    .A2(_12445_),
    .B1(_11919_),
    .X(_12453_));
 sky130_fd_sc_hd__nand3b_2 _34493_ (.A_N(_12447_),
    .B(_12453_),
    .C(_12451_),
    .Y(_12454_));
 sky130_fd_sc_hd__nor2_2 _34494_ (.A(_11761_),
    .B(_11916_),
    .Y(_12455_));
 sky130_fd_sc_hd__buf_1 _34495_ (.A(_12455_),
    .X(_12456_));
 sky130_fd_sc_hd__inv_2 _34496_ (.A(_12456_),
    .Y(_12457_));
 sky130_fd_sc_hd__and3_2 _34497_ (.A(_12452_),
    .B(_12454_),
    .C(_12457_),
    .X(_12458_));
 sky130_fd_sc_hd__a21oi_2 _34498_ (.A1(_12452_),
    .A2(_12454_),
    .B1(_12457_),
    .Y(_12459_));
 sky130_fd_sc_hd__o2bb2ai_2 _34499_ (.A1_N(_12430_),
    .A2_N(_12435_),
    .B1(_12458_),
    .B2(_12459_),
    .Y(_12460_));
 sky130_fd_sc_hd__nor2_2 _34500_ (.A(_12459_),
    .B(_12458_),
    .Y(_12461_));
 sky130_fd_sc_hd__nand3_2 _34501_ (.A(_12461_),
    .B(_12435_),
    .C(_12430_),
    .Y(_12462_));
 sky130_fd_sc_hd__nand2_2 _34502_ (.A(_12117_),
    .B(_12123_),
    .Y(_12463_));
 sky130_fd_sc_hd__nand2_2 _34503_ (.A(_12463_),
    .B(_12121_),
    .Y(_12464_));
 sky130_fd_sc_hd__a21o_2 _34504_ (.A1(_12460_),
    .A2(_12462_),
    .B1(_12464_),
    .X(_12465_));
 sky130_fd_sc_hd__nand3_2 _34505_ (.A(_12460_),
    .B(_12464_),
    .C(_12462_),
    .Y(_12466_));
 sky130_fd_sc_hd__a21bo_2 _34506_ (.A1(_11936_),
    .A2(_11892_),
    .B1_N(_11897_),
    .X(_12467_));
 sky130_fd_sc_hd__a21oi_2 _34507_ (.A1(_12465_),
    .A2(_12466_),
    .B1(_12467_),
    .Y(_12468_));
 sky130_fd_sc_hd__and3_2 _34508_ (.A(_12465_),
    .B(_12466_),
    .C(_12467_),
    .X(_12469_));
 sky130_fd_sc_hd__o2bb2ai_2 _34509_ (.A1_N(_12394_),
    .A2_N(_12401_),
    .B1(_12468_),
    .B2(_12469_),
    .Y(_12470_));
 sky130_fd_sc_hd__and3_2 _34510_ (.A(_12460_),
    .B(_12464_),
    .C(_12462_),
    .X(_12471_));
 sky130_fd_sc_hd__nand2_2 _34511_ (.A(_12465_),
    .B(_12467_),
    .Y(_12472_));
 sky130_fd_sc_hd__a21oi_2 _34512_ (.A1(_12460_),
    .A2(_12462_),
    .B1(_12464_),
    .Y(_12473_));
 sky130_fd_sc_hd__o21bai_2 _34513_ (.A1(_12473_),
    .A2(_12471_),
    .B1_N(_12467_),
    .Y(_12474_));
 sky130_fd_sc_hd__o2111ai_2 _34514_ (.A1(_12471_),
    .A2(_12472_),
    .B1(_12474_),
    .C1(_12394_),
    .D1(_12401_),
    .Y(_12475_));
 sky130_fd_sc_hd__inv_2 _34515_ (.A(_12138_),
    .Y(_12476_));
 sky130_fd_sc_hd__nand2_2 _34516_ (.A(_12131_),
    .B(_12134_),
    .Y(_12477_));
 sky130_fd_sc_hd__a21oi_2 _34517_ (.A1(_12134_),
    .A2(_12138_),
    .B1(_12131_),
    .Y(_12478_));
 sky130_fd_sc_hd__o22ai_2 _34518_ (.A1(_12476_),
    .A2(_12477_),
    .B1(_12147_),
    .B2(_12478_),
    .Y(_12479_));
 sky130_fd_sc_hd__a21oi_2 _34519_ (.A1(_12470_),
    .A2(_12475_),
    .B1(_12479_),
    .Y(_12480_));
 sky130_fd_sc_hd__a21oi_2 _34520_ (.A1(_12398_),
    .A2(_12400_),
    .B1(_12399_),
    .Y(_12481_));
 sky130_fd_sc_hd__nand3_2 _34521_ (.A(_12465_),
    .B(_12466_),
    .C(_12467_),
    .Y(_12482_));
 sky130_fd_sc_hd__nand3_2 _34522_ (.A(_12401_),
    .B(_12474_),
    .C(_12482_),
    .Y(_12483_));
 sky130_fd_sc_hd__o211a_2 _34523_ (.A1(_12481_),
    .A2(_12483_),
    .B1(_12479_),
    .C1(_12470_),
    .X(_12484_));
 sky130_fd_sc_hd__o22ai_2 _34524_ (.A1(_12194_),
    .A2(_12195_),
    .B1(_12480_),
    .B2(_12484_),
    .Y(_12485_));
 sky130_fd_sc_hd__a22oi_2 _34525_ (.A1(_12474_),
    .A2(_12482_),
    .B1(_12401_),
    .B2(_12394_),
    .Y(_12486_));
 sky130_fd_sc_hd__o2111a_2 _34526_ (.A1(_12471_),
    .A2(_12472_),
    .B1(_12474_),
    .C1(_12394_),
    .D1(_12401_),
    .X(_12487_));
 sky130_fd_sc_hd__o21bai_2 _34527_ (.A1(_12486_),
    .A2(_12487_),
    .B1_N(_12479_),
    .Y(_12488_));
 sky130_fd_sc_hd__nand3_2 _34528_ (.A(_12470_),
    .B(_12479_),
    .C(_12475_),
    .Y(_12489_));
 sky130_fd_sc_hd__nor2_2 _34529_ (.A(_12195_),
    .B(_12194_),
    .Y(_12490_));
 sky130_fd_sc_hd__nand3_2 _34530_ (.A(_12488_),
    .B(_12489_),
    .C(_12490_),
    .Y(_12491_));
 sky130_fd_sc_hd__nand2_2 _34531_ (.A(_12130_),
    .B(_12139_),
    .Y(_12492_));
 sky130_fd_sc_hd__and2_2 _34532_ (.A(_12492_),
    .B(_12147_),
    .X(_12493_));
 sky130_fd_sc_hd__nand2_2 _34533_ (.A(_11861_),
    .B(_12140_),
    .Y(_12494_));
 sky130_fd_sc_hd__a21oi_2 _34534_ (.A1(_12141_),
    .A2(_12140_),
    .B1(_11861_),
    .Y(_12495_));
 sky130_fd_sc_hd__o22ai_2 _34535_ (.A1(_12493_),
    .A2(_12494_),
    .B1(_12161_),
    .B2(_12495_),
    .Y(_12496_));
 sky130_fd_sc_hd__nand3_2 _34536_ (.A(_12485_),
    .B(_12491_),
    .C(_12496_),
    .Y(_12497_));
 sky130_fd_sc_hd__nor2_2 _34537_ (.A(_12190_),
    .B(_12193_),
    .Y(_12498_));
 sky130_fd_sc_hd__nor2_2 _34538_ (.A(_12191_),
    .B(_12192_),
    .Y(_12499_));
 sky130_fd_sc_hd__o22ai_2 _34539_ (.A1(_12498_),
    .A2(_12499_),
    .B1(_12480_),
    .B2(_12484_),
    .Y(_12500_));
 sky130_fd_sc_hd__a21boi_2 _34540_ (.A1(_12150_),
    .A2(_12170_),
    .B1_N(_12142_),
    .Y(_12501_));
 sky130_fd_sc_hd__nor2_2 _34541_ (.A(_12499_),
    .B(_12498_),
    .Y(_12502_));
 sky130_fd_sc_hd__nand3_2 _34542_ (.A(_12488_),
    .B(_12489_),
    .C(_12502_),
    .Y(_12503_));
 sky130_fd_sc_hd__nand3_2 _34543_ (.A(_12500_),
    .B(_12501_),
    .C(_12503_),
    .Y(_12504_));
 sky130_fd_sc_hd__o2bb2ai_2 _34544_ (.A1_N(_12497_),
    .A2_N(_12504_),
    .B1(_12157_),
    .B2(_12155_),
    .Y(_12505_));
 sky130_fd_sc_hd__nand3_2 _34545_ (.A(_12504_),
    .B(_12497_),
    .C(_12164_),
    .Y(_12506_));
 sky130_fd_sc_hd__inv_2 _34546_ (.A(_12171_),
    .Y(_12507_));
 sky130_fd_sc_hd__nand2_2 _34547_ (.A(_12166_),
    .B(_12169_),
    .Y(_12508_));
 sky130_fd_sc_hd__o2bb2ai_2 _34548_ (.A1_N(_11829_),
    .A2_N(_12163_),
    .B1(_12507_),
    .B2(_12508_),
    .Y(_12509_));
 sky130_fd_sc_hd__a21oi_2 _34549_ (.A1(_12505_),
    .A2(_12506_),
    .B1(_12509_),
    .Y(_12510_));
 sky130_fd_sc_hd__nand3_2 _34550_ (.A(_12505_),
    .B(_12509_),
    .C(_12506_),
    .Y(_12511_));
 sky130_fd_sc_hd__inv_2 _34551_ (.A(_12511_),
    .Y(_12512_));
 sky130_fd_sc_hd__nor2_2 _34552_ (.A(_12510_),
    .B(_12512_),
    .Y(_12513_));
 sky130_fd_sc_hd__inv_2 _34553_ (.A(_12513_),
    .Y(_12514_));
 sky130_fd_sc_hd__o22ai_2 _34554_ (.A1(_12185_),
    .A2(_12186_),
    .B1(_12180_),
    .B2(_12182_),
    .Y(_12515_));
 sky130_fd_sc_hd__a31oi_2 _34555_ (.A1(_11853_),
    .A2(_11854_),
    .A3(_12181_),
    .B1(_12515_),
    .Y(_12516_));
 sky130_fd_sc_hd__and3_2 _34556_ (.A(_12189_),
    .B(_12514_),
    .C(_12516_),
    .X(_12517_));
 sky130_fd_sc_hd__and2_2 _34557_ (.A(_12189_),
    .B(_12516_),
    .X(_12518_));
 sky130_fd_sc_hd__nor2_2 _34558_ (.A(_12514_),
    .B(_12518_),
    .Y(_12519_));
 sky130_fd_sc_hd__nor2_2 _34559_ (.A(_12517_),
    .B(_12519_),
    .Y(_02655_));
 sky130_fd_sc_hd__inv_2 _34560_ (.A(_12491_),
    .Y(_12520_));
 sky130_fd_sc_hd__nand2_2 _34561_ (.A(_12485_),
    .B(_12496_),
    .Y(_12521_));
 sky130_fd_sc_hd__o2bb2ai_2 _34562_ (.A1_N(_12164_),
    .A2_N(_12504_),
    .B1(_12520_),
    .B2(_12521_),
    .Y(_12522_));
 sky130_fd_sc_hd__a31oi_2 _34563_ (.A1(_12401_),
    .A2(_12474_),
    .A3(_12482_),
    .B1(_12481_),
    .Y(_12523_));
 sky130_fd_sc_hd__nand3_2 _34564_ (.A(_11514_),
    .B(_10822_),
    .C(_06609_),
    .Y(_12524_));
 sky130_fd_sc_hd__a22o_2 _34565_ (.A1(_10822_),
    .A2(_06609_),
    .B1(_05855_),
    .B2(_11514_),
    .X(_12525_));
 sky130_fd_sc_hd__o21ai_2 _34566_ (.A1(_19626_),
    .A2(_12524_),
    .B1(_12525_),
    .Y(_12526_));
 sky130_fd_sc_hd__nand2_2 _34567_ (.A(\pcpi_mul.rs2[30] ),
    .B(_05502_),
    .Y(_12527_));
 sky130_fd_sc_hd__inv_2 _34568_ (.A(_12527_),
    .Y(_12528_));
 sky130_fd_sc_hd__nand2_2 _34569_ (.A(_12526_),
    .B(_12528_),
    .Y(_12529_));
 sky130_fd_sc_hd__nor2_2 _34570_ (.A(_06502_),
    .B(_12524_),
    .Y(_12530_));
 sky130_fd_sc_hd__nand3b_2 _34571_ (.A_N(_12530_),
    .B(_12525_),
    .C(_12527_),
    .Y(_12531_));
 sky130_fd_sc_hd__o21ai_2 _34572_ (.A1(_06501_),
    .A2(_12209_),
    .B1(_12212_),
    .Y(_12532_));
 sky130_fd_sc_hd__nand2_2 _34573_ (.A(_12216_),
    .B(_12532_),
    .Y(_12533_));
 sky130_fd_sc_hd__nand3_2 _34574_ (.A(_12529_),
    .B(_12531_),
    .C(_12533_),
    .Y(_12534_));
 sky130_fd_sc_hd__nand2_2 _34575_ (.A(_12526_),
    .B(_12527_),
    .Y(_12535_));
 sky130_fd_sc_hd__nand3b_2 _34576_ (.A_N(_12530_),
    .B(_12525_),
    .C(_12528_),
    .Y(_12536_));
 sky130_fd_sc_hd__and2_2 _34577_ (.A(_12216_),
    .B(_12532_),
    .X(_12537_));
 sky130_fd_sc_hd__nand3_2 _34578_ (.A(_12535_),
    .B(_12536_),
    .C(_12537_),
    .Y(_12538_));
 sky130_fd_sc_hd__nor2_2 _34579_ (.A(_09356_),
    .B(_06694_),
    .Y(_12539_));
 sky130_fd_sc_hd__a22oi_2 _34580_ (.A1(_09842_),
    .A2(_06052_),
    .B1(_09838_),
    .B2(_05737_),
    .Y(_12540_));
 sky130_fd_sc_hd__nor2_2 _34581_ (.A(_05617_),
    .B(_10704_),
    .Y(_12541_));
 sky130_fd_sc_hd__nor2_2 _34582_ (.A(_12540_),
    .B(_12541_),
    .Y(_12542_));
 sky130_fd_sc_hd__nor2_2 _34583_ (.A(_12539_),
    .B(_12542_),
    .Y(_12543_));
 sky130_fd_sc_hd__a22o_2 _34584_ (.A1(_09842_),
    .A2(_19616_),
    .B1(_10141_),
    .B2(_07210_),
    .X(_12544_));
 sky130_fd_sc_hd__nand2_2 _34585_ (.A(_12539_),
    .B(_12544_),
    .Y(_12545_));
 sky130_fd_sc_hd__nor2_2 _34586_ (.A(_12541_),
    .B(_12545_),
    .Y(_12546_));
 sky130_fd_sc_hd__o2bb2ai_2 _34587_ (.A1_N(_12534_),
    .A2_N(_12538_),
    .B1(_12543_),
    .B2(_12546_),
    .Y(_12547_));
 sky130_fd_sc_hd__nand2_2 _34588_ (.A(_12218_),
    .B(_12235_),
    .Y(_12548_));
 sky130_fd_sc_hd__nand2_2 _34589_ (.A(_12548_),
    .B(_12222_),
    .Y(_12549_));
 sky130_fd_sc_hd__nor2_2 _34590_ (.A(_12546_),
    .B(_12543_),
    .Y(_12550_));
 sky130_fd_sc_hd__nand3_2 _34591_ (.A(_12538_),
    .B(_12534_),
    .C(_12550_),
    .Y(_12551_));
 sky130_fd_sc_hd__nand3_2 _34592_ (.A(_12547_),
    .B(_12549_),
    .C(_12551_),
    .Y(_12552_));
 sky130_fd_sc_hd__inv_2 _34593_ (.A(_12539_),
    .Y(_12553_));
 sky130_fd_sc_hd__nor2_2 _34594_ (.A(_12553_),
    .B(_12542_),
    .Y(_12554_));
 sky130_fd_sc_hd__and2_2 _34595_ (.A(_12542_),
    .B(_12553_),
    .X(_12555_));
 sky130_fd_sc_hd__o2bb2ai_2 _34596_ (.A1_N(_12534_),
    .A2_N(_12538_),
    .B1(_12554_),
    .B2(_12555_),
    .Y(_12556_));
 sky130_fd_sc_hd__a21boi_2 _34597_ (.A1(_12218_),
    .A2(_12235_),
    .B1_N(_12222_),
    .Y(_12557_));
 sky130_fd_sc_hd__o211ai_2 _34598_ (.A1(_12543_),
    .A2(_12546_),
    .B1(_12534_),
    .C1(_12538_),
    .Y(_12558_));
 sky130_fd_sc_hd__nand3_2 _34599_ (.A(_12556_),
    .B(_12557_),
    .C(_12558_),
    .Y(_12559_));
 sky130_fd_sc_hd__nand2_2 _34600_ (.A(_12552_),
    .B(_12559_),
    .Y(_12560_));
 sky130_fd_sc_hd__nand2_2 _34601_ (.A(_19327_),
    .B(_05910_),
    .Y(_12561_));
 sky130_fd_sc_hd__nand2_2 _34602_ (.A(_09120_),
    .B(_06732_),
    .Y(_12562_));
 sky130_fd_sc_hd__nor2_2 _34603_ (.A(_12561_),
    .B(_12562_),
    .Y(_12563_));
 sky130_fd_sc_hd__and2_2 _34604_ (.A(_12561_),
    .B(_12562_),
    .X(_12564_));
 sky130_fd_sc_hd__nand2_2 _34605_ (.A(_10862_),
    .B(_19600_),
    .Y(_12565_));
 sky130_fd_sc_hd__o21ai_2 _34606_ (.A1(_12563_),
    .A2(_12564_),
    .B1(_12565_),
    .Y(_12566_));
 sky130_fd_sc_hd__nand2_2 _34607_ (.A(_12561_),
    .B(_12562_),
    .Y(_12567_));
 sky130_fd_sc_hd__inv_2 _34608_ (.A(_12565_),
    .Y(_12568_));
 sky130_fd_sc_hd__nand3b_2 _34609_ (.A_N(_12563_),
    .B(_12567_),
    .C(_12568_),
    .Y(_12569_));
 sky130_fd_sc_hd__o21ai_2 _34610_ (.A1(_12223_),
    .A2(_12224_),
    .B1(_12232_),
    .Y(_12570_));
 sky130_fd_sc_hd__nand3_2 _34611_ (.A(_12566_),
    .B(_12569_),
    .C(_12570_),
    .Y(_12571_));
 sky130_fd_sc_hd__o21ai_2 _34612_ (.A1(_12563_),
    .A2(_12564_),
    .B1(_12568_),
    .Y(_12572_));
 sky130_fd_sc_hd__nand3b_2 _34613_ (.A_N(_12563_),
    .B(_12567_),
    .C(_12565_),
    .Y(_12573_));
 sky130_fd_sc_hd__a21oi_2 _34614_ (.A1(_12230_),
    .A2(_12231_),
    .B1(_12225_),
    .Y(_12574_));
 sky130_fd_sc_hd__nand3_2 _34615_ (.A(_12572_),
    .B(_12573_),
    .C(_12574_),
    .Y(_12575_));
 sky130_fd_sc_hd__a21oi_2 _34616_ (.A1(_12249_),
    .A2(_12247_),
    .B1(_12246_),
    .Y(_12576_));
 sky130_fd_sc_hd__inv_2 _34617_ (.A(_12576_),
    .Y(_12577_));
 sky130_fd_sc_hd__a21oi_2 _34618_ (.A1(_12571_),
    .A2(_12575_),
    .B1(_12577_),
    .Y(_12578_));
 sky130_fd_sc_hd__nand2_2 _34619_ (.A(_12571_),
    .B(_12575_),
    .Y(_12579_));
 sky130_fd_sc_hd__nor2_2 _34620_ (.A(_12576_),
    .B(_12579_),
    .Y(_12580_));
 sky130_fd_sc_hd__nor2_2 _34621_ (.A(_12578_),
    .B(_12580_),
    .Y(_12581_));
 sky130_fd_sc_hd__nand2_2 _34622_ (.A(_12560_),
    .B(_12581_),
    .Y(_12582_));
 sky130_fd_sc_hd__inv_2 _34623_ (.A(_12571_),
    .Y(_12583_));
 sky130_fd_sc_hd__nand2_2 _34624_ (.A(_12575_),
    .B(_12577_),
    .Y(_12584_));
 sky130_fd_sc_hd__nand2_2 _34625_ (.A(_12579_),
    .B(_12576_),
    .Y(_12585_));
 sky130_fd_sc_hd__o21ai_2 _34626_ (.A1(_12583_),
    .A2(_12584_),
    .B1(_12585_),
    .Y(_12586_));
 sky130_fd_sc_hd__nand3_2 _34627_ (.A(_12552_),
    .B(_12559_),
    .C(_12586_),
    .Y(_12587_));
 sky130_fd_sc_hd__a21boi_2 _34628_ (.A1(_12242_),
    .A2(_12261_),
    .B1_N(_12237_),
    .Y(_12588_));
 sky130_fd_sc_hd__a21oi_2 _34629_ (.A1(_12582_),
    .A2(_12587_),
    .B1(_12588_),
    .Y(_12589_));
 sky130_fd_sc_hd__inv_2 _34630_ (.A(_12253_),
    .Y(_12590_));
 sky130_fd_sc_hd__and2_2 _34631_ (.A(_12256_),
    .B(_12257_),
    .X(_12591_));
 sky130_fd_sc_hd__and4_2 _34632_ (.A(_07483_),
    .B(_07906_),
    .C(_08089_),
    .D(_06944_),
    .X(_12592_));
 sky130_fd_sc_hd__nor2_2 _34633_ (.A(_07052_),
    .B(_08946_),
    .Y(_12593_));
 sky130_fd_sc_hd__a22o_2 _34634_ (.A1(_07483_),
    .A2(_06944_),
    .B1(_07478_),
    .B2(_08089_),
    .X(_12594_));
 sky130_fd_sc_hd__nand2_2 _34635_ (.A(_12593_),
    .B(_12594_),
    .Y(_12595_));
 sky130_fd_sc_hd__inv_2 _34636_ (.A(_07480_),
    .Y(_12596_));
 sky130_fd_sc_hd__inv_2 _34637_ (.A(_07906_),
    .Y(_12597_));
 sky130_fd_sc_hd__o22a_2 _34638_ (.A1(_12596_),
    .A2(_07832_),
    .B1(_12597_),
    .B2(_08604_),
    .X(_12598_));
 sky130_fd_sc_hd__inv_2 _34639_ (.A(_12593_),
    .Y(_12599_));
 sky130_fd_sc_hd__o21ai_2 _34640_ (.A1(_12592_),
    .A2(_12598_),
    .B1(_12599_),
    .Y(_12600_));
 sky130_fd_sc_hd__o21ai_2 _34641_ (.A1(_12592_),
    .A2(_12595_),
    .B1(_12600_),
    .Y(_12601_));
 sky130_fd_sc_hd__buf_1 _34642_ (.A(_07717_),
    .X(_12602_));
 sky130_fd_sc_hd__nand3_2 _34643_ (.A(_08790_),
    .B(_09617_),
    .C(_07798_),
    .Y(_12603_));
 sky130_fd_sc_hd__a22o_2 _34644_ (.A1(_08382_),
    .A2(_07143_),
    .B1(_09617_),
    .B2(_06748_),
    .X(_12604_));
 sky130_fd_sc_hd__o21ai_2 _34645_ (.A1(_06401_),
    .A2(_12603_),
    .B1(_12604_),
    .Y(_12605_));
 sky130_fd_sc_hd__o21ai_2 _34646_ (.A1(_12602_),
    .A2(_10279_),
    .B1(_12605_),
    .Y(_12606_));
 sky130_fd_sc_hd__nor2_2 _34647_ (.A(_07718_),
    .B(_08053_),
    .Y(_12607_));
 sky130_fd_sc_hd__o211ai_2 _34648_ (.A1(_06397_),
    .A2(_12603_),
    .B1(_12604_),
    .C1(_12607_),
    .Y(_12608_));
 sky130_fd_sc_hd__nand2_2 _34649_ (.A(_12281_),
    .B(_12275_),
    .Y(_12609_));
 sky130_fd_sc_hd__a21o_2 _34650_ (.A1(_12606_),
    .A2(_12608_),
    .B1(_12609_),
    .X(_12610_));
 sky130_fd_sc_hd__nand3_2 _34651_ (.A(_12606_),
    .B(_12609_),
    .C(_12608_),
    .Y(_12611_));
 sky130_fd_sc_hd__nand3b_2 _34652_ (.A_N(_12601_),
    .B(_12610_),
    .C(_12611_),
    .Y(_12612_));
 sky130_fd_sc_hd__a21oi_2 _34653_ (.A1(_12606_),
    .A2(_12608_),
    .B1(_12609_),
    .Y(_12613_));
 sky130_fd_sc_hd__and3_2 _34654_ (.A(_12606_),
    .B(_12609_),
    .C(_12608_),
    .X(_12614_));
 sky130_fd_sc_hd__o21ai_2 _34655_ (.A1(_12613_),
    .A2(_12614_),
    .B1(_12601_),
    .Y(_12615_));
 sky130_fd_sc_hd__o211ai_2 _34656_ (.A1(_12590_),
    .A2(_12591_),
    .B1(_12612_),
    .C1(_12615_),
    .Y(_12616_));
 sky130_fd_sc_hd__o21bai_2 _34657_ (.A1(_12613_),
    .A2(_12614_),
    .B1_N(_12601_),
    .Y(_12617_));
 sky130_fd_sc_hd__a21boi_2 _34658_ (.A1(_12256_),
    .A2(_12257_),
    .B1_N(_12253_),
    .Y(_12618_));
 sky130_fd_sc_hd__nand3_2 _34659_ (.A(_12610_),
    .B(_12611_),
    .C(_12601_),
    .Y(_12619_));
 sky130_fd_sc_hd__nand3_2 _34660_ (.A(_12617_),
    .B(_12618_),
    .C(_12619_),
    .Y(_12620_));
 sky130_fd_sc_hd__a21bo_2 _34661_ (.A1(_12295_),
    .A2(_12284_),
    .B1_N(_12279_),
    .X(_12621_));
 sky130_fd_sc_hd__a21oi_2 _34662_ (.A1(_12616_),
    .A2(_12620_),
    .B1(_12621_),
    .Y(_12622_));
 sky130_fd_sc_hd__and3_2 _34663_ (.A(_12616_),
    .B(_12620_),
    .C(_12621_),
    .X(_12623_));
 sky130_fd_sc_hd__nor2_2 _34664_ (.A(_12622_),
    .B(_12623_),
    .Y(_12624_));
 sky130_fd_sc_hd__nand3_2 _34665_ (.A(_12582_),
    .B(_12588_),
    .C(_12587_),
    .Y(_12625_));
 sky130_fd_sc_hd__nand2_2 _34666_ (.A(_12624_),
    .B(_12625_),
    .Y(_12626_));
 sky130_fd_sc_hd__a21oi_2 _34667_ (.A1(_12260_),
    .A2(_12262_),
    .B1(_12205_),
    .Y(_12627_));
 sky130_fd_sc_hd__o21ai_2 _34668_ (.A1(_12318_),
    .A2(_12627_),
    .B1(_12263_),
    .Y(_12628_));
 sky130_fd_sc_hd__nand2_2 _34669_ (.A(_12242_),
    .B(_12261_),
    .Y(_12629_));
 sky130_fd_sc_hd__nand2_2 _34670_ (.A(_12629_),
    .B(_12237_),
    .Y(_12630_));
 sky130_fd_sc_hd__o2bb2ai_2 _34671_ (.A1_N(_12559_),
    .A2_N(_12552_),
    .B1(_12580_),
    .B2(_12578_),
    .Y(_12631_));
 sky130_fd_sc_hd__nand3_2 _34672_ (.A(_12552_),
    .B(_12559_),
    .C(_12581_),
    .Y(_12632_));
 sky130_fd_sc_hd__nand3_2 _34673_ (.A(_12630_),
    .B(_12631_),
    .C(_12632_),
    .Y(_12633_));
 sky130_fd_sc_hd__nand2_2 _34674_ (.A(_12625_),
    .B(_12633_),
    .Y(_12634_));
 sky130_fd_sc_hd__a21o_2 _34675_ (.A1(_12616_),
    .A2(_12620_),
    .B1(_12621_),
    .X(_12635_));
 sky130_fd_sc_hd__nand3_2 _34676_ (.A(_12616_),
    .B(_12620_),
    .C(_12621_),
    .Y(_12636_));
 sky130_fd_sc_hd__nand2_2 _34677_ (.A(_12635_),
    .B(_12636_),
    .Y(_12637_));
 sky130_fd_sc_hd__nand2_2 _34678_ (.A(_12634_),
    .B(_12637_),
    .Y(_12638_));
 sky130_fd_sc_hd__o211ai_2 _34679_ (.A1(_12589_),
    .A2(_12626_),
    .B1(_12628_),
    .C1(_12638_),
    .Y(_12639_));
 sky130_fd_sc_hd__nand2_2 _34680_ (.A(_12634_),
    .B(_12624_),
    .Y(_12640_));
 sky130_fd_sc_hd__a21boi_2 _34681_ (.A1(_12311_),
    .A2(_12268_),
    .B1_N(_12263_),
    .Y(_12641_));
 sky130_fd_sc_hd__nand3_2 _34682_ (.A(_12625_),
    .B(_12633_),
    .C(_12637_),
    .Y(_12642_));
 sky130_fd_sc_hd__nand3_2 _34683_ (.A(_12640_),
    .B(_12641_),
    .C(_12642_),
    .Y(_12643_));
 sky130_fd_sc_hd__nand2_2 _34684_ (.A(_07886_),
    .B(_07590_),
    .Y(_12644_));
 sky130_fd_sc_hd__nand2_2 _34685_ (.A(_06828_),
    .B(_09250_),
    .Y(_12645_));
 sky130_fd_sc_hd__nor2_2 _34686_ (.A(_12644_),
    .B(_12645_),
    .Y(_12646_));
 sky130_fd_sc_hd__and2_2 _34687_ (.A(_12644_),
    .B(_12645_),
    .X(_12647_));
 sky130_fd_sc_hd__nand2_2 _34688_ (.A(_19359_),
    .B(_19573_),
    .Y(_12648_));
 sky130_fd_sc_hd__o21ai_2 _34689_ (.A1(_12646_),
    .A2(_12647_),
    .B1(_12648_),
    .Y(_12649_));
 sky130_fd_sc_hd__nand2_2 _34690_ (.A(_12286_),
    .B(_12287_),
    .Y(_12650_));
 sky130_fd_sc_hd__a31o_2 _34691_ (.A1(_12650_),
    .A2(_12069_),
    .A3(_19586_),
    .B1(_12288_),
    .X(_12651_));
 sky130_fd_sc_hd__nand2_2 _34692_ (.A(_12644_),
    .B(_12645_),
    .Y(_12652_));
 sky130_fd_sc_hd__inv_2 _34693_ (.A(_12648_),
    .Y(_12653_));
 sky130_fd_sc_hd__nand3b_2 _34694_ (.A_N(_12646_),
    .B(_12652_),
    .C(_12653_),
    .Y(_12654_));
 sky130_fd_sc_hd__nand3_2 _34695_ (.A(_12649_),
    .B(_12651_),
    .C(_12654_),
    .Y(_12655_));
 sky130_fd_sc_hd__o21ai_2 _34696_ (.A1(_12646_),
    .A2(_12647_),
    .B1(_12653_),
    .Y(_12656_));
 sky130_fd_sc_hd__nand3b_2 _34697_ (.A_N(_12646_),
    .B(_12652_),
    .C(_12648_),
    .Y(_12657_));
 sky130_fd_sc_hd__a21oi_2 _34698_ (.A1(_12289_),
    .A2(_12650_),
    .B1(_12288_),
    .Y(_12658_));
 sky130_fd_sc_hd__nand3_2 _34699_ (.A(_12656_),
    .B(_12657_),
    .C(_12658_),
    .Y(_12659_));
 sky130_fd_sc_hd__a21o_2 _34700_ (.A1(_12334_),
    .A2(_12335_),
    .B1(_12329_),
    .X(_12660_));
 sky130_fd_sc_hd__a21o_2 _34701_ (.A1(_12655_),
    .A2(_12659_),
    .B1(_12660_),
    .X(_12661_));
 sky130_fd_sc_hd__nand3_2 _34702_ (.A(_12655_),
    .B(_12659_),
    .C(_12660_),
    .Y(_12662_));
 sky130_fd_sc_hd__nand2_2 _34703_ (.A(_12341_),
    .B(_12342_),
    .Y(_12663_));
 sky130_fd_sc_hd__nand2_2 _34704_ (.A(_12663_),
    .B(_12337_),
    .Y(_12664_));
 sky130_fd_sc_hd__a21oi_2 _34705_ (.A1(_12661_),
    .A2(_12662_),
    .B1(_12664_),
    .Y(_12665_));
 sky130_fd_sc_hd__inv_2 _34706_ (.A(_12655_),
    .Y(_12666_));
 sky130_fd_sc_hd__nand2_2 _34707_ (.A(_12659_),
    .B(_12660_),
    .Y(_12667_));
 sky130_fd_sc_hd__o211a_2 _34708_ (.A1(_12666_),
    .A2(_12667_),
    .B1(_12664_),
    .C1(_12661_),
    .X(_12668_));
 sky130_fd_sc_hd__a21oi_2 _34709_ (.A1(_12350_),
    .A2(_12354_),
    .B1(_12348_),
    .Y(_12669_));
 sky130_fd_sc_hd__nand2_2 _34710_ (.A(_19363_),
    .B(_19570_),
    .Y(_12670_));
 sky130_fd_sc_hd__nand2_2 _34711_ (.A(_07450_),
    .B(_19567_),
    .Y(_12671_));
 sky130_fd_sc_hd__nor2_2 _34712_ (.A(_12670_),
    .B(_12671_),
    .Y(_12672_));
 sky130_fd_sc_hd__and2_2 _34713_ (.A(_12670_),
    .B(_12671_),
    .X(_12673_));
 sky130_fd_sc_hd__nand2_2 _34714_ (.A(_06628_),
    .B(_19564_),
    .Y(_12674_));
 sky130_fd_sc_hd__o21ai_2 _34715_ (.A1(_12672_),
    .A2(_12673_),
    .B1(_12674_),
    .Y(_12675_));
 sky130_fd_sc_hd__nand2_2 _34716_ (.A(_12670_),
    .B(_12671_),
    .Y(_12676_));
 sky130_fd_sc_hd__inv_2 _34717_ (.A(_12674_),
    .Y(_12677_));
 sky130_fd_sc_hd__nand3b_2 _34718_ (.A_N(_12672_),
    .B(_12676_),
    .C(_12677_),
    .Y(_12678_));
 sky130_fd_sc_hd__nand3b_2 _34719_ (.A_N(_12669_),
    .B(_12675_),
    .C(_12678_),
    .Y(_12679_));
 sky130_fd_sc_hd__inv_2 _34720_ (.A(_12679_),
    .Y(_12680_));
 sky130_fd_sc_hd__nand2_2 _34721_ (.A(_12675_),
    .B(_12678_),
    .Y(_12681_));
 sky130_fd_sc_hd__nand2_2 _34722_ (.A(_05807_),
    .B(_08905_),
    .Y(_12682_));
 sky130_fd_sc_hd__nand2_2 _34723_ (.A(_08331_),
    .B(_09736_),
    .Y(_12683_));
 sky130_fd_sc_hd__nor2_2 _34724_ (.A(_12682_),
    .B(_12683_),
    .Y(_12684_));
 sky130_fd_sc_hd__nand2_2 _34725_ (.A(_12682_),
    .B(_12683_),
    .Y(_12685_));
 sky130_fd_sc_hd__or2b_2 _34726_ (.A(_12684_),
    .B_N(_12685_),
    .X(_12686_));
 sky130_fd_sc_hd__nor2_2 _34727_ (.A(_05498_),
    .B(_10542_),
    .Y(_12687_));
 sky130_fd_sc_hd__nand2_2 _34728_ (.A(_12686_),
    .B(_12687_),
    .Y(_12688_));
 sky130_fd_sc_hd__and2b_2 _34729_ (.A_N(_12684_),
    .B(_12685_),
    .X(_12689_));
 sky130_fd_sc_hd__o21ai_2 _34730_ (.A1(_05498_),
    .A2(_10543_),
    .B1(_12689_),
    .Y(_12690_));
 sky130_fd_sc_hd__a22o_2 _34731_ (.A1(_12681_),
    .A2(_12669_),
    .B1(_12688_),
    .B2(_12690_),
    .X(_12691_));
 sky130_fd_sc_hd__nand2_2 _34732_ (.A(_12681_),
    .B(_12669_),
    .Y(_12692_));
 sky130_fd_sc_hd__nand2_2 _34733_ (.A(_12690_),
    .B(_12688_),
    .Y(_12693_));
 sky130_fd_sc_hd__a21o_2 _34734_ (.A1(_12692_),
    .A2(_12679_),
    .B1(_12693_),
    .X(_12694_));
 sky130_fd_sc_hd__o21ai_2 _34735_ (.A1(_12680_),
    .A2(_12691_),
    .B1(_12694_),
    .Y(_12695_));
 sky130_fd_sc_hd__o21ai_2 _34736_ (.A1(_12665_),
    .A2(_12668_),
    .B1(_12695_),
    .Y(_12696_));
 sky130_fd_sc_hd__o21ai_2 _34737_ (.A1(_12305_),
    .A2(_12316_),
    .B1(_12300_),
    .Y(_12697_));
 sky130_fd_sc_hd__o21a_2 _34738_ (.A1(_12680_),
    .A2(_12691_),
    .B1(_12694_),
    .X(_12698_));
 sky130_fd_sc_hd__a21o_2 _34739_ (.A1(_12661_),
    .A2(_12662_),
    .B1(_12664_),
    .X(_12699_));
 sky130_fd_sc_hd__nand3_2 _34740_ (.A(_12661_),
    .B(_12664_),
    .C(_12662_),
    .Y(_12700_));
 sky130_fd_sc_hd__nand3_2 _34741_ (.A(_12698_),
    .B(_12699_),
    .C(_12700_),
    .Y(_12701_));
 sky130_fd_sc_hd__nand3_2 _34742_ (.A(_12696_),
    .B(_12697_),
    .C(_12701_),
    .Y(_12702_));
 sky130_fd_sc_hd__o21ai_2 _34743_ (.A1(_12665_),
    .A2(_12668_),
    .B1(_12698_),
    .Y(_12703_));
 sky130_fd_sc_hd__nand2_2 _34744_ (.A(_12305_),
    .B(_12300_),
    .Y(_12704_));
 sky130_fd_sc_hd__nand2_2 _34745_ (.A(_12704_),
    .B(_12299_),
    .Y(_12705_));
 sky130_fd_sc_hd__nand3_2 _34746_ (.A(_12699_),
    .B(_12695_),
    .C(_12700_),
    .Y(_12706_));
 sky130_fd_sc_hd__a32oi_2 _34747_ (.A1(_12703_),
    .A2(_12705_),
    .A3(_12706_),
    .B1(_12383_),
    .B2(_12374_),
    .Y(_12707_));
 sky130_fd_sc_hd__nand3_2 _34748_ (.A(_12703_),
    .B(_12705_),
    .C(_12706_),
    .Y(_12708_));
 sky130_fd_sc_hd__nand2_2 _34749_ (.A(_12374_),
    .B(_12383_),
    .Y(_12709_));
 sky130_fd_sc_hd__a21oi_2 _34750_ (.A1(_12702_),
    .A2(_12708_),
    .B1(_12709_),
    .Y(_12710_));
 sky130_fd_sc_hd__a21o_2 _34751_ (.A1(_12702_),
    .A2(_12707_),
    .B1(_12710_),
    .X(_12711_));
 sky130_fd_sc_hd__a21o_2 _34752_ (.A1(_12639_),
    .A2(_12643_),
    .B1(_12711_),
    .X(_12712_));
 sky130_fd_sc_hd__a21boi_2 _34753_ (.A1(_12392_),
    .A2(_12323_),
    .B1_N(_12313_),
    .Y(_12713_));
 sky130_fd_sc_hd__nand3_2 _34754_ (.A(_12711_),
    .B(_12639_),
    .C(_12643_),
    .Y(_12714_));
 sky130_fd_sc_hd__nand3_2 _34755_ (.A(_12712_),
    .B(_12713_),
    .C(_12714_),
    .Y(_12715_));
 sky130_fd_sc_hd__a21oi_2 _34756_ (.A1(_12308_),
    .A2(_12312_),
    .B1(_12203_),
    .Y(_12716_));
 sky130_fd_sc_hd__o21ai_2 _34757_ (.A1(_12397_),
    .A2(_12716_),
    .B1(_12313_),
    .Y(_12717_));
 sky130_fd_sc_hd__nand2_2 _34758_ (.A(_12707_),
    .B(_12702_),
    .Y(_12718_));
 sky130_fd_sc_hd__inv_2 _34759_ (.A(_12718_),
    .Y(_12719_));
 sky130_fd_sc_hd__o2bb2ai_2 _34760_ (.A1_N(_12643_),
    .A2_N(_12639_),
    .B1(_12710_),
    .B2(_12719_),
    .Y(_12720_));
 sky130_fd_sc_hd__a21oi_2 _34761_ (.A1(_12702_),
    .A2(_12707_),
    .B1(_12710_),
    .Y(_12721_));
 sky130_fd_sc_hd__nand3_2 _34762_ (.A(_12639_),
    .B(_12643_),
    .C(_12721_),
    .Y(_12722_));
 sky130_fd_sc_hd__nand3_2 _34763_ (.A(_12717_),
    .B(_12720_),
    .C(_12722_),
    .Y(_12723_));
 sky130_fd_sc_hd__nand2_2 _34764_ (.A(_12715_),
    .B(_12723_),
    .Y(_12724_));
 sky130_fd_sc_hd__nand2_2 _34765_ (.A(_12462_),
    .B(_12430_),
    .Y(_12725_));
 sky130_fd_sc_hd__inv_2 _34766_ (.A(_12725_),
    .Y(_12726_));
 sky130_fd_sc_hd__a21o_2 _34767_ (.A1(_12436_),
    .A2(_12437_),
    .B1(_04836_),
    .X(_12727_));
 sky130_fd_sc_hd__nand2_2 _34768_ (.A(_12727_),
    .B(_12438_),
    .Y(_12728_));
 sky130_fd_sc_hd__o21ai_2 _34769_ (.A1(_19389_),
    .A2(_19392_),
    .B1(_11429_),
    .Y(_12729_));
 sky130_fd_sc_hd__and3_2 _34770_ (.A(_11429_),
    .B(_05712_),
    .C(_05892_),
    .X(_12730_));
 sky130_fd_sc_hd__nor2_2 _34771_ (.A(_12729_),
    .B(_12730_),
    .Y(_12731_));
 sky130_fd_sc_hd__nand2_2 _34772_ (.A(_12728_),
    .B(_12731_),
    .Y(_12732_));
 sky130_fd_sc_hd__nand3b_2 _34773_ (.A_N(_12731_),
    .B(_12438_),
    .C(_12727_),
    .Y(_12733_));
 sky130_fd_sc_hd__a21o_2 _34774_ (.A1(_12732_),
    .A2(_12733_),
    .B1(_11919_),
    .X(_12734_));
 sky130_fd_sc_hd__nand3_2 _34775_ (.A(_11918_),
    .B(_12732_),
    .C(_12733_),
    .Y(_12735_));
 sky130_fd_sc_hd__a22o_2 _34776_ (.A1(_12446_),
    .A2(_12448_),
    .B1(_12734_),
    .B2(_12735_),
    .X(_12736_));
 sky130_fd_sc_hd__nand2_2 _34777_ (.A(_12446_),
    .B(_12448_),
    .Y(_12737_));
 sky130_fd_sc_hd__nand3b_2 _34778_ (.A_N(_12737_),
    .B(_12734_),
    .C(_12735_),
    .Y(_12738_));
 sky130_fd_sc_hd__nand2_2 _34779_ (.A(_12736_),
    .B(_12738_),
    .Y(_12739_));
 sky130_fd_sc_hd__and2_2 _34780_ (.A(_12739_),
    .B(_12456_),
    .X(_12740_));
 sky130_fd_sc_hd__nor2_2 _34781_ (.A(_12456_),
    .B(_12739_),
    .Y(_12741_));
 sky130_fd_sc_hd__and4_2 _34782_ (.A(_07797_),
    .B(_08949_),
    .C(_10537_),
    .D(_10538_),
    .X(_12742_));
 sky130_fd_sc_hd__inv_2 _34783_ (.A(_07797_),
    .Y(_12743_));
 sky130_fd_sc_hd__nand2_2 _34784_ (.A(_09254_),
    .B(_10537_),
    .Y(_12744_));
 sky130_fd_sc_hd__o21a_2 _34785_ (.A1(_12743_),
    .A2(_10533_),
    .B1(_12744_),
    .X(_12745_));
 sky130_fd_sc_hd__nand2_2 _34786_ (.A(_08953_),
    .B(_11901_),
    .Y(_12746_));
 sky130_fd_sc_hd__o21ai_2 _34787_ (.A1(_12742_),
    .A2(_12745_),
    .B1(_12746_),
    .Y(_12747_));
 sky130_fd_sc_hd__a21o_2 _34788_ (.A1(_12365_),
    .A2(_12362_),
    .B1(_12361_),
    .X(_12748_));
 sky130_fd_sc_hd__o21ai_2 _34789_ (.A1(_12743_),
    .A2(_10533_),
    .B1(_12744_),
    .Y(_12749_));
 sky130_fd_sc_hd__inv_2 _34790_ (.A(_12746_),
    .Y(_12750_));
 sky130_fd_sc_hd__nand3b_2 _34791_ (.A_N(_12742_),
    .B(_12749_),
    .C(_12750_),
    .Y(_12751_));
 sky130_fd_sc_hd__nand3_2 _34792_ (.A(_12747_),
    .B(_12748_),
    .C(_12751_),
    .Y(_12752_));
 sky130_fd_sc_hd__o21ai_2 _34793_ (.A1(_12742_),
    .A2(_12745_),
    .B1(_12750_),
    .Y(_12753_));
 sky130_fd_sc_hd__a21oi_2 _34794_ (.A1(_12365_),
    .A2(_12362_),
    .B1(_12361_),
    .Y(_12754_));
 sky130_fd_sc_hd__nand3b_2 _34795_ (.A_N(_12742_),
    .B(_12749_),
    .C(_12746_),
    .Y(_12755_));
 sky130_fd_sc_hd__nand3_2 _34796_ (.A(_12753_),
    .B(_12754_),
    .C(_12755_),
    .Y(_12756_));
 sky130_fd_sc_hd__nand2_2 _34797_ (.A(_12752_),
    .B(_12756_),
    .Y(_12757_));
 sky130_fd_sc_hd__a21oi_2 _34798_ (.A1(_12410_),
    .A2(_12409_),
    .B1(_12405_),
    .Y(_12758_));
 sky130_fd_sc_hd__nand2_2 _34799_ (.A(_12757_),
    .B(_12758_),
    .Y(_12759_));
 sky130_fd_sc_hd__nand3b_2 _34800_ (.A_N(_12758_),
    .B(_12752_),
    .C(_12756_),
    .Y(_12760_));
 sky130_fd_sc_hd__nand2_2 _34801_ (.A(_12370_),
    .B(_12357_),
    .Y(_12761_));
 sky130_fd_sc_hd__a21oi_2 _34802_ (.A1(_12759_),
    .A2(_12760_),
    .B1(_12761_),
    .Y(_12762_));
 sky130_fd_sc_hd__and3_2 _34803_ (.A(_12759_),
    .B(_12761_),
    .C(_12760_),
    .X(_12763_));
 sky130_fd_sc_hd__inv_2 _34804_ (.A(_12415_),
    .Y(_12764_));
 sky130_fd_sc_hd__o21a_2 _34805_ (.A1(_12416_),
    .A2(_12764_),
    .B1(_12412_),
    .X(_12765_));
 sky130_fd_sc_hd__o21ai_2 _34806_ (.A1(_12762_),
    .A2(_12763_),
    .B1(_12765_),
    .Y(_12766_));
 sky130_fd_sc_hd__nand2_2 _34807_ (.A(_12759_),
    .B(_12760_),
    .Y(_12767_));
 sky130_fd_sc_hd__and2_2 _34808_ (.A(_12370_),
    .B(_12357_),
    .X(_12768_));
 sky130_fd_sc_hd__nand2_2 _34809_ (.A(_12767_),
    .B(_12768_),
    .Y(_12769_));
 sky130_fd_sc_hd__nand3_2 _34810_ (.A(_12759_),
    .B(_12761_),
    .C(_12760_),
    .Y(_12770_));
 sky130_fd_sc_hd__nand3b_2 _34811_ (.A_N(_12765_),
    .B(_12769_),
    .C(_12770_),
    .Y(_12771_));
 sky130_fd_sc_hd__o21ai_2 _34812_ (.A1(_12432_),
    .A2(_12433_),
    .B1(_12425_),
    .Y(_12772_));
 sky130_fd_sc_hd__a21oi_2 _34813_ (.A1(_12766_),
    .A2(_12771_),
    .B1(_12772_),
    .Y(_12773_));
 sky130_fd_sc_hd__and3_2 _34814_ (.A(_12766_),
    .B(_12771_),
    .C(_12772_),
    .X(_12774_));
 sky130_fd_sc_hd__o22ai_2 _34815_ (.A1(_12740_),
    .A2(_12741_),
    .B1(_12773_),
    .B2(_12774_),
    .Y(_12775_));
 sky130_fd_sc_hd__a21o_2 _34816_ (.A1(_12766_),
    .A2(_12771_),
    .B1(_12772_),
    .X(_12776_));
 sky130_fd_sc_hd__nand3_2 _34817_ (.A(_12766_),
    .B(_12772_),
    .C(_12771_),
    .Y(_12777_));
 sky130_fd_sc_hd__o2bb2ai_2 _34818_ (.A1_N(_12736_),
    .A2_N(_12738_),
    .B1(_11761_),
    .B2(_11916_),
    .Y(_12778_));
 sky130_fd_sc_hd__nand3_2 _34819_ (.A(_12736_),
    .B(_12738_),
    .C(_12456_),
    .Y(_12779_));
 sky130_fd_sc_hd__nand2_2 _34820_ (.A(_12778_),
    .B(_12779_),
    .Y(_12780_));
 sky130_fd_sc_hd__nand3_2 _34821_ (.A(_12776_),
    .B(_12777_),
    .C(_12780_),
    .Y(_12781_));
 sky130_fd_sc_hd__nand2_2 _34822_ (.A(_12385_),
    .B(_12388_),
    .Y(_12782_));
 sky130_fd_sc_hd__nand2_2 _34823_ (.A(_12782_),
    .B(_12380_),
    .Y(_12783_));
 sky130_fd_sc_hd__a21oi_2 _34824_ (.A1(_12775_),
    .A2(_12781_),
    .B1(_12783_),
    .Y(_12784_));
 sky130_fd_sc_hd__nor2_2 _34825_ (.A(_12726_),
    .B(_12784_),
    .Y(_12785_));
 sky130_fd_sc_hd__nand3_2 _34826_ (.A(_12775_),
    .B(_12783_),
    .C(_12781_),
    .Y(_12786_));
 sky130_fd_sc_hd__nand2_2 _34827_ (.A(_12777_),
    .B(_12780_),
    .Y(_12787_));
 sky130_fd_sc_hd__nor2_2 _34828_ (.A(_12773_),
    .B(_12787_),
    .Y(_12788_));
 sky130_fd_sc_hd__a21oi_2 _34829_ (.A1(_12776_),
    .A2(_12777_),
    .B1(_12780_),
    .Y(_12789_));
 sky130_fd_sc_hd__o21bai_2 _34830_ (.A1(_12788_),
    .A2(_12789_),
    .B1_N(_12783_),
    .Y(_12790_));
 sky130_fd_sc_hd__a21oi_2 _34831_ (.A1(_12790_),
    .A2(_12786_),
    .B1(_12725_),
    .Y(_12791_));
 sky130_fd_sc_hd__a21oi_2 _34832_ (.A1(_12785_),
    .A2(_12786_),
    .B1(_12791_),
    .Y(_12792_));
 sky130_fd_sc_hd__nand2_2 _34833_ (.A(_12724_),
    .B(_12792_),
    .Y(_12793_));
 sky130_fd_sc_hd__and3_2 _34834_ (.A(_12775_),
    .B(_12781_),
    .C(_12783_),
    .X(_12794_));
 sky130_fd_sc_hd__o21ai_2 _34835_ (.A1(_12784_),
    .A2(_12794_),
    .B1(_12726_),
    .Y(_12795_));
 sky130_fd_sc_hd__nand3_2 _34836_ (.A(_12790_),
    .B(_12725_),
    .C(_12786_),
    .Y(_12796_));
 sky130_fd_sc_hd__nand2_2 _34837_ (.A(_12795_),
    .B(_12796_),
    .Y(_12797_));
 sky130_fd_sc_hd__nand3_2 _34838_ (.A(_12797_),
    .B(_12715_),
    .C(_12723_),
    .Y(_12798_));
 sky130_fd_sc_hd__nand3_2 _34839_ (.A(_12523_),
    .B(_12793_),
    .C(_12798_),
    .Y(_12799_));
 sky130_fd_sc_hd__nand2_2 _34840_ (.A(_12483_),
    .B(_12394_),
    .Y(_12800_));
 sky130_fd_sc_hd__inv_2 _34841_ (.A(_12796_),
    .Y(_12801_));
 sky130_fd_sc_hd__o2bb2ai_2 _34842_ (.A1_N(_12723_),
    .A2_N(_12715_),
    .B1(_12791_),
    .B2(_12801_),
    .Y(_12802_));
 sky130_fd_sc_hd__nand2_2 _34843_ (.A(_12790_),
    .B(_12725_),
    .Y(_12803_));
 sky130_fd_sc_hd__o2111ai_2 _34844_ (.A1(_12794_),
    .A2(_12803_),
    .B1(_12795_),
    .C1(_12723_),
    .D1(_12715_),
    .Y(_12804_));
 sky130_fd_sc_hd__nand3_2 _34845_ (.A(_12800_),
    .B(_12802_),
    .C(_12804_),
    .Y(_12805_));
 sky130_fd_sc_hd__nand2_2 _34846_ (.A(_12472_),
    .B(_12466_),
    .Y(_12806_));
 sky130_fd_sc_hd__and2_2 _34847_ (.A(_12452_),
    .B(_12457_),
    .X(_12807_));
 sky130_fd_sc_hd__inv_2 _34848_ (.A(_12807_),
    .Y(_12808_));
 sky130_fd_sc_hd__nand2_2 _34849_ (.A(_12808_),
    .B(_12454_),
    .Y(_12809_));
 sky130_fd_sc_hd__nand2_2 _34850_ (.A(_12806_),
    .B(_12809_),
    .Y(_12810_));
 sky130_fd_sc_hd__inv_2 _34851_ (.A(_12809_),
    .Y(_12811_));
 sky130_fd_sc_hd__nand3_2 _34852_ (.A(_12472_),
    .B(_12466_),
    .C(_12811_),
    .Y(_12812_));
 sky130_fd_sc_hd__nand2_2 _34853_ (.A(_12810_),
    .B(_12812_),
    .Y(_12813_));
 sky130_fd_sc_hd__inv_2 _34854_ (.A(_12813_),
    .Y(_12814_));
 sky130_fd_sc_hd__a21o_2 _34855_ (.A1(_12799_),
    .A2(_12805_),
    .B1(_12814_),
    .X(_12815_));
 sky130_fd_sc_hd__o21ai_2 _34856_ (.A1(_12502_),
    .A2(_12480_),
    .B1(_12489_),
    .Y(_12816_));
 sky130_fd_sc_hd__nand3_2 _34857_ (.A(_12799_),
    .B(_12805_),
    .C(_12814_),
    .Y(_12817_));
 sky130_fd_sc_hd__nand3_2 _34858_ (.A(_12815_),
    .B(_12816_),
    .C(_12817_),
    .Y(_12818_));
 sky130_fd_sc_hd__a21oi_2 _34859_ (.A1(_12488_),
    .A2(_12490_),
    .B1(_12484_),
    .Y(_12819_));
 sky130_fd_sc_hd__inv_2 _34860_ (.A(_12806_),
    .Y(_12820_));
 sky130_fd_sc_hd__nor2_2 _34861_ (.A(_12809_),
    .B(_12820_),
    .Y(_12821_));
 sky130_fd_sc_hd__nor2_2 _34862_ (.A(_12811_),
    .B(_12806_),
    .Y(_12822_));
 sky130_fd_sc_hd__o2bb2ai_2 _34863_ (.A1_N(_12805_),
    .A2_N(_12799_),
    .B1(_12821_),
    .B2(_12822_),
    .Y(_12823_));
 sky130_fd_sc_hd__nand3_2 _34864_ (.A(_12799_),
    .B(_12805_),
    .C(_12813_),
    .Y(_12824_));
 sky130_fd_sc_hd__nand3_2 _34865_ (.A(_12819_),
    .B(_12823_),
    .C(_12824_),
    .Y(_12825_));
 sky130_fd_sc_hd__inv_2 _34866_ (.A(_12194_),
    .Y(_12826_));
 sky130_fd_sc_hd__nand3_2 _34867_ (.A(_12818_),
    .B(_12825_),
    .C(_12826_),
    .Y(_12827_));
 sky130_fd_sc_hd__a21o_2 _34868_ (.A1(_12818_),
    .A2(_12825_),
    .B1(_12826_),
    .X(_12828_));
 sky130_fd_sc_hd__nand3b_2 _34869_ (.A_N(_12522_),
    .B(_12827_),
    .C(_12828_),
    .Y(_12829_));
 sky130_fd_sc_hd__o2bb2ai_2 _34870_ (.A1_N(_12825_),
    .A2_N(_12818_),
    .B1(_12191_),
    .B2(_12193_),
    .Y(_12830_));
 sky130_fd_sc_hd__nand3_2 _34871_ (.A(_12818_),
    .B(_12825_),
    .C(_12194_),
    .Y(_12831_));
 sky130_fd_sc_hd__nand3_2 _34872_ (.A(_12830_),
    .B(_12522_),
    .C(_12831_),
    .Y(_12832_));
 sky130_fd_sc_hd__and2_2 _34873_ (.A(_12829_),
    .B(_12832_),
    .X(_12833_));
 sky130_fd_sc_hd__nand3b_2 _34874_ (.A_N(_12519_),
    .B(_12511_),
    .C(_12833_),
    .Y(_12834_));
 sky130_fd_sc_hd__o21bai_2 _34875_ (.A1(_12512_),
    .A2(_12519_),
    .B1_N(_12833_),
    .Y(_12835_));
 sky130_fd_sc_hd__nand2_2 _34876_ (.A(_12834_),
    .B(_12835_),
    .Y(_02656_));
 sky130_fd_sc_hd__a21oi_2 _34877_ (.A1(_12823_),
    .A2(_12824_),
    .B1(_12819_),
    .Y(_12836_));
 sky130_fd_sc_hd__a31oi_2 _34878_ (.A1(_12819_),
    .A2(_12823_),
    .A3(_12824_),
    .B1(_12826_),
    .Y(_12837_));
 sky130_fd_sc_hd__a21oi_2 _34879_ (.A1(_12793_),
    .A2(_12798_),
    .B1(_12523_),
    .Y(_12838_));
 sky130_fd_sc_hd__a31oi_2 _34880_ (.A1(_12523_),
    .A2(_12793_),
    .A3(_12798_),
    .B1(_12813_),
    .Y(_12839_));
 sky130_fd_sc_hd__a21oi_2 _34881_ (.A1(_12712_),
    .A2(_12714_),
    .B1(_12713_),
    .Y(_12840_));
 sky130_fd_sc_hd__a31oi_2 _34882_ (.A1(_12715_),
    .A2(_12795_),
    .A3(_12796_),
    .B1(_12840_),
    .Y(_12841_));
 sky130_fd_sc_hd__nand2_2 _34883_ (.A(_12534_),
    .B(_12550_),
    .Y(_12842_));
 sky130_fd_sc_hd__nand2_2 _34884_ (.A(_12842_),
    .B(_12538_),
    .Y(_12843_));
 sky130_fd_sc_hd__o21ai_2 _34885_ (.A1(_19626_),
    .A2(_12524_),
    .B1(_12527_),
    .Y(_12844_));
 sky130_fd_sc_hd__nand2_2 _34886_ (.A(_12525_),
    .B(_12844_),
    .Y(_12845_));
 sky130_fd_sc_hd__nand2_2 _34887_ (.A(_19307_),
    .B(_06808_),
    .Y(_12846_));
 sky130_fd_sc_hd__nand3b_2 _34888_ (.A_N(_12846_),
    .B(_10824_),
    .C(_05261_),
    .Y(_12847_));
 sky130_fd_sc_hd__o21ai_2 _34889_ (.A1(_06614_),
    .A2(_11509_),
    .B1(_12846_),
    .Y(_12848_));
 sky130_fd_sc_hd__nand2_2 _34890_ (.A(_12847_),
    .B(_12848_),
    .Y(_12849_));
 sky130_fd_sc_hd__nand2_2 _34891_ (.A(_19311_),
    .B(_05613_),
    .Y(_12850_));
 sky130_fd_sc_hd__nand2_2 _34892_ (.A(_12849_),
    .B(_12850_),
    .Y(_12851_));
 sky130_fd_sc_hd__inv_2 _34893_ (.A(_12850_),
    .Y(_12852_));
 sky130_fd_sc_hd__nand3_2 _34894_ (.A(_12847_),
    .B(_12848_),
    .C(_12852_),
    .Y(_12853_));
 sky130_fd_sc_hd__nand3b_2 _34895_ (.A_N(_12845_),
    .B(_12851_),
    .C(_12853_),
    .Y(_12854_));
 sky130_fd_sc_hd__nand2_2 _34896_ (.A(_12849_),
    .B(_12852_),
    .Y(_12855_));
 sky130_fd_sc_hd__nand3_2 _34897_ (.A(_12847_),
    .B(_12848_),
    .C(_12850_),
    .Y(_12856_));
 sky130_fd_sc_hd__nand3_2 _34898_ (.A(_12855_),
    .B(_12856_),
    .C(_12845_),
    .Y(_12857_));
 sky130_fd_sc_hd__nor2_2 _34899_ (.A(_05735_),
    .B(_10704_),
    .Y(_12858_));
 sky130_fd_sc_hd__a22o_2 _34900_ (.A1(_19316_),
    .A2(_05615_),
    .B1(_10136_),
    .B2(_05738_),
    .X(_12859_));
 sky130_fd_sc_hd__nand2_2 _34901_ (.A(_19322_),
    .B(_19606_),
    .Y(_12860_));
 sky130_fd_sc_hd__inv_2 _34902_ (.A(_12860_),
    .Y(_12861_));
 sky130_fd_sc_hd__nand2_2 _34903_ (.A(_12859_),
    .B(_12861_),
    .Y(_12862_));
 sky130_fd_sc_hd__o21ai_2 _34904_ (.A1(_05735_),
    .A2(_11178_),
    .B1(_12859_),
    .Y(_12863_));
 sky130_fd_sc_hd__nand2_2 _34905_ (.A(_12863_),
    .B(_12860_),
    .Y(_12864_));
 sky130_fd_sc_hd__o21a_2 _34906_ (.A1(_12858_),
    .A2(_12862_),
    .B1(_12864_),
    .X(_12865_));
 sky130_fd_sc_hd__a21o_2 _34907_ (.A1(_12854_),
    .A2(_12857_),
    .B1(_12865_),
    .X(_12866_));
 sky130_fd_sc_hd__nand3_2 _34908_ (.A(_12854_),
    .B(_12865_),
    .C(_12857_),
    .Y(_12867_));
 sky130_fd_sc_hd__nand3_2 _34909_ (.A(_12843_),
    .B(_12866_),
    .C(_12867_),
    .Y(_12868_));
 sky130_fd_sc_hd__a21boi_2 _34910_ (.A1(_12534_),
    .A2(_12550_),
    .B1_N(_12538_),
    .Y(_12869_));
 sky130_fd_sc_hd__nand2_2 _34911_ (.A(_12854_),
    .B(_12857_),
    .Y(_12870_));
 sky130_fd_sc_hd__nand2_2 _34912_ (.A(_12870_),
    .B(_12865_),
    .Y(_12871_));
 sky130_fd_sc_hd__nand3b_2 _34913_ (.A_N(_12865_),
    .B(_12857_),
    .C(_12854_),
    .Y(_12872_));
 sky130_fd_sc_hd__nand3_2 _34914_ (.A(_12869_),
    .B(_12871_),
    .C(_12872_),
    .Y(_12873_));
 sky130_fd_sc_hd__nand2_2 _34915_ (.A(_12868_),
    .B(_12873_),
    .Y(_12874_));
 sky130_fd_sc_hd__o21ai_2 _34916_ (.A1(_05617_),
    .A2(_10705_),
    .B1(_12545_),
    .Y(_12875_));
 sky130_fd_sc_hd__nand2_2 _34917_ (.A(_09826_),
    .B(_07939_),
    .Y(_12876_));
 sky130_fd_sc_hd__nand2_2 _34918_ (.A(_10158_),
    .B(_19600_),
    .Y(_12877_));
 sky130_fd_sc_hd__nor2_2 _34919_ (.A(_12876_),
    .B(_12877_),
    .Y(_12878_));
 sky130_fd_sc_hd__and2_2 _34920_ (.A(_12876_),
    .B(_12877_),
    .X(_12879_));
 sky130_fd_sc_hd__nand2_2 _34921_ (.A(_19333_),
    .B(_08761_),
    .Y(_12880_));
 sky130_fd_sc_hd__o21ai_2 _34922_ (.A1(_12878_),
    .A2(_12879_),
    .B1(_12880_),
    .Y(_12881_));
 sky130_fd_sc_hd__nand2_2 _34923_ (.A(_12876_),
    .B(_12877_),
    .Y(_12882_));
 sky130_fd_sc_hd__inv_2 _34924_ (.A(_12880_),
    .Y(_12883_));
 sky130_fd_sc_hd__nand3b_2 _34925_ (.A_N(_12878_),
    .B(_12882_),
    .C(_12883_),
    .Y(_12884_));
 sky130_fd_sc_hd__nand3_2 _34926_ (.A(_12875_),
    .B(_12881_),
    .C(_12884_),
    .Y(_12885_));
 sky130_fd_sc_hd__o21ai_2 _34927_ (.A1(_12878_),
    .A2(_12879_),
    .B1(_12883_),
    .Y(_12886_));
 sky130_fd_sc_hd__nand3b_2 _34928_ (.A_N(_12878_),
    .B(_12882_),
    .C(_12880_),
    .Y(_12887_));
 sky130_fd_sc_hd__a21oi_2 _34929_ (.A1(_12539_),
    .A2(_12544_),
    .B1(_12541_),
    .Y(_12888_));
 sky130_fd_sc_hd__nand3_2 _34930_ (.A(_12886_),
    .B(_12887_),
    .C(_12888_),
    .Y(_12889_));
 sky130_fd_sc_hd__a21o_2 _34931_ (.A1(_12568_),
    .A2(_12567_),
    .B1(_12563_),
    .X(_12890_));
 sky130_fd_sc_hd__a21oi_2 _34932_ (.A1(_12885_),
    .A2(_12889_),
    .B1(_12890_),
    .Y(_12891_));
 sky130_fd_sc_hd__and3_2 _34933_ (.A(_12885_),
    .B(_12889_),
    .C(_12890_),
    .X(_12892_));
 sky130_fd_sc_hd__nor2_2 _34934_ (.A(_12891_),
    .B(_12892_),
    .Y(_12893_));
 sky130_fd_sc_hd__nand2_2 _34935_ (.A(_12874_),
    .B(_12893_),
    .Y(_12894_));
 sky130_fd_sc_hd__a21oi_2 _34936_ (.A1(_12556_),
    .A2(_12558_),
    .B1(_12557_),
    .Y(_12895_));
 sky130_fd_sc_hd__a21oi_2 _34937_ (.A1(_12559_),
    .A2(_12581_),
    .B1(_12895_),
    .Y(_12896_));
 sky130_fd_sc_hd__nand3b_2 _34938_ (.A_N(_12893_),
    .B(_12873_),
    .C(_12868_),
    .Y(_12897_));
 sky130_fd_sc_hd__nand3_2 _34939_ (.A(_12894_),
    .B(_12896_),
    .C(_12897_),
    .Y(_12898_));
 sky130_fd_sc_hd__a31oi_2 _34940_ (.A1(_12557_),
    .A2(_12556_),
    .A3(_12558_),
    .B1(_12586_),
    .Y(_12899_));
 sky130_fd_sc_hd__nand3_2 _34941_ (.A(_12868_),
    .B(_12873_),
    .C(_12893_),
    .Y(_12900_));
 sky130_fd_sc_hd__o2bb2ai_2 _34942_ (.A1_N(_12873_),
    .A2_N(_12868_),
    .B1(_12891_),
    .B2(_12892_),
    .Y(_12901_));
 sky130_fd_sc_hd__o211ai_2 _34943_ (.A1(_12895_),
    .A2(_12899_),
    .B1(_12900_),
    .C1(_12901_),
    .Y(_12902_));
 sky130_fd_sc_hd__nor2_2 _34944_ (.A(_07052_),
    .B(_09245_),
    .Y(_12903_));
 sky130_fd_sc_hd__a22oi_2 _34945_ (.A1(_07481_),
    .A2(_08950_),
    .B1(_07907_),
    .B2(_09933_),
    .Y(_12904_));
 sky130_fd_sc_hd__and4_2 _34946_ (.A(_07903_),
    .B(_07723_),
    .C(_07377_),
    .D(_08089_),
    .X(_12905_));
 sky130_fd_sc_hd__nor2_2 _34947_ (.A(_12904_),
    .B(_12905_),
    .Y(_12906_));
 sky130_fd_sc_hd__nor2_2 _34948_ (.A(_12903_),
    .B(_12906_),
    .Y(_12907_));
 sky130_fd_sc_hd__and2_2 _34949_ (.A(_12906_),
    .B(_12903_),
    .X(_12908_));
 sky130_fd_sc_hd__nand2_2 _34950_ (.A(_09094_),
    .B(_06957_),
    .Y(_12909_));
 sky130_fd_sc_hd__nand2_2 _34951_ (.A(_09614_),
    .B(_06949_),
    .Y(_12910_));
 sky130_fd_sc_hd__nor2_2 _34952_ (.A(_12909_),
    .B(_12910_),
    .Y(_12911_));
 sky130_fd_sc_hd__and2_2 _34953_ (.A(_12909_),
    .B(_12910_),
    .X(_12912_));
 sky130_fd_sc_hd__nand2_2 _34954_ (.A(_19342_),
    .B(_06951_),
    .Y(_12913_));
 sky130_fd_sc_hd__inv_2 _34955_ (.A(_12913_),
    .Y(_12914_));
 sky130_fd_sc_hd__o21ai_2 _34956_ (.A1(_12911_),
    .A2(_12912_),
    .B1(_12914_),
    .Y(_12915_));
 sky130_fd_sc_hd__nand2_2 _34957_ (.A(_12909_),
    .B(_12910_),
    .Y(_12916_));
 sky130_fd_sc_hd__nand3b_2 _34958_ (.A_N(_12911_),
    .B(_12916_),
    .C(_12913_),
    .Y(_12917_));
 sky130_fd_sc_hd__nor2_2 _34959_ (.A(_06401_),
    .B(_12603_),
    .Y(_12918_));
 sky130_fd_sc_hd__a21oi_2 _34960_ (.A1(_12607_),
    .A2(_12604_),
    .B1(_12918_),
    .Y(_12919_));
 sky130_fd_sc_hd__nand3_2 _34961_ (.A(_12915_),
    .B(_12917_),
    .C(_12919_),
    .Y(_12920_));
 sky130_fd_sc_hd__a21o_2 _34962_ (.A1(_12607_),
    .A2(_12604_),
    .B1(_12918_),
    .X(_12921_));
 sky130_fd_sc_hd__o21ai_2 _34963_ (.A1(_12911_),
    .A2(_12912_),
    .B1(_12913_),
    .Y(_12922_));
 sky130_fd_sc_hd__nand3b_2 _34964_ (.A_N(_12911_),
    .B(_12916_),
    .C(_12914_),
    .Y(_12923_));
 sky130_fd_sc_hd__nand3_2 _34965_ (.A(_12921_),
    .B(_12922_),
    .C(_12923_),
    .Y(_12924_));
 sky130_fd_sc_hd__o211ai_2 _34966_ (.A1(_12907_),
    .A2(_12908_),
    .B1(_12920_),
    .C1(_12924_),
    .Y(_12925_));
 sky130_fd_sc_hd__xor2_2 _34967_ (.A(_12903_),
    .B(_12906_),
    .X(_12926_));
 sky130_fd_sc_hd__nand2_2 _34968_ (.A(_12924_),
    .B(_12920_),
    .Y(_12927_));
 sky130_fd_sc_hd__nand2_2 _34969_ (.A(_12926_),
    .B(_12927_),
    .Y(_12928_));
 sky130_fd_sc_hd__inv_2 _34970_ (.A(_12584_),
    .Y(_12929_));
 sky130_fd_sc_hd__o2bb2a_2 _34971_ (.A1_N(_12925_),
    .A2_N(_12928_),
    .B1(_12583_),
    .B2(_12929_),
    .X(_12930_));
 sky130_fd_sc_hd__inv_2 _34972_ (.A(_12575_),
    .Y(_12931_));
 sky130_fd_sc_hd__a31oi_2 _34973_ (.A1(_12566_),
    .A2(_12570_),
    .A3(_12569_),
    .B1(_12577_),
    .Y(_12932_));
 sky130_fd_sc_hd__o211ai_2 _34974_ (.A1(_12931_),
    .A2(_12932_),
    .B1(_12925_),
    .C1(_12928_),
    .Y(_12933_));
 sky130_fd_sc_hd__o21ai_2 _34975_ (.A1(_12613_),
    .A2(_12601_),
    .B1(_12611_),
    .Y(_12934_));
 sky130_fd_sc_hd__nand2_2 _34976_ (.A(_12933_),
    .B(_12934_),
    .Y(_12935_));
 sky130_fd_sc_hd__o2bb2ai_2 _34977_ (.A1_N(_12925_),
    .A2_N(_12928_),
    .B1(_12583_),
    .B2(_12929_),
    .Y(_12936_));
 sky130_fd_sc_hd__a21o_2 _34978_ (.A1(_12936_),
    .A2(_12933_),
    .B1(_12934_),
    .X(_12937_));
 sky130_fd_sc_hd__o21ai_2 _34979_ (.A1(_12930_),
    .A2(_12935_),
    .B1(_12937_),
    .Y(_12938_));
 sky130_fd_sc_hd__a21o_2 _34980_ (.A1(_12898_),
    .A2(_12902_),
    .B1(_12938_),
    .X(_12939_));
 sky130_fd_sc_hd__a21oi_2 _34981_ (.A1(_12624_),
    .A2(_12625_),
    .B1(_12589_),
    .Y(_12940_));
 sky130_fd_sc_hd__nand3_2 _34982_ (.A(_12938_),
    .B(_12898_),
    .C(_12902_),
    .Y(_12941_));
 sky130_fd_sc_hd__nand3_2 _34983_ (.A(_12939_),
    .B(_12940_),
    .C(_12941_),
    .Y(_12942_));
 sky130_fd_sc_hd__a21oi_2 _34984_ (.A1(_12631_),
    .A2(_12632_),
    .B1(_12630_),
    .Y(_12943_));
 sky130_fd_sc_hd__o21ai_2 _34985_ (.A1(_12637_),
    .A2(_12943_),
    .B1(_12633_),
    .Y(_12944_));
 sky130_fd_sc_hd__nor2_2 _34986_ (.A(_12935_),
    .B(_12930_),
    .Y(_12945_));
 sky130_fd_sc_hd__a21oi_2 _34987_ (.A1(_12936_),
    .A2(_12933_),
    .B1(_12934_),
    .Y(_12946_));
 sky130_fd_sc_hd__o2bb2ai_2 _34988_ (.A1_N(_12902_),
    .A2_N(_12898_),
    .B1(_12945_),
    .B2(_12946_),
    .Y(_12947_));
 sky130_fd_sc_hd__nor2_2 _34989_ (.A(_12946_),
    .B(_12945_),
    .Y(_12948_));
 sky130_fd_sc_hd__nand3_2 _34990_ (.A(_12948_),
    .B(_12898_),
    .C(_12902_),
    .Y(_12949_));
 sky130_fd_sc_hd__nand3_2 _34991_ (.A(_12944_),
    .B(_12947_),
    .C(_12949_),
    .Y(_12950_));
 sky130_fd_sc_hd__nand2_2 _34992_ (.A(_12942_),
    .B(_12950_),
    .Y(_12951_));
 sky130_fd_sc_hd__a21oi_2 _34993_ (.A1(_12677_),
    .A2(_12676_),
    .B1(_12672_),
    .Y(_12952_));
 sky130_fd_sc_hd__nand2_2 _34994_ (.A(_07012_),
    .B(_08661_),
    .Y(_12953_));
 sky130_fd_sc_hd__nand2_2 _34995_ (.A(_06443_),
    .B(_08645_),
    .Y(_12954_));
 sky130_fd_sc_hd__nor2_2 _34996_ (.A(_12953_),
    .B(_12954_),
    .Y(_12955_));
 sky130_fd_sc_hd__and2_2 _34997_ (.A(_12953_),
    .B(_12954_),
    .X(_12956_));
 sky130_fd_sc_hd__nor2_2 _34998_ (.A(_06119_),
    .B(_10513_),
    .Y(_12957_));
 sky130_fd_sc_hd__o21bai_2 _34999_ (.A1(_12955_),
    .A2(_12956_),
    .B1_N(_12957_),
    .Y(_12958_));
 sky130_fd_sc_hd__nand2_2 _35000_ (.A(_12953_),
    .B(_12954_),
    .Y(_12959_));
 sky130_fd_sc_hd__nand3b_2 _35001_ (.A_N(_12955_),
    .B(_12957_),
    .C(_12959_),
    .Y(_12960_));
 sky130_fd_sc_hd__nand3b_2 _35002_ (.A_N(_12952_),
    .B(_12958_),
    .C(_12960_),
    .Y(_12961_));
 sky130_fd_sc_hd__inv_2 _35003_ (.A(_12961_),
    .Y(_12962_));
 sky130_fd_sc_hd__nand2_2 _35004_ (.A(_06500_),
    .B(_09203_),
    .Y(_12963_));
 sky130_fd_sc_hd__nand2_2 _35005_ (.A(_05670_),
    .B(_11410_),
    .Y(_12964_));
 sky130_fd_sc_hd__nor2_2 _35006_ (.A(_12963_),
    .B(_12964_),
    .Y(_12965_));
 sky130_fd_sc_hd__nand2_2 _35007_ (.A(_12963_),
    .B(_12964_),
    .Y(_12966_));
 sky130_fd_sc_hd__inv_2 _35008_ (.A(_12966_),
    .Y(_12967_));
 sky130_fd_sc_hd__nor2_2 _35009_ (.A(_05497_),
    .B(_10533_),
    .Y(_12968_));
 sky130_fd_sc_hd__o21bai_2 _35010_ (.A1(_12965_),
    .A2(_12967_),
    .B1_N(_12968_),
    .Y(_12969_));
 sky130_fd_sc_hd__nand3b_2 _35011_ (.A_N(_12965_),
    .B(_12968_),
    .C(_12966_),
    .Y(_12970_));
 sky130_fd_sc_hd__and2_2 _35012_ (.A(_12969_),
    .B(_12970_),
    .X(_12971_));
 sky130_fd_sc_hd__a21bo_2 _35013_ (.A1(_12958_),
    .A2(_12960_),
    .B1_N(_12952_),
    .X(_12972_));
 sky130_fd_sc_hd__nand2_2 _35014_ (.A(_12971_),
    .B(_12972_),
    .Y(_12973_));
 sky130_fd_sc_hd__nor2_2 _35015_ (.A(_12962_),
    .B(_12973_),
    .Y(_12974_));
 sky130_fd_sc_hd__a21oi_2 _35016_ (.A1(_12972_),
    .A2(_12961_),
    .B1(_12971_),
    .Y(_12975_));
 sky130_fd_sc_hd__a31o_2 _35017_ (.A1(_12649_),
    .A2(_12651_),
    .A3(_12654_),
    .B1(_12660_),
    .X(_12976_));
 sky130_fd_sc_hd__a21o_2 _35018_ (.A1(_12593_),
    .A2(_12594_),
    .B1(_12592_),
    .X(_12977_));
 sky130_fd_sc_hd__nand3_2 _35019_ (.A(_06821_),
    .B(_06827_),
    .C(_07837_),
    .Y(_12978_));
 sky130_fd_sc_hd__a22o_2 _35020_ (.A1(_06821_),
    .A2(_07605_),
    .B1(_06827_),
    .B2(_07837_),
    .X(_12979_));
 sky130_fd_sc_hd__o21ai_2 _35021_ (.A1(_09677_),
    .A2(_12978_),
    .B1(_12979_),
    .Y(_12980_));
 sky130_fd_sc_hd__nand2_2 _35022_ (.A(_07890_),
    .B(_08085_),
    .Y(_12981_));
 sky130_fd_sc_hd__nand2_2 _35023_ (.A(_12980_),
    .B(_12981_),
    .Y(_12982_));
 sky130_fd_sc_hd__nor2_2 _35024_ (.A(_09677_),
    .B(_12978_),
    .Y(_12983_));
 sky130_fd_sc_hd__inv_2 _35025_ (.A(_12981_),
    .Y(_12984_));
 sky130_fd_sc_hd__nand3b_2 _35026_ (.A_N(_12983_),
    .B(_12979_),
    .C(_12984_),
    .Y(_12985_));
 sky130_fd_sc_hd__nand3_2 _35027_ (.A(_12977_),
    .B(_12982_),
    .C(_12985_),
    .Y(_12986_));
 sky130_fd_sc_hd__nand2_2 _35028_ (.A(_12980_),
    .B(_12984_),
    .Y(_12987_));
 sky130_fd_sc_hd__nand3b_2 _35029_ (.A_N(_12983_),
    .B(_12979_),
    .C(_12981_),
    .Y(_12988_));
 sky130_fd_sc_hd__a21oi_2 _35030_ (.A1(_12593_),
    .A2(_12594_),
    .B1(_12592_),
    .Y(_12989_));
 sky130_fd_sc_hd__nand3_2 _35031_ (.A(_12987_),
    .B(_12988_),
    .C(_12989_),
    .Y(_12990_));
 sky130_fd_sc_hd__a21o_2 _35032_ (.A1(_12653_),
    .A2(_12652_),
    .B1(_12646_),
    .X(_12991_));
 sky130_fd_sc_hd__a21o_2 _35033_ (.A1(_12986_),
    .A2(_12990_),
    .B1(_12991_),
    .X(_12992_));
 sky130_fd_sc_hd__nand3_2 _35034_ (.A(_12986_),
    .B(_12990_),
    .C(_12991_),
    .Y(_12993_));
 sky130_fd_sc_hd__a22oi_2 _35035_ (.A1(_12659_),
    .A2(_12976_),
    .B1(_12992_),
    .B2(_12993_),
    .Y(_12994_));
 sky130_fd_sc_hd__nand2_2 _35036_ (.A(_12976_),
    .B(_12659_),
    .Y(_12995_));
 sky130_fd_sc_hd__nand2_2 _35037_ (.A(_12992_),
    .B(_12993_),
    .Y(_12996_));
 sky130_fd_sc_hd__nor2_2 _35038_ (.A(_12995_),
    .B(_12996_),
    .Y(_12997_));
 sky130_fd_sc_hd__o22ai_2 _35039_ (.A1(_12974_),
    .A2(_12975_),
    .B1(_12994_),
    .B2(_12997_),
    .Y(_12998_));
 sky130_fd_sc_hd__nand2_2 _35040_ (.A(_12620_),
    .B(_12621_),
    .Y(_12999_));
 sky130_fd_sc_hd__nand2_2 _35041_ (.A(_12999_),
    .B(_12616_),
    .Y(_13000_));
 sky130_fd_sc_hd__nor2_2 _35042_ (.A(_12975_),
    .B(_12974_),
    .Y(_13001_));
 sky130_fd_sc_hd__nand2_2 _35043_ (.A(_12996_),
    .B(_12995_),
    .Y(_13002_));
 sky130_fd_sc_hd__nand3b_2 _35044_ (.A_N(_12995_),
    .B(_12992_),
    .C(_12993_),
    .Y(_13003_));
 sky130_fd_sc_hd__nand3_2 _35045_ (.A(_13001_),
    .B(_13002_),
    .C(_13003_),
    .Y(_13004_));
 sky130_fd_sc_hd__nand3_2 _35046_ (.A(_12998_),
    .B(_13000_),
    .C(_13004_),
    .Y(_13005_));
 sky130_fd_sc_hd__a21o_2 _35047_ (.A1(_12972_),
    .A2(_12961_),
    .B1(_12971_),
    .X(_13006_));
 sky130_fd_sc_hd__o21ai_2 _35048_ (.A1(_12962_),
    .A2(_12973_),
    .B1(_13006_),
    .Y(_13007_));
 sky130_fd_sc_hd__o21bai_2 _35049_ (.A1(_12994_),
    .A2(_12997_),
    .B1_N(_13007_),
    .Y(_13008_));
 sky130_fd_sc_hd__a21boi_2 _35050_ (.A1(_12620_),
    .A2(_12621_),
    .B1_N(_12616_),
    .Y(_13009_));
 sky130_fd_sc_hd__nand3_2 _35051_ (.A(_13002_),
    .B(_13003_),
    .C(_13007_),
    .Y(_13010_));
 sky130_fd_sc_hd__o21a_2 _35052_ (.A1(_12665_),
    .A2(_12695_),
    .B1(_12700_),
    .X(_13011_));
 sky130_fd_sc_hd__a31oi_2 _35053_ (.A1(_13008_),
    .A2(_13009_),
    .A3(_13010_),
    .B1(_13011_),
    .Y(_13012_));
 sky130_fd_sc_hd__nand3_2 _35054_ (.A(_13008_),
    .B(_13009_),
    .C(_13010_),
    .Y(_13013_));
 sky130_fd_sc_hd__inv_2 _35055_ (.A(_13011_),
    .Y(_13014_));
 sky130_fd_sc_hd__a21oi_2 _35056_ (.A1(_13013_),
    .A2(_13005_),
    .B1(_13014_),
    .Y(_13015_));
 sky130_fd_sc_hd__a21oi_2 _35057_ (.A1(_13005_),
    .A2(_13012_),
    .B1(_13015_),
    .Y(_13016_));
 sky130_fd_sc_hd__nand2_2 _35058_ (.A(_12951_),
    .B(_13016_),
    .Y(_13017_));
 sky130_fd_sc_hd__a21oi_2 _35059_ (.A1(_12640_),
    .A2(_12642_),
    .B1(_12641_),
    .Y(_13018_));
 sky130_fd_sc_hd__a21oi_2 _35060_ (.A1(_12643_),
    .A2(_12721_),
    .B1(_13018_),
    .Y(_13019_));
 sky130_fd_sc_hd__a21o_2 _35061_ (.A1(_13013_),
    .A2(_13005_),
    .B1(_13014_),
    .X(_13020_));
 sky130_fd_sc_hd__nand2_2 _35062_ (.A(_13012_),
    .B(_13005_),
    .Y(_13021_));
 sky130_fd_sc_hd__nand2_2 _35063_ (.A(_13020_),
    .B(_13021_),
    .Y(_13022_));
 sky130_fd_sc_hd__nand3_2 _35064_ (.A(_13022_),
    .B(_12942_),
    .C(_12950_),
    .Y(_13023_));
 sky130_fd_sc_hd__nand3_2 _35065_ (.A(_13017_),
    .B(_13019_),
    .C(_13023_),
    .Y(_13024_));
 sky130_fd_sc_hd__nand2_2 _35066_ (.A(_12643_),
    .B(_12721_),
    .Y(_13025_));
 sky130_fd_sc_hd__nand2_2 _35067_ (.A(_13025_),
    .B(_12639_),
    .Y(_13026_));
 sky130_fd_sc_hd__and3_2 _35068_ (.A(_13014_),
    .B(_13013_),
    .C(_13005_),
    .X(_13027_));
 sky130_fd_sc_hd__o2bb2ai_2 _35069_ (.A1_N(_12950_),
    .A2_N(_12942_),
    .B1(_13027_),
    .B2(_13015_),
    .Y(_13028_));
 sky130_fd_sc_hd__nand3_2 _35070_ (.A(_13016_),
    .B(_12942_),
    .C(_12950_),
    .Y(_13029_));
 sky130_fd_sc_hd__nand3_2 _35071_ (.A(_13026_),
    .B(_13028_),
    .C(_13029_),
    .Y(_13030_));
 sky130_fd_sc_hd__nand2_2 _35072_ (.A(_13024_),
    .B(_13030_),
    .Y(_13031_));
 sky130_fd_sc_hd__a21o_2 _35073_ (.A1(_11030_),
    .A2(_12729_),
    .B1(_12735_),
    .X(_13032_));
 sky130_fd_sc_hd__nand2_2 _35074_ (.A(_12729_),
    .B(_11029_),
    .Y(_13033_));
 sky130_fd_sc_hd__nor2_2 _35075_ (.A(_13033_),
    .B(_11918_),
    .Y(_13034_));
 sky130_fd_sc_hd__inv_2 _35076_ (.A(_13034_),
    .Y(_13035_));
 sky130_fd_sc_hd__nand2_2 _35077_ (.A(_13032_),
    .B(_13035_),
    .Y(_13036_));
 sky130_fd_sc_hd__nor2_2 _35078_ (.A(_12456_),
    .B(_13036_),
    .Y(_13037_));
 sky130_fd_sc_hd__nand2_2 _35079_ (.A(_13036_),
    .B(_12456_),
    .Y(_13038_));
 sky130_fd_sc_hd__inv_2 _35080_ (.A(_13038_),
    .Y(_13039_));
 sky130_fd_sc_hd__nand3_2 _35081_ (.A(_12679_),
    .B(_12688_),
    .C(_12690_),
    .Y(_13040_));
 sky130_fd_sc_hd__nand2_2 _35082_ (.A(_05851_),
    .B(_19544_),
    .Y(_13041_));
 sky130_fd_sc_hd__nand2_2 _35083_ (.A(_09247_),
    .B(_19540_),
    .Y(_13042_));
 sky130_fd_sc_hd__nor2_2 _35084_ (.A(_13041_),
    .B(_13042_),
    .Y(_13043_));
 sky130_fd_sc_hd__and2_2 _35085_ (.A(_13041_),
    .B(_13042_),
    .X(_13044_));
 sky130_fd_sc_hd__nand2_2 _35086_ (.A(\pcpi_mul.rs1[32] ),
    .B(\pcpi_mul.rs2[6] ),
    .Y(_13045_));
 sky130_fd_sc_hd__buf_1 _35087_ (.A(_13045_),
    .X(_13046_));
 sky130_fd_sc_hd__o21ai_2 _35088_ (.A1(_13043_),
    .A2(_13044_),
    .B1(_13046_),
    .Y(_13047_));
 sky130_fd_sc_hd__a31o_2 _35089_ (.A1(_12685_),
    .A2(_19377_),
    .A3(_19554_),
    .B1(_12684_),
    .X(_13048_));
 sky130_fd_sc_hd__nand2_2 _35090_ (.A(_13041_),
    .B(_13042_),
    .Y(_13049_));
 sky130_fd_sc_hd__inv_2 _35091_ (.A(_13045_),
    .Y(_13050_));
 sky130_fd_sc_hd__buf_1 _35092_ (.A(_13050_),
    .X(_13051_));
 sky130_fd_sc_hd__nand3b_2 _35093_ (.A_N(_13043_),
    .B(_13049_),
    .C(_13051_),
    .Y(_13052_));
 sky130_fd_sc_hd__nand3_2 _35094_ (.A(_13047_),
    .B(_13048_),
    .C(_13052_),
    .Y(_13053_));
 sky130_fd_sc_hd__o21ai_2 _35095_ (.A1(_13043_),
    .A2(_13044_),
    .B1(_13051_),
    .Y(_13054_));
 sky130_fd_sc_hd__nand3b_2 _35096_ (.A_N(_13043_),
    .B(_13049_),
    .C(_13046_),
    .Y(_13055_));
 sky130_fd_sc_hd__a21oi_2 _35097_ (.A1(_12687_),
    .A2(_12685_),
    .B1(_12684_),
    .Y(_13056_));
 sky130_fd_sc_hd__nand3_2 _35098_ (.A(_13054_),
    .B(_13055_),
    .C(_13056_),
    .Y(_13057_));
 sky130_fd_sc_hd__a21o_2 _35099_ (.A1(_12749_),
    .A2(_12750_),
    .B1(_12742_),
    .X(_13058_));
 sky130_fd_sc_hd__a21o_2 _35100_ (.A1(_13053_),
    .A2(_13057_),
    .B1(_13058_),
    .X(_13059_));
 sky130_fd_sc_hd__nand3_2 _35101_ (.A(_13053_),
    .B(_13057_),
    .C(_13058_),
    .Y(_13060_));
 sky130_fd_sc_hd__a22oi_2 _35102_ (.A1(_13040_),
    .A2(_12692_),
    .B1(_13059_),
    .B2(_13060_),
    .Y(_13061_));
 sky130_fd_sc_hd__a21oi_2 _35103_ (.A1(_13053_),
    .A2(_13057_),
    .B1(_13058_),
    .Y(_13062_));
 sky130_fd_sc_hd__nand3_2 _35104_ (.A(_13040_),
    .B(_13060_),
    .C(_12692_),
    .Y(_13063_));
 sky130_fd_sc_hd__nor2_2 _35105_ (.A(_13062_),
    .B(_13063_),
    .Y(_13064_));
 sky130_fd_sc_hd__and2_2 _35106_ (.A(_12760_),
    .B(_12752_),
    .X(_13065_));
 sky130_fd_sc_hd__o21ai_2 _35107_ (.A1(_13061_),
    .A2(_13064_),
    .B1(_13065_),
    .Y(_13066_));
 sky130_fd_sc_hd__nand2_2 _35108_ (.A(_13059_),
    .B(_13060_),
    .Y(_13067_));
 sky130_fd_sc_hd__nand2_2 _35109_ (.A(_13040_),
    .B(_12692_),
    .Y(_13068_));
 sky130_fd_sc_hd__nand2_2 _35110_ (.A(_13067_),
    .B(_13068_),
    .Y(_13069_));
 sky130_fd_sc_hd__nand2_2 _35111_ (.A(_13057_),
    .B(_13058_),
    .Y(_13070_));
 sky130_fd_sc_hd__inv_2 _35112_ (.A(_13053_),
    .Y(_13071_));
 sky130_fd_sc_hd__o2111ai_2 _35113_ (.A1(_13070_),
    .A2(_13071_),
    .B1(_12692_),
    .C1(_13040_),
    .D1(_13059_),
    .Y(_13072_));
 sky130_fd_sc_hd__nand3b_2 _35114_ (.A_N(_13065_),
    .B(_13069_),
    .C(_13072_),
    .Y(_13073_));
 sky130_fd_sc_hd__o21ai_2 _35115_ (.A1(_12765_),
    .A2(_12762_),
    .B1(_12770_),
    .Y(_13074_));
 sky130_fd_sc_hd__a21oi_2 _35116_ (.A1(_13066_),
    .A2(_13073_),
    .B1(_13074_),
    .Y(_13075_));
 sky130_fd_sc_hd__a21oi_2 _35117_ (.A1(_12767_),
    .A2(_12768_),
    .B1(_12765_),
    .Y(_13076_));
 sky130_fd_sc_hd__o211a_2 _35118_ (.A1(_12763_),
    .A2(_13076_),
    .B1(_13073_),
    .C1(_13066_),
    .X(_13077_));
 sky130_fd_sc_hd__o22ai_2 _35119_ (.A1(_13037_),
    .A2(_13039_),
    .B1(_13075_),
    .B2(_13077_),
    .Y(_13078_));
 sky130_fd_sc_hd__nand2_2 _35120_ (.A(_12708_),
    .B(_12709_),
    .Y(_13079_));
 sky130_fd_sc_hd__nand2_2 _35121_ (.A(_13079_),
    .B(_12702_),
    .Y(_13080_));
 sky130_fd_sc_hd__a21o_2 _35122_ (.A1(_13066_),
    .A2(_13073_),
    .B1(_13074_),
    .X(_13081_));
 sky130_fd_sc_hd__nor2_2 _35123_ (.A(_13037_),
    .B(_13039_),
    .Y(_13082_));
 sky130_fd_sc_hd__nand3_2 _35124_ (.A(_13074_),
    .B(_13066_),
    .C(_13073_),
    .Y(_13083_));
 sky130_fd_sc_hd__nand3_2 _35125_ (.A(_13081_),
    .B(_13082_),
    .C(_13083_),
    .Y(_13084_));
 sky130_fd_sc_hd__nand3_2 _35126_ (.A(_13078_),
    .B(_13080_),
    .C(_13084_),
    .Y(_13085_));
 sky130_fd_sc_hd__o21ai_2 _35127_ (.A1(_13075_),
    .A2(_13077_),
    .B1(_13082_),
    .Y(_13086_));
 sky130_fd_sc_hd__a21boi_2 _35128_ (.A1(_12709_),
    .A2(_12708_),
    .B1_N(_12702_),
    .Y(_13087_));
 sky130_fd_sc_hd__or2b_2 _35129_ (.A(_13037_),
    .B_N(_13038_),
    .X(_13088_));
 sky130_fd_sc_hd__nand3_2 _35130_ (.A(_13081_),
    .B(_13083_),
    .C(_13088_),
    .Y(_13089_));
 sky130_fd_sc_hd__a32oi_2 _35131_ (.A1(_13086_),
    .A2(_13087_),
    .A3(_13089_),
    .B1(_12777_),
    .B2(_12781_),
    .Y(_13090_));
 sky130_fd_sc_hd__nand3_2 _35132_ (.A(_13086_),
    .B(_13087_),
    .C(_13089_),
    .Y(_13091_));
 sky130_fd_sc_hd__nand2_2 _35133_ (.A(_12781_),
    .B(_12777_),
    .Y(_13092_));
 sky130_fd_sc_hd__a21oi_2 _35134_ (.A1(_13091_),
    .A2(_13085_),
    .B1(_13092_),
    .Y(_13093_));
 sky130_fd_sc_hd__a21oi_2 _35135_ (.A1(_13085_),
    .A2(_13090_),
    .B1(_13093_),
    .Y(_13094_));
 sky130_fd_sc_hd__nand2_2 _35136_ (.A(_13031_),
    .B(_13094_),
    .Y(_13095_));
 sky130_fd_sc_hd__a21o_2 _35137_ (.A1(_13091_),
    .A2(_13085_),
    .B1(_13092_),
    .X(_13096_));
 sky130_fd_sc_hd__nand3_2 _35138_ (.A(_13091_),
    .B(_13085_),
    .C(_13092_),
    .Y(_13097_));
 sky130_fd_sc_hd__nand2_2 _35139_ (.A(_13096_),
    .B(_13097_),
    .Y(_13098_));
 sky130_fd_sc_hd__nand3_2 _35140_ (.A(_13098_),
    .B(_13024_),
    .C(_13030_),
    .Y(_13099_));
 sky130_fd_sc_hd__nor2_2 _35141_ (.A(_12794_),
    .B(_12785_),
    .Y(_13100_));
 sky130_fd_sc_hd__nand2_2 _35142_ (.A(_12738_),
    .B(_12457_),
    .Y(_13101_));
 sky130_fd_sc_hd__nand2_2 _35143_ (.A(_13101_),
    .B(_12736_),
    .Y(_13102_));
 sky130_fd_sc_hd__inv_2 _35144_ (.A(_13102_),
    .Y(_13103_));
 sky130_fd_sc_hd__nand2_2 _35145_ (.A(_13100_),
    .B(_13103_),
    .Y(_13104_));
 sky130_fd_sc_hd__o21ai_2 _35146_ (.A1(_12794_),
    .A2(_12785_),
    .B1(_13102_),
    .Y(_13105_));
 sky130_fd_sc_hd__nand2_2 _35147_ (.A(_13104_),
    .B(_13105_),
    .Y(_13106_));
 sky130_fd_sc_hd__a31oi_2 _35148_ (.A1(_12841_),
    .A2(_13095_),
    .A3(_13099_),
    .B1(_13106_),
    .Y(_13107_));
 sky130_fd_sc_hd__nand3_2 _35149_ (.A(_12715_),
    .B(_12795_),
    .C(_12796_),
    .Y(_13108_));
 sky130_fd_sc_hd__nand2_2 _35150_ (.A(_13108_),
    .B(_12723_),
    .Y(_13109_));
 sky130_fd_sc_hd__nand2_2 _35151_ (.A(_13031_),
    .B(_13098_),
    .Y(_13110_));
 sky130_fd_sc_hd__nand3_2 _35152_ (.A(_13094_),
    .B(_13024_),
    .C(_13030_),
    .Y(_13111_));
 sky130_fd_sc_hd__nand3_2 _35153_ (.A(_13109_),
    .B(_13110_),
    .C(_13111_),
    .Y(_13112_));
 sky130_fd_sc_hd__nand2_2 _35154_ (.A(_13107_),
    .B(_13112_),
    .Y(_13113_));
 sky130_fd_sc_hd__nand3_2 _35155_ (.A(_12841_),
    .B(_13095_),
    .C(_13099_),
    .Y(_13114_));
 sky130_fd_sc_hd__nand2_2 _35156_ (.A(_13114_),
    .B(_13112_),
    .Y(_13115_));
 sky130_fd_sc_hd__nand2_2 _35157_ (.A(_13115_),
    .B(_13106_),
    .Y(_13116_));
 sky130_fd_sc_hd__o211ai_2 _35158_ (.A1(_12838_),
    .A2(_12839_),
    .B1(_13113_),
    .C1(_13116_),
    .Y(_13117_));
 sky130_fd_sc_hd__and3_2 _35159_ (.A(_12803_),
    .B(_12786_),
    .C(_13103_),
    .X(_13118_));
 sky130_fd_sc_hd__nor2_2 _35160_ (.A(_13103_),
    .B(_13100_),
    .Y(_13119_));
 sky130_fd_sc_hd__nor2_2 _35161_ (.A(_13118_),
    .B(_13119_),
    .Y(_13120_));
 sky130_fd_sc_hd__nand2_2 _35162_ (.A(_13115_),
    .B(_13120_),
    .Y(_13121_));
 sky130_fd_sc_hd__a21oi_2 _35163_ (.A1(_12799_),
    .A2(_12814_),
    .B1(_12838_),
    .Y(_13122_));
 sky130_fd_sc_hd__nand3_2 _35164_ (.A(_13114_),
    .B(_13112_),
    .C(_13106_),
    .Y(_13123_));
 sky130_fd_sc_hd__nand3_2 _35165_ (.A(_13121_),
    .B(_13122_),
    .C(_13123_),
    .Y(_13124_));
 sky130_fd_sc_hd__inv_2 _35166_ (.A(_12810_),
    .Y(_13125_));
 sky130_fd_sc_hd__nand3_2 _35167_ (.A(_13117_),
    .B(_13124_),
    .C(_13125_),
    .Y(_13126_));
 sky130_fd_sc_hd__o2bb2ai_2 _35168_ (.A1_N(_13117_),
    .A2_N(_13124_),
    .B1(_12820_),
    .B2(_12811_),
    .Y(_13127_));
 sky130_fd_sc_hd__o211ai_2 _35169_ (.A1(_12836_),
    .A2(_12837_),
    .B1(_13126_),
    .C1(_13127_),
    .Y(_13128_));
 sky130_fd_sc_hd__nand2_2 _35170_ (.A(_13117_),
    .B(_13124_),
    .Y(_13129_));
 sky130_fd_sc_hd__nand2_2 _35171_ (.A(_13129_),
    .B(_13125_),
    .Y(_13130_));
 sky130_fd_sc_hd__a21oi_2 _35172_ (.A1(_12825_),
    .A2(_12194_),
    .B1(_12836_),
    .Y(_13131_));
 sky130_fd_sc_hd__nand3_2 _35173_ (.A(_13117_),
    .B(_13124_),
    .C(_12810_),
    .Y(_13132_));
 sky130_fd_sc_hd__nand3_2 _35174_ (.A(_13130_),
    .B(_13131_),
    .C(_13132_),
    .Y(_13133_));
 sky130_fd_sc_hd__and2_2 _35175_ (.A(_13128_),
    .B(_13133_),
    .X(_13134_));
 sky130_fd_sc_hd__nand2_2 _35176_ (.A(_12832_),
    .B(_12511_),
    .Y(_13135_));
 sky130_fd_sc_hd__nand2_2 _35177_ (.A(_13135_),
    .B(_12829_),
    .Y(_13136_));
 sky130_fd_sc_hd__inv_2 _35178_ (.A(_13136_),
    .Y(_13137_));
 sky130_fd_sc_hd__nand2_2 _35179_ (.A(_12833_),
    .B(_12513_),
    .Y(_13138_));
 sky130_fd_sc_hd__nor2_2 _35180_ (.A(_13138_),
    .B(_12518_),
    .Y(_13139_));
 sky130_fd_sc_hd__nor3_2 _35181_ (.A(_13134_),
    .B(_13137_),
    .C(_13139_),
    .Y(_13140_));
 sky130_fd_sc_hd__o21a_2 _35182_ (.A1(_13137_),
    .A2(_13139_),
    .B1(_13134_),
    .X(_13141_));
 sky130_fd_sc_hd__nor2_2 _35183_ (.A(_13140_),
    .B(_13141_),
    .Y(_02657_));
 sky130_fd_sc_hd__o211ai_2 _35184_ (.A1(_13138_),
    .A2(_12518_),
    .B1(_13128_),
    .C1(_13136_),
    .Y(_13142_));
 sky130_fd_sc_hd__nand2_2 _35185_ (.A(_12847_),
    .B(_12850_),
    .Y(_13143_));
 sky130_fd_sc_hd__nand3_2 _35186_ (.A(_10824_),
    .B(_10823_),
    .C(_06052_),
    .Y(_13144_));
 sky130_fd_sc_hd__nor2_2 _35187_ (.A(_19620_),
    .B(_13144_),
    .Y(_13145_));
 sky130_fd_sc_hd__buf_1 _35188_ (.A(_10822_),
    .X(_13146_));
 sky130_fd_sc_hd__nand2_2 _35189_ (.A(_13146_),
    .B(_05613_),
    .Y(_13147_));
 sky130_fd_sc_hd__o21a_2 _35190_ (.A1(_19620_),
    .A2(_18182_),
    .B1(_13147_),
    .X(_13148_));
 sky130_fd_sc_hd__nand2_2 _35191_ (.A(_19311_),
    .B(_05734_),
    .Y(_13149_));
 sky130_fd_sc_hd__o21ai_2 _35192_ (.A1(_13145_),
    .A2(_13148_),
    .B1(_13149_),
    .Y(_13150_));
 sky130_fd_sc_hd__nand3b_2 _35193_ (.A_N(_13147_),
    .B(_11122_),
    .C(_06333_),
    .Y(_13151_));
 sky130_fd_sc_hd__o21ai_2 _35194_ (.A1(_05421_),
    .A2(_10830_),
    .B1(_13147_),
    .Y(_13152_));
 sky130_fd_sc_hd__inv_2 _35195_ (.A(_13149_),
    .Y(_13153_));
 sky130_fd_sc_hd__nand3_2 _35196_ (.A(_13151_),
    .B(_13152_),
    .C(_13153_),
    .Y(_13154_));
 sky130_fd_sc_hd__a22oi_2 _35197_ (.A1(_12848_),
    .A2(_13143_),
    .B1(_13150_),
    .B2(_13154_),
    .Y(_13155_));
 sky130_fd_sc_hd__o211a_2 _35198_ (.A1(_19620_),
    .A2(_13144_),
    .B1(_13153_),
    .C1(_13152_),
    .X(_13156_));
 sky130_fd_sc_hd__a21oi_2 _35199_ (.A1(_13151_),
    .A2(_13152_),
    .B1(_13153_),
    .Y(_13157_));
 sky130_fd_sc_hd__nand2_2 _35200_ (.A(_13143_),
    .B(_12848_),
    .Y(_13158_));
 sky130_fd_sc_hd__nor3_2 _35201_ (.A(_13156_),
    .B(_13157_),
    .C(_13158_),
    .Y(_13159_));
 sky130_fd_sc_hd__nand2_2 _35202_ (.A(_10138_),
    .B(_05733_),
    .Y(_13160_));
 sky130_fd_sc_hd__nand2_2 _35203_ (.A(_09602_),
    .B(_06369_),
    .Y(_13161_));
 sky130_fd_sc_hd__nor2_2 _35204_ (.A(_13160_),
    .B(_13161_),
    .Y(_13162_));
 sky130_fd_sc_hd__nand2_2 _35205_ (.A(_13160_),
    .B(_13161_),
    .Y(_13163_));
 sky130_fd_sc_hd__inv_2 _35206_ (.A(_13163_),
    .Y(_13164_));
 sky130_fd_sc_hd__nor2_2 _35207_ (.A(_09357_),
    .B(_06391_),
    .Y(_13165_));
 sky130_fd_sc_hd__o21ai_2 _35208_ (.A1(_13162_),
    .A2(_13164_),
    .B1(_13165_),
    .Y(_13166_));
 sky130_fd_sc_hd__inv_2 _35209_ (.A(_13165_),
    .Y(_13167_));
 sky130_fd_sc_hd__or2_2 _35210_ (.A(_13160_),
    .B(_13161_),
    .X(_13168_));
 sky130_fd_sc_hd__nand3_2 _35211_ (.A(_13167_),
    .B(_13163_),
    .C(_13168_),
    .Y(_13169_));
 sky130_fd_sc_hd__nand2_2 _35212_ (.A(_13166_),
    .B(_13169_),
    .Y(_13170_));
 sky130_fd_sc_hd__o21ai_2 _35213_ (.A1(_13155_),
    .A2(_13159_),
    .B1(_13170_),
    .Y(_13171_));
 sky130_fd_sc_hd__a21boi_2 _35214_ (.A1(_12857_),
    .A2(_12865_),
    .B1_N(_12854_),
    .Y(_13172_));
 sky130_fd_sc_hd__nand3b_2 _35215_ (.A_N(_13158_),
    .B(_13150_),
    .C(_13154_),
    .Y(_13173_));
 sky130_fd_sc_hd__o21ai_2 _35216_ (.A1(_13156_),
    .A2(_13157_),
    .B1(_13158_),
    .Y(_13174_));
 sky130_fd_sc_hd__nand2_2 _35217_ (.A(_13168_),
    .B(_13165_),
    .Y(_13175_));
 sky130_fd_sc_hd__o21ai_2 _35218_ (.A1(_13162_),
    .A2(_13164_),
    .B1(_13167_),
    .Y(_13176_));
 sky130_fd_sc_hd__o21ai_2 _35219_ (.A1(_13164_),
    .A2(_13175_),
    .B1(_13176_),
    .Y(_13177_));
 sky130_fd_sc_hd__nand3_2 _35220_ (.A(_13173_),
    .B(_13174_),
    .C(_13177_),
    .Y(_13178_));
 sky130_fd_sc_hd__nand3_2 _35221_ (.A(_13171_),
    .B(_13172_),
    .C(_13178_),
    .Y(_13179_));
 sky130_fd_sc_hd__o21ai_2 _35222_ (.A1(_13155_),
    .A2(_13159_),
    .B1(_13177_),
    .Y(_13180_));
 sky130_fd_sc_hd__nand2_2 _35223_ (.A(_12865_),
    .B(_12857_),
    .Y(_13181_));
 sky130_fd_sc_hd__nand2_2 _35224_ (.A(_13181_),
    .B(_12854_),
    .Y(_13182_));
 sky130_fd_sc_hd__nand3_2 _35225_ (.A(_13173_),
    .B(_13174_),
    .C(_13170_),
    .Y(_13183_));
 sky130_fd_sc_hd__nand3_2 _35226_ (.A(_13180_),
    .B(_13182_),
    .C(_13183_),
    .Y(_13184_));
 sky130_fd_sc_hd__nand2_2 _35227_ (.A(_19327_),
    .B(_07311_),
    .Y(_13185_));
 sky130_fd_sc_hd__nand2_2 _35228_ (.A(_10158_),
    .B(_08761_),
    .Y(_13186_));
 sky130_fd_sc_hd__nor2_2 _35229_ (.A(_13185_),
    .B(_13186_),
    .Y(_13187_));
 sky130_fd_sc_hd__and2_2 _35230_ (.A(_13185_),
    .B(_13186_),
    .X(_13188_));
 sky130_fd_sc_hd__nand2_2 _35231_ (.A(_10862_),
    .B(_19594_),
    .Y(_13189_));
 sky130_fd_sc_hd__o21ai_2 _35232_ (.A1(_13187_),
    .A2(_13188_),
    .B1(_13189_),
    .Y(_13190_));
 sky130_fd_sc_hd__a21o_2 _35233_ (.A1(_12859_),
    .A2(_12861_),
    .B1(_12858_),
    .X(_13191_));
 sky130_fd_sc_hd__nand2_2 _35234_ (.A(_13185_),
    .B(_13186_),
    .Y(_13192_));
 sky130_fd_sc_hd__inv_2 _35235_ (.A(_13189_),
    .Y(_13193_));
 sky130_fd_sc_hd__nand3b_2 _35236_ (.A_N(_13187_),
    .B(_13192_),
    .C(_13193_),
    .Y(_13194_));
 sky130_fd_sc_hd__nand3_2 _35237_ (.A(_13190_),
    .B(_13191_),
    .C(_13194_),
    .Y(_13195_));
 sky130_fd_sc_hd__o21ai_2 _35238_ (.A1(_13187_),
    .A2(_13188_),
    .B1(_13193_),
    .Y(_13196_));
 sky130_fd_sc_hd__nand3b_2 _35239_ (.A_N(_13187_),
    .B(_13192_),
    .C(_13189_),
    .Y(_13197_));
 sky130_fd_sc_hd__a21oi_2 _35240_ (.A1(_12859_),
    .A2(_12861_),
    .B1(_12858_),
    .Y(_13198_));
 sky130_fd_sc_hd__nand3_2 _35241_ (.A(_13196_),
    .B(_13197_),
    .C(_13198_),
    .Y(_13199_));
 sky130_fd_sc_hd__a21oi_2 _35242_ (.A1(_12883_),
    .A2(_12882_),
    .B1(_12878_),
    .Y(_13200_));
 sky130_fd_sc_hd__inv_2 _35243_ (.A(_13200_),
    .Y(_13201_));
 sky130_fd_sc_hd__a21oi_2 _35244_ (.A1(_13195_),
    .A2(_13199_),
    .B1(_13201_),
    .Y(_13202_));
 sky130_fd_sc_hd__nand2_2 _35245_ (.A(_13195_),
    .B(_13199_),
    .Y(_13203_));
 sky130_fd_sc_hd__nor2_2 _35246_ (.A(_13200_),
    .B(_13203_),
    .Y(_13204_));
 sky130_fd_sc_hd__o2bb2ai_2 _35247_ (.A1_N(_13179_),
    .A2_N(_13184_),
    .B1(_13202_),
    .B2(_13204_),
    .Y(_13205_));
 sky130_fd_sc_hd__nor2_2 _35248_ (.A(_13202_),
    .B(_13204_),
    .Y(_13206_));
 sky130_fd_sc_hd__nand3_2 _35249_ (.A(_13184_),
    .B(_13179_),
    .C(_13206_),
    .Y(_13207_));
 sky130_fd_sc_hd__nand2_2 _35250_ (.A(_12873_),
    .B(_12893_),
    .Y(_13208_));
 sky130_fd_sc_hd__nand2_2 _35251_ (.A(_13208_),
    .B(_12868_),
    .Y(_13209_));
 sky130_fd_sc_hd__a21oi_2 _35252_ (.A1(_13205_),
    .A2(_13207_),
    .B1(_13209_),
    .Y(_13210_));
 sky130_fd_sc_hd__and3_2 _35253_ (.A(_13180_),
    .B(_13182_),
    .C(_13183_),
    .X(_13211_));
 sky130_fd_sc_hd__nand2_2 _35254_ (.A(_13179_),
    .B(_13206_),
    .Y(_13212_));
 sky130_fd_sc_hd__o211a_2 _35255_ (.A1(_13211_),
    .A2(_13212_),
    .B1(_13205_),
    .C1(_13209_),
    .X(_13213_));
 sky130_fd_sc_hd__a21oi_2 _35256_ (.A1(_12914_),
    .A2(_12916_),
    .B1(_12911_),
    .Y(_13214_));
 sky130_fd_sc_hd__nand2_2 _35257_ (.A(_08391_),
    .B(_06542_),
    .Y(_13215_));
 sky130_fd_sc_hd__nand2_2 _35258_ (.A(_08386_),
    .B(_06951_),
    .Y(_13216_));
 sky130_fd_sc_hd__nor2_2 _35259_ (.A(_13215_),
    .B(_13216_),
    .Y(_13217_));
 sky130_fd_sc_hd__and2_2 _35260_ (.A(_13215_),
    .B(_13216_),
    .X(_13218_));
 sky130_fd_sc_hd__nand2_2 _35261_ (.A(_07976_),
    .B(_19585_),
    .Y(_13219_));
 sky130_fd_sc_hd__o21ai_2 _35262_ (.A1(_13217_),
    .A2(_13218_),
    .B1(_13219_),
    .Y(_13220_));
 sky130_fd_sc_hd__inv_2 _35263_ (.A(_13219_),
    .Y(_13221_));
 sky130_fd_sc_hd__nand2_2 _35264_ (.A(_13215_),
    .B(_13216_),
    .Y(_13222_));
 sky130_fd_sc_hd__nand3b_2 _35265_ (.A_N(_13217_),
    .B(_13221_),
    .C(_13222_),
    .Y(_13223_));
 sky130_fd_sc_hd__nand3b_2 _35266_ (.A_N(_13214_),
    .B(_13220_),
    .C(_13223_),
    .Y(_13224_));
 sky130_fd_sc_hd__o21ai_2 _35267_ (.A1(_13217_),
    .A2(_13218_),
    .B1(_13221_),
    .Y(_13225_));
 sky130_fd_sc_hd__nand3b_2 _35268_ (.A_N(_13217_),
    .B(_13219_),
    .C(_13222_),
    .Y(_13226_));
 sky130_fd_sc_hd__nand3_2 _35269_ (.A(_13225_),
    .B(_13226_),
    .C(_13214_),
    .Y(_13227_));
 sky130_fd_sc_hd__nand2_2 _35270_ (.A(_19347_),
    .B(_07593_),
    .Y(_13228_));
 sky130_fd_sc_hd__nand2_2 _35271_ (.A(_07895_),
    .B(_07358_),
    .Y(_13229_));
 sky130_fd_sc_hd__nor2_2 _35272_ (.A(_13228_),
    .B(_13229_),
    .Y(_13230_));
 sky130_fd_sc_hd__nand2_2 _35273_ (.A(_13228_),
    .B(_13229_),
    .Y(_13231_));
 sky130_fd_sc_hd__inv_2 _35274_ (.A(_13231_),
    .Y(_13232_));
 sky130_fd_sc_hd__nor2_2 _35275_ (.A(_07053_),
    .B(_11660_),
    .Y(_13233_));
 sky130_fd_sc_hd__o21ai_2 _35276_ (.A1(_13230_),
    .A2(_13232_),
    .B1(_13233_),
    .Y(_13234_));
 sky130_fd_sc_hd__or2_2 _35277_ (.A(_13228_),
    .B(_13229_),
    .X(_13235_));
 sky130_fd_sc_hd__nand3b_2 _35278_ (.A_N(_13233_),
    .B(_13235_),
    .C(_13231_),
    .Y(_13236_));
 sky130_fd_sc_hd__nand2_2 _35279_ (.A(_13234_),
    .B(_13236_),
    .Y(_13237_));
 sky130_fd_sc_hd__a21o_2 _35280_ (.A1(_13224_),
    .A2(_13227_),
    .B1(_13237_),
    .X(_13238_));
 sky130_fd_sc_hd__nand3_2 _35281_ (.A(_13224_),
    .B(_13237_),
    .C(_13227_),
    .Y(_13239_));
 sky130_fd_sc_hd__nand2_2 _35282_ (.A(_12889_),
    .B(_12890_),
    .Y(_13240_));
 sky130_fd_sc_hd__nand2_2 _35283_ (.A(_13240_),
    .B(_12885_),
    .Y(_13241_));
 sky130_fd_sc_hd__a21o_2 _35284_ (.A1(_13238_),
    .A2(_13239_),
    .B1(_13241_),
    .X(_13242_));
 sky130_fd_sc_hd__nand3_2 _35285_ (.A(_13238_),
    .B(_13241_),
    .C(_13239_),
    .Y(_13243_));
 sky130_fd_sc_hd__nand2_2 _35286_ (.A(_12926_),
    .B(_12920_),
    .Y(_13244_));
 sky130_fd_sc_hd__nand2_2 _35287_ (.A(_13244_),
    .B(_12924_),
    .Y(_13245_));
 sky130_fd_sc_hd__a21oi_2 _35288_ (.A1(_13242_),
    .A2(_13243_),
    .B1(_13245_),
    .Y(_13246_));
 sky130_fd_sc_hd__and3_2 _35289_ (.A(_13242_),
    .B(_13243_),
    .C(_13245_),
    .X(_13247_));
 sky130_fd_sc_hd__nor2_2 _35290_ (.A(_13246_),
    .B(_13247_),
    .Y(_13248_));
 sky130_fd_sc_hd__o21ai_2 _35291_ (.A1(_13210_),
    .A2(_13213_),
    .B1(_13248_),
    .Y(_13249_));
 sky130_fd_sc_hd__a21boi_2 _35292_ (.A1(_12948_),
    .A2(_12898_),
    .B1_N(_12902_),
    .Y(_13250_));
 sky130_fd_sc_hd__nand2_2 _35293_ (.A(_13205_),
    .B(_13207_),
    .Y(_13251_));
 sky130_fd_sc_hd__and2_2 _35294_ (.A(_13208_),
    .B(_12868_),
    .X(_13252_));
 sky130_fd_sc_hd__nand2_2 _35295_ (.A(_13251_),
    .B(_13252_),
    .Y(_13253_));
 sky130_fd_sc_hd__nand3_2 _35296_ (.A(_13209_),
    .B(_13205_),
    .C(_13207_),
    .Y(_13254_));
 sky130_fd_sc_hd__and3_2 _35297_ (.A(_13238_),
    .B(_13241_),
    .C(_13239_),
    .X(_13255_));
 sky130_fd_sc_hd__nand2_2 _35298_ (.A(_13242_),
    .B(_13245_),
    .Y(_13256_));
 sky130_fd_sc_hd__a21oi_2 _35299_ (.A1(_13238_),
    .A2(_13239_),
    .B1(_13241_),
    .Y(_13257_));
 sky130_fd_sc_hd__inv_2 _35300_ (.A(_13245_),
    .Y(_13258_));
 sky130_fd_sc_hd__o21ai_2 _35301_ (.A1(_13257_),
    .A2(_13255_),
    .B1(_13258_),
    .Y(_13259_));
 sky130_fd_sc_hd__o21ai_2 _35302_ (.A1(_13255_),
    .A2(_13256_),
    .B1(_13259_),
    .Y(_13260_));
 sky130_fd_sc_hd__nand3_2 _35303_ (.A(_13253_),
    .B(_13254_),
    .C(_13260_),
    .Y(_13261_));
 sky130_fd_sc_hd__nand3_2 _35304_ (.A(_13249_),
    .B(_13250_),
    .C(_13261_),
    .Y(_13262_));
 sky130_fd_sc_hd__o22ai_2 _35305_ (.A1(_13247_),
    .A2(_13246_),
    .B1(_13210_),
    .B2(_13213_),
    .Y(_13263_));
 sky130_fd_sc_hd__nand2_2 _35306_ (.A(_12552_),
    .B(_12586_),
    .Y(_13264_));
 sky130_fd_sc_hd__a22oi_2 _35307_ (.A1(_12559_),
    .A2(_13264_),
    .B1(_12901_),
    .B2(_12900_),
    .Y(_13265_));
 sky130_fd_sc_hd__o21ai_2 _35308_ (.A1(_12938_),
    .A2(_13265_),
    .B1(_12902_),
    .Y(_13266_));
 sky130_fd_sc_hd__nand3_2 _35309_ (.A(_13253_),
    .B(_13248_),
    .C(_13254_),
    .Y(_13267_));
 sky130_fd_sc_hd__nand3_2 _35310_ (.A(_13263_),
    .B(_13266_),
    .C(_13267_),
    .Y(_13268_));
 sky130_fd_sc_hd__nand2_2 _35311_ (.A(_13262_),
    .B(_13268_),
    .Y(_13269_));
 sky130_fd_sc_hd__and4_2 _35312_ (.A(_06441_),
    .B(_06272_),
    .C(\pcpi_mul.rs1[26] ),
    .D(_08645_),
    .X(_13270_));
 sky130_fd_sc_hd__nor2_2 _35313_ (.A(_06118_),
    .B(_11374_),
    .Y(_13271_));
 sky130_fd_sc_hd__a22o_2 _35314_ (.A1(_06278_),
    .A2(_19564_),
    .B1(_06276_),
    .B2(_08905_),
    .X(_13272_));
 sky130_fd_sc_hd__nand3b_2 _35315_ (.A_N(_13270_),
    .B(_13271_),
    .C(_13272_),
    .Y(_13273_));
 sky130_fd_sc_hd__buf_1 _35316_ (.A(_11374_),
    .X(_13274_));
 sky130_fd_sc_hd__a22oi_2 _35317_ (.A1(_06790_),
    .A2(_08920_),
    .B1(_06115_),
    .B2(_09220_),
    .Y(_13275_));
 sky130_fd_sc_hd__o22ai_2 _35318_ (.A1(_06119_),
    .A2(_13274_),
    .B1(_13275_),
    .B2(_13270_),
    .Y(_13276_));
 sky130_fd_sc_hd__nand2_2 _35319_ (.A(_13273_),
    .B(_13276_),
    .Y(_13277_));
 sky130_fd_sc_hd__a21oi_2 _35320_ (.A1(_12957_),
    .A2(_12959_),
    .B1(_12955_),
    .Y(_13278_));
 sky130_fd_sc_hd__nand2_2 _35321_ (.A(_13277_),
    .B(_13278_),
    .Y(_13279_));
 sky130_fd_sc_hd__a31o_2 _35322_ (.A1(_12959_),
    .A2(_19368_),
    .A3(_09216_),
    .B1(_12955_),
    .X(_13280_));
 sky130_fd_sc_hd__nand3_2 _35323_ (.A(_13280_),
    .B(_13273_),
    .C(_13276_),
    .Y(_13281_));
 sky130_fd_sc_hd__and4_2 _35324_ (.A(_19370_),
    .B(_05958_),
    .C(_19548_),
    .D(_19552_),
    .X(_13282_));
 sky130_fd_sc_hd__nor2_2 _35325_ (.A(_05496_),
    .B(_10534_),
    .Y(_13283_));
 sky130_fd_sc_hd__a22o_2 _35326_ (.A1(_09051_),
    .A2(_11410_),
    .B1(_05803_),
    .B2(_10538_),
    .X(_13284_));
 sky130_fd_sc_hd__nand3b_2 _35327_ (.A_N(_13282_),
    .B(_13283_),
    .C(_13284_),
    .Y(_13285_));
 sky130_fd_sc_hd__a22oi_2 _35328_ (.A1(_05807_),
    .A2(_09722_),
    .B1(_05808_),
    .B2(_11765_),
    .Y(_13286_));
 sky130_fd_sc_hd__o21bai_2 _35329_ (.A1(_13286_),
    .A2(_13282_),
    .B1_N(_13283_),
    .Y(_13287_));
 sky130_fd_sc_hd__nand2_2 _35330_ (.A(_13285_),
    .B(_13287_),
    .Y(_13288_));
 sky130_fd_sc_hd__inv_2 _35331_ (.A(_13288_),
    .Y(_13289_));
 sky130_fd_sc_hd__a21oi_2 _35332_ (.A1(_13279_),
    .A2(_13281_),
    .B1(_13289_),
    .Y(_13290_));
 sky130_fd_sc_hd__and3_2 _35333_ (.A(_13289_),
    .B(_13279_),
    .C(_13281_),
    .X(_13291_));
 sky130_fd_sc_hd__a22o_2 _35334_ (.A1(_07903_),
    .A2(_08596_),
    .B1(_07895_),
    .B2(_07593_),
    .X(_13292_));
 sky130_fd_sc_hd__a21o_2 _35335_ (.A1(_12903_),
    .A2(_13292_),
    .B1(_12905_),
    .X(_13293_));
 sky130_fd_sc_hd__nand2_2 _35336_ (.A(_06821_),
    .B(_07837_),
    .Y(_13294_));
 sky130_fd_sc_hd__nand2_2 _35337_ (.A(_07417_),
    .B(_08085_),
    .Y(_13295_));
 sky130_fd_sc_hd__nor2_2 _35338_ (.A(_13294_),
    .B(_13295_),
    .Y(_13296_));
 sky130_fd_sc_hd__and2_2 _35339_ (.A(_13294_),
    .B(_13295_),
    .X(_13297_));
 sky130_fd_sc_hd__nand2_2 _35340_ (.A(_19359_),
    .B(_08661_),
    .Y(_13298_));
 sky130_fd_sc_hd__o21ai_2 _35341_ (.A1(_13296_),
    .A2(_13297_),
    .B1(_13298_),
    .Y(_13299_));
 sky130_fd_sc_hd__nand2_2 _35342_ (.A(_13294_),
    .B(_13295_),
    .Y(_13300_));
 sky130_fd_sc_hd__inv_2 _35343_ (.A(_13298_),
    .Y(_13301_));
 sky130_fd_sc_hd__nand3b_2 _35344_ (.A_N(_13296_),
    .B(_13300_),
    .C(_13301_),
    .Y(_13302_));
 sky130_fd_sc_hd__nand3_2 _35345_ (.A(_13293_),
    .B(_13299_),
    .C(_13302_),
    .Y(_13303_));
 sky130_fd_sc_hd__o21ai_2 _35346_ (.A1(_13296_),
    .A2(_13297_),
    .B1(_13301_),
    .Y(_13304_));
 sky130_fd_sc_hd__nand3b_2 _35347_ (.A_N(_13296_),
    .B(_13300_),
    .C(_13298_),
    .Y(_13305_));
 sky130_fd_sc_hd__a21oi_2 _35348_ (.A1(_12903_),
    .A2(_13292_),
    .B1(_12905_),
    .Y(_13306_));
 sky130_fd_sc_hd__nand3_2 _35349_ (.A(_13304_),
    .B(_13305_),
    .C(_13306_),
    .Y(_13307_));
 sky130_fd_sc_hd__nand2_2 _35350_ (.A(_13303_),
    .B(_13307_),
    .Y(_13308_));
 sky130_fd_sc_hd__a21oi_2 _35351_ (.A1(_12979_),
    .A2(_12984_),
    .B1(_12983_),
    .Y(_13309_));
 sky130_fd_sc_hd__nand2_2 _35352_ (.A(_13308_),
    .B(_13309_),
    .Y(_13310_));
 sky130_fd_sc_hd__inv_2 _35353_ (.A(_13309_),
    .Y(_13311_));
 sky130_fd_sc_hd__nand3_2 _35354_ (.A(_13303_),
    .B(_13307_),
    .C(_13311_),
    .Y(_13312_));
 sky130_fd_sc_hd__nand2_2 _35355_ (.A(_12993_),
    .B(_12986_),
    .Y(_13313_));
 sky130_fd_sc_hd__a21oi_2 _35356_ (.A1(_13310_),
    .A2(_13312_),
    .B1(_13313_),
    .Y(_13314_));
 sky130_fd_sc_hd__inv_2 _35357_ (.A(_12986_),
    .Y(_13315_));
 sky130_fd_sc_hd__nand2_2 _35358_ (.A(_12982_),
    .B(_12985_),
    .Y(_13316_));
 sky130_fd_sc_hd__a21boi_2 _35359_ (.A1(_13316_),
    .A2(_12989_),
    .B1_N(_12991_),
    .Y(_13317_));
 sky130_fd_sc_hd__o211a_2 _35360_ (.A1(_13315_),
    .A2(_13317_),
    .B1(_13312_),
    .C1(_13310_),
    .X(_13318_));
 sky130_fd_sc_hd__o22ai_2 _35361_ (.A1(_13290_),
    .A2(_13291_),
    .B1(_13314_),
    .B2(_13318_),
    .Y(_13319_));
 sky130_fd_sc_hd__a21o_2 _35362_ (.A1(_13310_),
    .A2(_13312_),
    .B1(_13313_),
    .X(_13320_));
 sky130_fd_sc_hd__and3_2 _35363_ (.A(_13281_),
    .B(_13285_),
    .C(_13287_),
    .X(_13321_));
 sky130_fd_sc_hd__a21oi_2 _35364_ (.A1(_13321_),
    .A2(_13279_),
    .B1(_13290_),
    .Y(_13322_));
 sky130_fd_sc_hd__nand3_2 _35365_ (.A(_13313_),
    .B(_13310_),
    .C(_13312_),
    .Y(_13323_));
 sky130_fd_sc_hd__nand3_2 _35366_ (.A(_13320_),
    .B(_13322_),
    .C(_13323_),
    .Y(_13324_));
 sky130_fd_sc_hd__nand2_2 _35367_ (.A(_12935_),
    .B(_12936_),
    .Y(_13325_));
 sky130_fd_sc_hd__a21oi_2 _35368_ (.A1(_13319_),
    .A2(_13324_),
    .B1(_13325_),
    .Y(_13326_));
 sky130_fd_sc_hd__and3_2 _35369_ (.A(_13319_),
    .B(_13325_),
    .C(_13324_),
    .X(_13327_));
 sky130_fd_sc_hd__nor2_2 _35370_ (.A(_12994_),
    .B(_13007_),
    .Y(_13328_));
 sky130_fd_sc_hd__nor2_2 _35371_ (.A(_12997_),
    .B(_13328_),
    .Y(_13329_));
 sky130_fd_sc_hd__inv_2 _35372_ (.A(_13329_),
    .Y(_13330_));
 sky130_fd_sc_hd__o21ai_2 _35373_ (.A1(_13326_),
    .A2(_13327_),
    .B1(_13330_),
    .Y(_13331_));
 sky130_fd_sc_hd__a21o_2 _35374_ (.A1(_13319_),
    .A2(_13324_),
    .B1(_13325_),
    .X(_13332_));
 sky130_fd_sc_hd__nand3_2 _35375_ (.A(_13319_),
    .B(_13325_),
    .C(_13324_),
    .Y(_13333_));
 sky130_fd_sc_hd__nand3_2 _35376_ (.A(_13332_),
    .B(_13333_),
    .C(_13329_),
    .Y(_13334_));
 sky130_fd_sc_hd__nand2_2 _35377_ (.A(_13331_),
    .B(_13334_),
    .Y(_13335_));
 sky130_fd_sc_hd__nand2_2 _35378_ (.A(_13269_),
    .B(_13335_),
    .Y(_13336_));
 sky130_fd_sc_hd__a21boi_2 _35379_ (.A1(_13016_),
    .A2(_12942_),
    .B1_N(_12950_),
    .Y(_13337_));
 sky130_fd_sc_hd__o21ai_2 _35380_ (.A1(_13326_),
    .A2(_13327_),
    .B1(_13329_),
    .Y(_13338_));
 sky130_fd_sc_hd__nand3_2 _35381_ (.A(_13330_),
    .B(_13332_),
    .C(_13333_),
    .Y(_13339_));
 sky130_fd_sc_hd__nand2_2 _35382_ (.A(_13338_),
    .B(_13339_),
    .Y(_13340_));
 sky130_fd_sc_hd__nand3_2 _35383_ (.A(_13262_),
    .B(_13340_),
    .C(_13268_),
    .Y(_13341_));
 sky130_fd_sc_hd__nand3_2 _35384_ (.A(_13336_),
    .B(_13337_),
    .C(_13341_),
    .Y(_13342_));
 sky130_fd_sc_hd__inv_2 _35385_ (.A(_13339_),
    .Y(_13343_));
 sky130_fd_sc_hd__inv_2 _35386_ (.A(_13338_),
    .Y(_13344_));
 sky130_fd_sc_hd__o2bb2ai_2 _35387_ (.A1_N(_13268_),
    .A2_N(_13262_),
    .B1(_13343_),
    .B2(_13344_),
    .Y(_13345_));
 sky130_fd_sc_hd__a21oi_2 _35388_ (.A1(_12947_),
    .A2(_12949_),
    .B1(_12944_),
    .Y(_13346_));
 sky130_fd_sc_hd__o21ai_2 _35389_ (.A1(_13022_),
    .A2(_13346_),
    .B1(_12950_),
    .Y(_13347_));
 sky130_fd_sc_hd__nand3_2 _35390_ (.A(_13262_),
    .B(_13335_),
    .C(_13268_),
    .Y(_13348_));
 sky130_fd_sc_hd__nand3_2 _35391_ (.A(_13345_),
    .B(_13347_),
    .C(_13348_),
    .Y(_13349_));
 sky130_fd_sc_hd__nand2_2 _35392_ (.A(_13342_),
    .B(_13349_),
    .Y(_13350_));
 sky130_fd_sc_hd__and3_2 _35393_ (.A(_11918_),
    .B(_19404_),
    .C(_12730_),
    .X(_13351_));
 sky130_fd_sc_hd__o21a_2 _35394_ (.A1(_13034_),
    .A2(_13351_),
    .B1(_12455_),
    .X(_13352_));
 sky130_fd_sc_hd__nor3_2 _35395_ (.A(_12455_),
    .B(_13034_),
    .C(_13351_),
    .Y(_13353_));
 sky130_fd_sc_hd__buf_1 _35396_ (.A(_13353_),
    .X(_13354_));
 sky130_fd_sc_hd__inv_2 _35397_ (.A(_13057_),
    .Y(_13355_));
 sky130_fd_sc_hd__nor2_2 _35398_ (.A(_13058_),
    .B(_13071_),
    .Y(_13356_));
 sky130_fd_sc_hd__nand2_2 _35399_ (.A(_19380_),
    .B(_19540_),
    .Y(_13357_));
 sky130_fd_sc_hd__nand2_2 _35400_ (.A(_18156_),
    .B(_06508_),
    .Y(_13358_));
 sky130_fd_sc_hd__nor2_2 _35401_ (.A(_13357_),
    .B(_13358_),
    .Y(_13359_));
 sky130_fd_sc_hd__and2_2 _35402_ (.A(_13357_),
    .B(_13358_),
    .X(_13360_));
 sky130_fd_sc_hd__buf_1 _35403_ (.A(_13360_),
    .X(_13361_));
 sky130_fd_sc_hd__o21ai_2 _35404_ (.A1(_13359_),
    .A2(_13361_),
    .B1(_13046_),
    .Y(_13362_));
 sky130_fd_sc_hd__or2_2 _35405_ (.A(_13357_),
    .B(_13358_),
    .X(_13363_));
 sky130_fd_sc_hd__nand2_2 _35406_ (.A(_13357_),
    .B(_13358_),
    .Y(_13364_));
 sky130_fd_sc_hd__nand3_2 _35407_ (.A(_13363_),
    .B(_13051_),
    .C(_13364_),
    .Y(_13365_));
 sky130_fd_sc_hd__a31o_2 _35408_ (.A1(_12966_),
    .A2(_19377_),
    .A3(_19550_),
    .B1(_12965_),
    .X(_13366_));
 sky130_fd_sc_hd__nand3_2 _35409_ (.A(_13362_),
    .B(_13365_),
    .C(_13366_),
    .Y(_13367_));
 sky130_fd_sc_hd__o21ai_2 _35410_ (.A1(_13359_),
    .A2(_13361_),
    .B1(_13051_),
    .Y(_13368_));
 sky130_fd_sc_hd__nand3_2 _35411_ (.A(_13363_),
    .B(_13046_),
    .C(_13364_),
    .Y(_13369_));
 sky130_fd_sc_hd__a21oi_2 _35412_ (.A1(_12968_),
    .A2(_12966_),
    .B1(_12965_),
    .Y(_13370_));
 sky130_fd_sc_hd__nand3_2 _35413_ (.A(_13368_),
    .B(_13369_),
    .C(_13370_),
    .Y(_13371_));
 sky130_fd_sc_hd__nor2_2 _35414_ (.A(_13051_),
    .B(_13043_),
    .Y(_13372_));
 sky130_fd_sc_hd__o2bb2ai_2 _35415_ (.A1_N(_13367_),
    .A2_N(_13371_),
    .B1(_13044_),
    .B2(_13372_),
    .Y(_13373_));
 sky130_fd_sc_hd__nor2_2 _35416_ (.A(_13044_),
    .B(_13372_),
    .Y(_13374_));
 sky130_fd_sc_hd__nand3_2 _35417_ (.A(_13367_),
    .B(_13371_),
    .C(_13374_),
    .Y(_13375_));
 sky130_fd_sc_hd__nand2_2 _35418_ (.A(_12969_),
    .B(_12970_),
    .Y(_13376_));
 sky130_fd_sc_hd__a21boi_2 _35419_ (.A1(_12958_),
    .A2(_12960_),
    .B1_N(_12952_),
    .Y(_13377_));
 sky130_fd_sc_hd__o21ai_2 _35420_ (.A1(_13376_),
    .A2(_13377_),
    .B1(_12961_),
    .Y(_13378_));
 sky130_fd_sc_hd__a21oi_2 _35421_ (.A1(_13373_),
    .A2(_13375_),
    .B1(_13378_),
    .Y(_13379_));
 sky130_fd_sc_hd__and3_2 _35422_ (.A(_13378_),
    .B(_13373_),
    .C(_13375_),
    .X(_13380_));
 sky130_fd_sc_hd__o22ai_2 _35423_ (.A1(_13355_),
    .A2(_13356_),
    .B1(_13379_),
    .B2(_13380_),
    .Y(_13381_));
 sky130_fd_sc_hd__nand2_2 _35424_ (.A(_13373_),
    .B(_13375_),
    .Y(_13382_));
 sky130_fd_sc_hd__o21a_2 _35425_ (.A1(_13376_),
    .A2(_13377_),
    .B1(_12961_),
    .X(_13383_));
 sky130_fd_sc_hd__nand2_2 _35426_ (.A(_13382_),
    .B(_13383_),
    .Y(_13384_));
 sky130_fd_sc_hd__nand3_2 _35427_ (.A(_13378_),
    .B(_13373_),
    .C(_13375_),
    .Y(_13385_));
 sky130_fd_sc_hd__nand2_2 _35428_ (.A(_13070_),
    .B(_13053_),
    .Y(_13386_));
 sky130_fd_sc_hd__nand3_2 _35429_ (.A(_13384_),
    .B(_13385_),
    .C(_13386_),
    .Y(_13387_));
 sky130_fd_sc_hd__o21ai_2 _35430_ (.A1(_13065_),
    .A2(_13061_),
    .B1(_13072_),
    .Y(_13388_));
 sky130_fd_sc_hd__a21oi_2 _35431_ (.A1(_13381_),
    .A2(_13387_),
    .B1(_13388_),
    .Y(_13389_));
 sky130_fd_sc_hd__nand2_2 _35432_ (.A(_13384_),
    .B(_13386_),
    .Y(_13390_));
 sky130_fd_sc_hd__o211a_2 _35433_ (.A1(_13380_),
    .A2(_13390_),
    .B1(_13388_),
    .C1(_13381_),
    .X(_13391_));
 sky130_fd_sc_hd__o22ai_2 _35434_ (.A1(_13352_),
    .A2(_13354_),
    .B1(_13389_),
    .B2(_13391_),
    .Y(_13392_));
 sky130_fd_sc_hd__inv_2 _35435_ (.A(_13004_),
    .Y(_13393_));
 sky130_fd_sc_hd__nand2_2 _35436_ (.A(_12998_),
    .B(_13000_),
    .Y(_13394_));
 sky130_fd_sc_hd__o2bb2ai_2 _35437_ (.A1_N(_13013_),
    .A2_N(_13014_),
    .B1(_13393_),
    .B2(_13394_),
    .Y(_13395_));
 sky130_fd_sc_hd__a21o_2 _35438_ (.A1(_13381_),
    .A2(_13387_),
    .B1(_13388_),
    .X(_13396_));
 sky130_fd_sc_hd__nor2_2 _35439_ (.A(_13353_),
    .B(_13352_),
    .Y(_13397_));
 sky130_fd_sc_hd__buf_1 _35440_ (.A(_13397_),
    .X(_13398_));
 sky130_fd_sc_hd__nand3_2 _35441_ (.A(_13381_),
    .B(_13388_),
    .C(_13387_),
    .Y(_13399_));
 sky130_fd_sc_hd__nand3_2 _35442_ (.A(_13396_),
    .B(_13398_),
    .C(_13399_),
    .Y(_13400_));
 sky130_fd_sc_hd__nand3_2 _35443_ (.A(_13392_),
    .B(_13395_),
    .C(_13400_),
    .Y(_13401_));
 sky130_fd_sc_hd__buf_1 _35444_ (.A(_13397_),
    .X(_13402_));
 sky130_fd_sc_hd__o21ai_2 _35445_ (.A1(_13389_),
    .A2(_13391_),
    .B1(_13402_),
    .Y(_13403_));
 sky130_fd_sc_hd__a21boi_2 _35446_ (.A1(_13014_),
    .A2(_13013_),
    .B1_N(_13005_),
    .Y(_13404_));
 sky130_fd_sc_hd__inv_2 _35447_ (.A(_13397_),
    .Y(_13405_));
 sky130_fd_sc_hd__buf_1 _35448_ (.A(_13405_),
    .X(_13406_));
 sky130_fd_sc_hd__nand3_2 _35449_ (.A(_13396_),
    .B(_13406_),
    .C(_13399_),
    .Y(_13407_));
 sky130_fd_sc_hd__a21oi_2 _35450_ (.A1(_13081_),
    .A2(_13082_),
    .B1(_13077_),
    .Y(_13408_));
 sky130_fd_sc_hd__a31oi_2 _35451_ (.A1(_13403_),
    .A2(_13404_),
    .A3(_13407_),
    .B1(_13408_),
    .Y(_13409_));
 sky130_fd_sc_hd__nand3_2 _35452_ (.A(_13403_),
    .B(_13404_),
    .C(_13407_),
    .Y(_13410_));
 sky130_fd_sc_hd__inv_2 _35453_ (.A(_13408_),
    .Y(_13411_));
 sky130_fd_sc_hd__a21oi_2 _35454_ (.A1(_13410_),
    .A2(_13401_),
    .B1(_13411_),
    .Y(_13412_));
 sky130_fd_sc_hd__a21oi_2 _35455_ (.A1(_13401_),
    .A2(_13409_),
    .B1(_13412_),
    .Y(_13413_));
 sky130_fd_sc_hd__nand2_2 _35456_ (.A(_13350_),
    .B(_13413_),
    .Y(_13414_));
 sky130_fd_sc_hd__a21boi_2 _35457_ (.A1(_13094_),
    .A2(_13024_),
    .B1_N(_13030_),
    .Y(_13415_));
 sky130_fd_sc_hd__and3_2 _35458_ (.A(_13410_),
    .B(_13401_),
    .C(_13411_),
    .X(_13416_));
 sky130_fd_sc_hd__o211ai_2 _35459_ (.A1(_13412_),
    .A2(_13416_),
    .B1(_13349_),
    .C1(_13342_),
    .Y(_13417_));
 sky130_fd_sc_hd__nand3_2 _35460_ (.A(_13414_),
    .B(_13415_),
    .C(_13417_),
    .Y(_13418_));
 sky130_fd_sc_hd__o2bb2ai_2 _35461_ (.A1_N(_13342_),
    .A2_N(_13349_),
    .B1(_13412_),
    .B2(_13416_),
    .Y(_13419_));
 sky130_fd_sc_hd__inv_2 _35462_ (.A(_13029_),
    .Y(_13420_));
 sky130_fd_sc_hd__nand2_2 _35463_ (.A(_13026_),
    .B(_13028_),
    .Y(_13421_));
 sky130_fd_sc_hd__a21oi_2 _35464_ (.A1(_13028_),
    .A2(_13029_),
    .B1(_13026_),
    .Y(_13422_));
 sky130_fd_sc_hd__o22ai_2 _35465_ (.A1(_13420_),
    .A2(_13421_),
    .B1(_13098_),
    .B2(_13422_),
    .Y(_13423_));
 sky130_fd_sc_hd__nand3_2 _35466_ (.A(_13413_),
    .B(_13342_),
    .C(_13349_),
    .Y(_13424_));
 sky130_fd_sc_hd__nand3_2 _35467_ (.A(_13419_),
    .B(_13423_),
    .C(_13424_),
    .Y(_13425_));
 sky130_fd_sc_hd__nor2_2 _35468_ (.A(_13351_),
    .B(_13037_),
    .Y(_13426_));
 sky130_fd_sc_hd__and3_2 _35469_ (.A(_13097_),
    .B(_13085_),
    .C(_13426_),
    .X(_13427_));
 sky130_fd_sc_hd__and2_2 _35470_ (.A(_13097_),
    .B(_13085_),
    .X(_13428_));
 sky130_fd_sc_hd__nor2_2 _35471_ (.A(_13426_),
    .B(_13428_),
    .Y(_13429_));
 sky130_fd_sc_hd__or2_2 _35472_ (.A(_13427_),
    .B(_13429_),
    .X(_13430_));
 sky130_fd_sc_hd__a21o_2 _35473_ (.A1(_13418_),
    .A2(_13425_),
    .B1(_13430_),
    .X(_13431_));
 sky130_fd_sc_hd__a21oi_2 _35474_ (.A1(_13095_),
    .A2(_13099_),
    .B1(_12841_),
    .Y(_13432_));
 sky130_fd_sc_hd__a21oi_2 _35475_ (.A1(_13114_),
    .A2(_13120_),
    .B1(_13432_),
    .Y(_13433_));
 sky130_fd_sc_hd__nand3_2 _35476_ (.A(_13430_),
    .B(_13418_),
    .C(_13425_),
    .Y(_13434_));
 sky130_fd_sc_hd__nand3_2 _35477_ (.A(_13431_),
    .B(_13433_),
    .C(_13434_),
    .Y(_13435_));
 sky130_fd_sc_hd__nor2_2 _35478_ (.A(_13427_),
    .B(_13429_),
    .Y(_13436_));
 sky130_fd_sc_hd__nand3_2 _35479_ (.A(_13418_),
    .B(_13425_),
    .C(_13436_),
    .Y(_13437_));
 sky130_fd_sc_hd__o2bb2ai_2 _35480_ (.A1_N(_13425_),
    .A2_N(_13418_),
    .B1(_13429_),
    .B2(_13427_),
    .Y(_13438_));
 sky130_fd_sc_hd__o211ai_2 _35481_ (.A1(_13432_),
    .A2(_13107_),
    .B1(_13437_),
    .C1(_13438_),
    .Y(_13439_));
 sky130_fd_sc_hd__a21oi_2 _35482_ (.A1(_13435_),
    .A2(_13439_),
    .B1(_13119_),
    .Y(_13440_));
 sky130_fd_sc_hd__and3_2 _35483_ (.A(_13435_),
    .B(_13439_),
    .C(_13119_),
    .X(_13441_));
 sky130_fd_sc_hd__o21ai_2 _35484_ (.A1(_12838_),
    .A2(_12839_),
    .B1(_13116_),
    .Y(_13442_));
 sky130_fd_sc_hd__inv_2 _35485_ (.A(_13113_),
    .Y(_13443_));
 sky130_fd_sc_hd__o2bb2ai_2 _35486_ (.A1_N(_13125_),
    .A2_N(_13124_),
    .B1(_13442_),
    .B2(_13443_),
    .Y(_13444_));
 sky130_fd_sc_hd__o21bai_2 _35487_ (.A1(_13440_),
    .A2(_13441_),
    .B1_N(_13444_),
    .Y(_13445_));
 sky130_fd_sc_hd__nand2_2 _35488_ (.A(_13435_),
    .B(_13439_),
    .Y(_13446_));
 sky130_fd_sc_hd__nand2_2 _35489_ (.A(_13446_),
    .B(_13105_),
    .Y(_13447_));
 sky130_fd_sc_hd__nand3_2 _35490_ (.A(_13435_),
    .B(_13439_),
    .C(_13119_),
    .Y(_13448_));
 sky130_fd_sc_hd__nand3_2 _35491_ (.A(_13447_),
    .B(_13444_),
    .C(_13448_),
    .Y(_13449_));
 sky130_fd_sc_hd__nand2_2 _35492_ (.A(_13445_),
    .B(_13449_),
    .Y(_13450_));
 sky130_fd_sc_hd__a21o_2 _35493_ (.A1(_13142_),
    .A2(_13133_),
    .B1(_13450_),
    .X(_13451_));
 sky130_fd_sc_hd__nand3_2 _35494_ (.A(_13142_),
    .B(_13133_),
    .C(_13450_),
    .Y(_13452_));
 sky130_fd_sc_hd__nand2_2 _35495_ (.A(_13451_),
    .B(_13452_),
    .Y(_02658_));
 sky130_fd_sc_hd__and4_2 _35496_ (.A(_19337_),
    .B(_19340_),
    .C(_07153_),
    .D(_06945_),
    .X(_13453_));
 sky130_fd_sc_hd__buf_1 _35497_ (.A(_07974_),
    .X(_13454_));
 sky130_fd_sc_hd__a22o_2 _35498_ (.A1(_10193_),
    .A2(_07380_),
    .B1(_13454_),
    .B2(_08959_),
    .X(_13455_));
 sky130_fd_sc_hd__nand2_2 _35499_ (.A(_07976_),
    .B(_09248_),
    .Y(_13456_));
 sky130_fd_sc_hd__inv_2 _35500_ (.A(_13456_),
    .Y(_13457_));
 sky130_fd_sc_hd__nand3b_2 _35501_ (.A_N(_13453_),
    .B(_13455_),
    .C(_13457_),
    .Y(_13458_));
 sky130_fd_sc_hd__a21o_2 _35502_ (.A1(_13221_),
    .A2(_13222_),
    .B1(_13217_),
    .X(_13459_));
 sky130_fd_sc_hd__a22oi_2 _35503_ (.A1(_10655_),
    .A2(_19589_),
    .B1(_13454_),
    .B2(_08959_),
    .Y(_13460_));
 sky130_fd_sc_hd__o21ai_2 _35504_ (.A1(_13460_),
    .A2(_13453_),
    .B1(_13456_),
    .Y(_13461_));
 sky130_fd_sc_hd__nand3_2 _35505_ (.A(_13458_),
    .B(_13459_),
    .C(_13461_),
    .Y(_13462_));
 sky130_fd_sc_hd__nand3b_2 _35506_ (.A_N(_13453_),
    .B(_13455_),
    .C(_13456_),
    .Y(_13463_));
 sky130_fd_sc_hd__a21oi_2 _35507_ (.A1(_13221_),
    .A2(_13222_),
    .B1(_13217_),
    .Y(_13464_));
 sky130_fd_sc_hd__o21ai_2 _35508_ (.A1(_13460_),
    .A2(_13453_),
    .B1(_13457_),
    .Y(_13465_));
 sky130_fd_sc_hd__nand3_2 _35509_ (.A(_13463_),
    .B(_13464_),
    .C(_13465_),
    .Y(_13466_));
 sky130_fd_sc_hd__nand2_2 _35510_ (.A(_07894_),
    .B(_07358_),
    .Y(_13467_));
 sky130_fd_sc_hd__nand2_2 _35511_ (.A(_07895_),
    .B(_09250_),
    .Y(_13468_));
 sky130_fd_sc_hd__nor2_2 _35512_ (.A(_13467_),
    .B(_13468_),
    .Y(_13469_));
 sky130_fd_sc_hd__and2_2 _35513_ (.A(_13467_),
    .B(_13468_),
    .X(_13470_));
 sky130_fd_sc_hd__nand2_2 _35514_ (.A(_19352_),
    .B(_08910_),
    .Y(_13471_));
 sky130_fd_sc_hd__o21bai_2 _35515_ (.A1(_13469_),
    .A2(_13470_),
    .B1_N(_13471_),
    .Y(_13472_));
 sky130_fd_sc_hd__nand2_2 _35516_ (.A(_13467_),
    .B(_13468_),
    .Y(_13473_));
 sky130_fd_sc_hd__nand3b_2 _35517_ (.A_N(_13469_),
    .B(_13471_),
    .C(_13473_),
    .Y(_13474_));
 sky130_fd_sc_hd__nand2_2 _35518_ (.A(_13472_),
    .B(_13474_),
    .Y(_13475_));
 sky130_fd_sc_hd__a21o_2 _35519_ (.A1(_13462_),
    .A2(_13466_),
    .B1(_13475_),
    .X(_13476_));
 sky130_fd_sc_hd__nand3_2 _35520_ (.A(_13462_),
    .B(_13466_),
    .C(_13475_),
    .Y(_13477_));
 sky130_fd_sc_hd__nand3_2 _35521_ (.A(_13195_),
    .B(_13199_),
    .C(_13201_),
    .Y(_13478_));
 sky130_fd_sc_hd__nand2_2 _35522_ (.A(_13478_),
    .B(_13195_),
    .Y(_13479_));
 sky130_fd_sc_hd__a21o_2 _35523_ (.A1(_13476_),
    .A2(_13477_),
    .B1(_13479_),
    .X(_13480_));
 sky130_fd_sc_hd__nand3_2 _35524_ (.A(_13479_),
    .B(_13476_),
    .C(_13477_),
    .Y(_13481_));
 sky130_fd_sc_hd__and3_2 _35525_ (.A(_13224_),
    .B(_13234_),
    .C(_13236_),
    .X(_13482_));
 sky130_fd_sc_hd__and2b_2 _35526_ (.A_N(_13482_),
    .B(_13227_),
    .X(_13483_));
 sky130_fd_sc_hd__a21oi_2 _35527_ (.A1(_13480_),
    .A2(_13481_),
    .B1(_13483_),
    .Y(_13484_));
 sky130_fd_sc_hd__nand3_2 _35528_ (.A(_13483_),
    .B(_13480_),
    .C(_13481_),
    .Y(_13485_));
 sky130_fd_sc_hd__inv_2 _35529_ (.A(_13485_),
    .Y(_13486_));
 sky130_fd_sc_hd__nand2_2 _35530_ (.A(_10138_),
    .B(_19606_),
    .Y(_13487_));
 sky130_fd_sc_hd__nand2_2 _35531_ (.A(_10141_),
    .B(_07939_),
    .Y(_13488_));
 sky130_fd_sc_hd__nor2_2 _35532_ (.A(_13487_),
    .B(_13488_),
    .Y(_13489_));
 sky130_fd_sc_hd__and2_2 _35533_ (.A(_13487_),
    .B(_13488_),
    .X(_13490_));
 sky130_fd_sc_hd__nor2_2 _35534_ (.A(_09357_),
    .B(_07313_),
    .Y(_13491_));
 sky130_fd_sc_hd__inv_2 _35535_ (.A(_13491_),
    .Y(_13492_));
 sky130_fd_sc_hd__o21ai_2 _35536_ (.A1(_13489_),
    .A2(_13490_),
    .B1(_13492_),
    .Y(_13493_));
 sky130_fd_sc_hd__inv_2 _35537_ (.A(_13493_),
    .Y(_13494_));
 sky130_fd_sc_hd__or2_2 _35538_ (.A(_13487_),
    .B(_13488_),
    .X(_13495_));
 sky130_fd_sc_hd__nand2_2 _35539_ (.A(_13487_),
    .B(_13488_),
    .Y(_13496_));
 sky130_fd_sc_hd__nand3_2 _35540_ (.A(_13495_),
    .B(_13491_),
    .C(_13496_),
    .Y(_13497_));
 sky130_fd_sc_hd__inv_2 _35541_ (.A(_13497_),
    .Y(_13498_));
 sky130_fd_sc_hd__nand3_2 _35542_ (.A(_10818_),
    .B(_10699_),
    .C(_05734_),
    .Y(_13499_));
 sky130_fd_sc_hd__nor2_2 _35543_ (.A(_05893_),
    .B(_13499_),
    .Y(_13500_));
 sky130_fd_sc_hd__nand2_2 _35544_ (.A(_13146_),
    .B(_07210_),
    .Y(_13501_));
 sky130_fd_sc_hd__o21a_2 _35545_ (.A1(_05893_),
    .A2(_10830_),
    .B1(_13501_),
    .X(_13502_));
 sky130_fd_sc_hd__nor2_2 _35546_ (.A(_10150_),
    .B(_06694_),
    .Y(_13503_));
 sky130_fd_sc_hd__o21bai_2 _35547_ (.A1(_13500_),
    .A2(_13502_),
    .B1_N(_13503_),
    .Y(_13504_));
 sky130_fd_sc_hd__o21ai_2 _35548_ (.A1(_19617_),
    .A2(_18182_),
    .B1(_13501_),
    .Y(_13505_));
 sky130_fd_sc_hd__nand3b_2 _35549_ (.A_N(_13500_),
    .B(_13505_),
    .C(_13503_),
    .Y(_13506_));
 sky130_fd_sc_hd__a21o_2 _35550_ (.A1(_13152_),
    .A2(_13153_),
    .B1(_13145_),
    .X(_13507_));
 sky130_fd_sc_hd__a21oi_2 _35551_ (.A1(_13504_),
    .A2(_13506_),
    .B1(_13507_),
    .Y(_13508_));
 sky130_fd_sc_hd__o21ai_2 _35552_ (.A1(_19617_),
    .A2(_13499_),
    .B1(_13503_),
    .Y(_13509_));
 sky130_fd_sc_hd__o211a_2 _35553_ (.A1(_13502_),
    .A2(_13509_),
    .B1(_13504_),
    .C1(_13507_),
    .X(_13510_));
 sky130_fd_sc_hd__o22ai_2 _35554_ (.A1(_13494_),
    .A2(_13498_),
    .B1(_13508_),
    .B2(_13510_),
    .Y(_13511_));
 sky130_fd_sc_hd__o21ai_2 _35555_ (.A1(_13177_),
    .A2(_13155_),
    .B1(_13173_),
    .Y(_13512_));
 sky130_fd_sc_hd__a21o_2 _35556_ (.A1(_13504_),
    .A2(_13506_),
    .B1(_13507_),
    .X(_13513_));
 sky130_fd_sc_hd__and2_2 _35557_ (.A(_13493_),
    .B(_13497_),
    .X(_13514_));
 sky130_fd_sc_hd__nand3_2 _35558_ (.A(_13507_),
    .B(_13504_),
    .C(_13506_),
    .Y(_13515_));
 sky130_fd_sc_hd__nand3_2 _35559_ (.A(_13513_),
    .B(_13514_),
    .C(_13515_),
    .Y(_13516_));
 sky130_fd_sc_hd__nand3_2 _35560_ (.A(_13511_),
    .B(_13512_),
    .C(_13516_),
    .Y(_13517_));
 sky130_fd_sc_hd__o21ai_2 _35561_ (.A1(_13508_),
    .A2(_13510_),
    .B1(_13514_),
    .Y(_13518_));
 sky130_fd_sc_hd__a21oi_2 _35562_ (.A1(_13174_),
    .A2(_13170_),
    .B1(_13159_),
    .Y(_13519_));
 sky130_fd_sc_hd__nand2_2 _35563_ (.A(_13493_),
    .B(_13497_),
    .Y(_13520_));
 sky130_fd_sc_hd__nand3_2 _35564_ (.A(_13513_),
    .B(_13515_),
    .C(_13520_),
    .Y(_13521_));
 sky130_fd_sc_hd__nand3_2 _35565_ (.A(_13518_),
    .B(_13519_),
    .C(_13521_),
    .Y(_13522_));
 sky130_fd_sc_hd__nand2_2 _35566_ (.A(_09819_),
    .B(_07143_),
    .Y(_13523_));
 sky130_fd_sc_hd__nand2_2 _35567_ (.A(_09827_),
    .B(_19594_),
    .Y(_13524_));
 sky130_fd_sc_hd__nor2_2 _35568_ (.A(_13523_),
    .B(_13524_),
    .Y(_13525_));
 sky130_fd_sc_hd__and2_2 _35569_ (.A(_13523_),
    .B(_13524_),
    .X(_13526_));
 sky130_fd_sc_hd__nor2_2 _35570_ (.A(_08423_),
    .B(_10268_),
    .Y(_13527_));
 sky130_fd_sc_hd__o21bai_2 _35571_ (.A1(_13525_),
    .A2(_13526_),
    .B1_N(_13527_),
    .Y(_13528_));
 sky130_fd_sc_hd__or2_2 _35572_ (.A(_13523_),
    .B(_13524_),
    .X(_13529_));
 sky130_fd_sc_hd__nand2_2 _35573_ (.A(_13523_),
    .B(_13524_),
    .Y(_13530_));
 sky130_fd_sc_hd__nand3_2 _35574_ (.A(_13529_),
    .B(_13527_),
    .C(_13530_),
    .Y(_13531_));
 sky130_fd_sc_hd__a31o_2 _35575_ (.A1(_13163_),
    .A2(_19324_),
    .A3(_19604_),
    .B1(_13162_),
    .X(_13532_));
 sky130_fd_sc_hd__a21o_2 _35576_ (.A1(_13528_),
    .A2(_13531_),
    .B1(_13532_),
    .X(_13533_));
 sky130_fd_sc_hd__nand3_2 _35577_ (.A(_13528_),
    .B(_13531_),
    .C(_13532_),
    .Y(_13534_));
 sky130_fd_sc_hd__nor2_2 _35578_ (.A(_13189_),
    .B(_13188_),
    .Y(_13535_));
 sky130_fd_sc_hd__nor2_2 _35579_ (.A(_13187_),
    .B(_13535_),
    .Y(_13536_));
 sky130_fd_sc_hd__inv_2 _35580_ (.A(_13536_),
    .Y(_13537_));
 sky130_fd_sc_hd__a21oi_2 _35581_ (.A1(_13533_),
    .A2(_13534_),
    .B1(_13537_),
    .Y(_13538_));
 sky130_fd_sc_hd__and3_2 _35582_ (.A(_13533_),
    .B(_13537_),
    .C(_13534_),
    .X(_13539_));
 sky130_fd_sc_hd__o2bb2ai_2 _35583_ (.A1_N(_13517_),
    .A2_N(_13522_),
    .B1(_13538_),
    .B2(_13539_),
    .Y(_13540_));
 sky130_fd_sc_hd__nand2_2 _35584_ (.A(_13533_),
    .B(_13534_),
    .Y(_13541_));
 sky130_fd_sc_hd__a21oi_2 _35585_ (.A1(_13528_),
    .A2(_13531_),
    .B1(_13532_),
    .Y(_13542_));
 sky130_fd_sc_hd__nand2_2 _35586_ (.A(_13534_),
    .B(_13536_),
    .Y(_13543_));
 sky130_fd_sc_hd__o2bb2ai_2 _35587_ (.A1_N(_13541_),
    .A2_N(_13537_),
    .B1(_13542_),
    .B2(_13543_),
    .Y(_13544_));
 sky130_fd_sc_hd__nand3_2 _35588_ (.A(_13544_),
    .B(_13522_),
    .C(_13517_),
    .Y(_13545_));
 sky130_fd_sc_hd__nand2_2 _35589_ (.A(_13212_),
    .B(_13184_),
    .Y(_13546_));
 sky130_fd_sc_hd__a21oi_2 _35590_ (.A1(_13540_),
    .A2(_13545_),
    .B1(_13546_),
    .Y(_13547_));
 sky130_fd_sc_hd__nand2_2 _35591_ (.A(_13203_),
    .B(_13200_),
    .Y(_13548_));
 sky130_fd_sc_hd__nand2_2 _35592_ (.A(_13548_),
    .B(_13478_),
    .Y(_13549_));
 sky130_fd_sc_hd__a31oi_2 _35593_ (.A1(_13171_),
    .A2(_13172_),
    .A3(_13178_),
    .B1(_13549_),
    .Y(_13550_));
 sky130_fd_sc_hd__o211a_2 _35594_ (.A1(_13211_),
    .A2(_13550_),
    .B1(_13545_),
    .C1(_13540_),
    .X(_13551_));
 sky130_fd_sc_hd__o22ai_2 _35595_ (.A1(_13484_),
    .A2(_13486_),
    .B1(_13547_),
    .B2(_13551_),
    .Y(_13552_));
 sky130_fd_sc_hd__a21oi_2 _35596_ (.A1(_13476_),
    .A2(_13477_),
    .B1(_13479_),
    .Y(_13553_));
 sky130_fd_sc_hd__and3_2 _35597_ (.A(_13479_),
    .B(_13476_),
    .C(_13477_),
    .X(_13554_));
 sky130_fd_sc_hd__a31o_2 _35598_ (.A1(_13214_),
    .A2(_13225_),
    .A3(_13226_),
    .B1(_13482_),
    .X(_13555_));
 sky130_fd_sc_hd__o21ai_2 _35599_ (.A1(_13553_),
    .A2(_13554_),
    .B1(_13555_),
    .Y(_13556_));
 sky130_fd_sc_hd__nand2_2 _35600_ (.A(_13556_),
    .B(_13485_),
    .Y(_13557_));
 sky130_fd_sc_hd__a21oi_2 _35601_ (.A1(_13522_),
    .A2(_13517_),
    .B1(_13544_),
    .Y(_13558_));
 sky130_fd_sc_hd__a21oi_2 _35602_ (.A1(_13533_),
    .A2(_13534_),
    .B1(_13536_),
    .Y(_13559_));
 sky130_fd_sc_hd__nor2_2 _35603_ (.A(_13542_),
    .B(_13543_),
    .Y(_13560_));
 sky130_fd_sc_hd__o211a_2 _35604_ (.A1(_13559_),
    .A2(_13560_),
    .B1(_13517_),
    .C1(_13522_),
    .X(_13561_));
 sky130_fd_sc_hd__nor2_2 _35605_ (.A(_13211_),
    .B(_13550_),
    .Y(_13562_));
 sky130_fd_sc_hd__o21ai_2 _35606_ (.A1(_13558_),
    .A2(_13561_),
    .B1(_13562_),
    .Y(_13563_));
 sky130_fd_sc_hd__nand3_2 _35607_ (.A(_13546_),
    .B(_13540_),
    .C(_13545_),
    .Y(_13564_));
 sky130_fd_sc_hd__nand3b_2 _35608_ (.A_N(_13557_),
    .B(_13563_),
    .C(_13564_),
    .Y(_13565_));
 sky130_fd_sc_hd__o21ai_2 _35609_ (.A1(_13260_),
    .A2(_13210_),
    .B1(_13254_),
    .Y(_13566_));
 sky130_fd_sc_hd__a21oi_2 _35610_ (.A1(_13552_),
    .A2(_13565_),
    .B1(_13566_),
    .Y(_13567_));
 sky130_fd_sc_hd__a21oi_2 _35611_ (.A1(_13251_),
    .A2(_13252_),
    .B1(_13260_),
    .Y(_13568_));
 sky130_fd_sc_hd__o211a_2 _35612_ (.A1(_13213_),
    .A2(_13568_),
    .B1(_13565_),
    .C1(_13552_),
    .X(_13569_));
 sky130_fd_sc_hd__nand2_2 _35613_ (.A(_06624_),
    .B(\pcpi_mul.rs1[26] ),
    .Y(_13570_));
 sky130_fd_sc_hd__nand2_2 _35614_ (.A(_07015_),
    .B(_19557_),
    .Y(_13571_));
 sky130_fd_sc_hd__nor2_2 _35615_ (.A(_13570_),
    .B(_13571_),
    .Y(_13572_));
 sky130_fd_sc_hd__and2_2 _35616_ (.A(_13570_),
    .B(_13571_),
    .X(_13573_));
 sky130_fd_sc_hd__nor2_2 _35617_ (.A(_06118_),
    .B(_10542_),
    .Y(_13574_));
 sky130_fd_sc_hd__o21bai_2 _35618_ (.A1(_13572_),
    .A2(_13573_),
    .B1_N(_13574_),
    .Y(_13575_));
 sky130_fd_sc_hd__nand2_2 _35619_ (.A(_13570_),
    .B(_13571_),
    .Y(_13576_));
 sky130_fd_sc_hd__nand3b_2 _35620_ (.A_N(_13572_),
    .B(_13574_),
    .C(_13576_),
    .Y(_13577_));
 sky130_fd_sc_hd__a21o_2 _35621_ (.A1(_13271_),
    .A2(_13272_),
    .B1(_13270_),
    .X(_13578_));
 sky130_fd_sc_hd__a21oi_2 _35622_ (.A1(_13575_),
    .A2(_13577_),
    .B1(_13578_),
    .Y(_13579_));
 sky130_fd_sc_hd__nand3_2 _35623_ (.A(_13578_),
    .B(_13575_),
    .C(_13577_),
    .Y(_13580_));
 sky130_fd_sc_hd__inv_2 _35624_ (.A(_13580_),
    .Y(_13581_));
 sky130_fd_sc_hd__nor2_2 _35625_ (.A(_13579_),
    .B(_13581_),
    .Y(_13582_));
 sky130_fd_sc_hd__nand2_2 _35626_ (.A(_05956_),
    .B(_19548_),
    .Y(_13583_));
 sky130_fd_sc_hd__nand2_2 _35627_ (.A(_07034_),
    .B(_19544_),
    .Y(_13584_));
 sky130_fd_sc_hd__nor2_2 _35628_ (.A(_13583_),
    .B(_13584_),
    .Y(_13585_));
 sky130_fd_sc_hd__and2_2 _35629_ (.A(_13583_),
    .B(_13584_),
    .X(_13586_));
 sky130_fd_sc_hd__nand2_2 _35630_ (.A(_06616_),
    .B(_11901_),
    .Y(_13587_));
 sky130_fd_sc_hd__o21ai_2 _35631_ (.A1(_13585_),
    .A2(_13586_),
    .B1(_13587_),
    .Y(_13588_));
 sky130_fd_sc_hd__inv_2 _35632_ (.A(_13587_),
    .Y(_13589_));
 sky130_fd_sc_hd__nand2_2 _35633_ (.A(_13583_),
    .B(_13584_),
    .Y(_13590_));
 sky130_fd_sc_hd__nand3b_2 _35634_ (.A_N(_13585_),
    .B(_13589_),
    .C(_13590_),
    .Y(_13591_));
 sky130_fd_sc_hd__and2_2 _35635_ (.A(_13588_),
    .B(_13591_),
    .X(_13592_));
 sky130_fd_sc_hd__nand2_2 _35636_ (.A(_13582_),
    .B(_13592_),
    .Y(_13593_));
 sky130_fd_sc_hd__a21o_2 _35637_ (.A1(_13575_),
    .A2(_13577_),
    .B1(_13578_),
    .X(_13594_));
 sky130_fd_sc_hd__buf_1 _35638_ (.A(_13580_),
    .X(_13595_));
 sky130_fd_sc_hd__a21o_2 _35639_ (.A1(_13594_),
    .A2(_13595_),
    .B1(_13592_),
    .X(_13596_));
 sky130_fd_sc_hd__nand2_2 _35640_ (.A(_08182_),
    .B(_08085_),
    .Y(_13597_));
 sky130_fd_sc_hd__nand2_2 _35641_ (.A(_07652_),
    .B(_08661_),
    .Y(_13598_));
 sky130_fd_sc_hd__nor2_2 _35642_ (.A(_13597_),
    .B(_13598_),
    .Y(_13599_));
 sky130_fd_sc_hd__and2_2 _35643_ (.A(_13597_),
    .B(_13598_),
    .X(_13600_));
 sky130_fd_sc_hd__nor2_2 _35644_ (.A(_06831_),
    .B(_11671_),
    .Y(_13601_));
 sky130_fd_sc_hd__o21bai_2 _35645_ (.A1(_13599_),
    .A2(_13600_),
    .B1_N(_13601_),
    .Y(_13602_));
 sky130_fd_sc_hd__nand2_2 _35646_ (.A(_13597_),
    .B(_13598_),
    .Y(_13603_));
 sky130_fd_sc_hd__nand3b_2 _35647_ (.A_N(_13599_),
    .B(_13601_),
    .C(_13603_),
    .Y(_13604_));
 sky130_fd_sc_hd__a31o_2 _35648_ (.A1(_13231_),
    .A2(_12069_),
    .A3(_07845_),
    .B1(_13230_),
    .X(_13605_));
 sky130_fd_sc_hd__a21oi_2 _35649_ (.A1(_13602_),
    .A2(_13604_),
    .B1(_13605_),
    .Y(_13606_));
 sky130_fd_sc_hd__nand3_2 _35650_ (.A(_13602_),
    .B(_13605_),
    .C(_13604_),
    .Y(_13607_));
 sky130_fd_sc_hd__a21oi_2 _35651_ (.A1(_13301_),
    .A2(_13300_),
    .B1(_13296_),
    .Y(_13608_));
 sky130_fd_sc_hd__nand2_2 _35652_ (.A(_13607_),
    .B(_13608_),
    .Y(_13609_));
 sky130_fd_sc_hd__a21boi_2 _35653_ (.A1(_13307_),
    .A2(_13311_),
    .B1_N(_13303_),
    .Y(_13610_));
 sky130_fd_sc_hd__and3_2 _35654_ (.A(_13602_),
    .B(_13605_),
    .C(_13604_),
    .X(_13611_));
 sky130_fd_sc_hd__inv_2 _35655_ (.A(_13608_),
    .Y(_13612_));
 sky130_fd_sc_hd__o21ai_2 _35656_ (.A1(_13606_),
    .A2(_13611_),
    .B1(_13612_),
    .Y(_13613_));
 sky130_fd_sc_hd__o211ai_2 _35657_ (.A1(_13606_),
    .A2(_13609_),
    .B1(_13610_),
    .C1(_13613_),
    .Y(_13614_));
 sky130_fd_sc_hd__o21ai_2 _35658_ (.A1(_13606_),
    .A2(_13611_),
    .B1(_13608_),
    .Y(_13615_));
 sky130_fd_sc_hd__nand2_2 _35659_ (.A(_13312_),
    .B(_13303_),
    .Y(_13616_));
 sky130_fd_sc_hd__nand3b_2 _35660_ (.A_N(_13606_),
    .B(_13607_),
    .C(_13612_),
    .Y(_13617_));
 sky130_fd_sc_hd__nand3_2 _35661_ (.A(_13615_),
    .B(_13616_),
    .C(_13617_),
    .Y(_13618_));
 sky130_fd_sc_hd__a22oi_2 _35662_ (.A1(_13593_),
    .A2(_13596_),
    .B1(_13614_),
    .B2(_13618_),
    .Y(_13619_));
 sky130_fd_sc_hd__nand2_2 _35663_ (.A(_13588_),
    .B(_13591_),
    .Y(_13620_));
 sky130_fd_sc_hd__a21oi_2 _35664_ (.A1(_13594_),
    .A2(_13595_),
    .B1(_13620_),
    .Y(_13621_));
 sky130_fd_sc_hd__and3_2 _35665_ (.A(_13594_),
    .B(_13595_),
    .C(_13620_),
    .X(_13622_));
 sky130_fd_sc_hd__o211a_2 _35666_ (.A1(_13621_),
    .A2(_13622_),
    .B1(_13618_),
    .C1(_13614_),
    .X(_13623_));
 sky130_fd_sc_hd__a21oi_2 _35667_ (.A1(_13242_),
    .A2(_13245_),
    .B1(_13255_),
    .Y(_13624_));
 sky130_fd_sc_hd__o21ai_2 _35668_ (.A1(_13619_),
    .A2(_13623_),
    .B1(_13624_),
    .Y(_13625_));
 sky130_fd_sc_hd__a22o_2 _35669_ (.A1(_13593_),
    .A2(_13596_),
    .B1(_13614_),
    .B2(_13618_),
    .X(_13626_));
 sky130_fd_sc_hd__o21ai_2 _35670_ (.A1(_13257_),
    .A2(_13258_),
    .B1(_13243_),
    .Y(_13627_));
 sky130_fd_sc_hd__nand2_2 _35671_ (.A(_13582_),
    .B(_13620_),
    .Y(_13628_));
 sky130_fd_sc_hd__a21o_2 _35672_ (.A1(_13594_),
    .A2(_13595_),
    .B1(_13620_),
    .X(_13629_));
 sky130_fd_sc_hd__nand2_2 _35673_ (.A(_13628_),
    .B(_13629_),
    .Y(_13630_));
 sky130_fd_sc_hd__nand3_2 _35674_ (.A(_13630_),
    .B(_13614_),
    .C(_13618_),
    .Y(_13631_));
 sky130_fd_sc_hd__nand3_2 _35675_ (.A(_13626_),
    .B(_13627_),
    .C(_13631_),
    .Y(_13632_));
 sky130_fd_sc_hd__nand2_2 _35676_ (.A(_13324_),
    .B(_13323_),
    .Y(_13633_));
 sky130_fd_sc_hd__a21o_2 _35677_ (.A1(_13625_),
    .A2(_13632_),
    .B1(_13633_),
    .X(_13634_));
 sky130_fd_sc_hd__buf_1 _35678_ (.A(_13632_),
    .X(_13635_));
 sky130_fd_sc_hd__nand3_2 _35679_ (.A(_13625_),
    .B(_13635_),
    .C(_13633_),
    .Y(_13636_));
 sky130_fd_sc_hd__nand2_2 _35680_ (.A(_13634_),
    .B(_13636_),
    .Y(_13637_));
 sky130_fd_sc_hd__o21ai_2 _35681_ (.A1(_13567_),
    .A2(_13569_),
    .B1(_13637_),
    .Y(_13638_));
 sky130_fd_sc_hd__nand2_2 _35682_ (.A(_13262_),
    .B(_13335_),
    .Y(_13639_));
 sky130_fd_sc_hd__nand2_2 _35683_ (.A(_13639_),
    .B(_13268_),
    .Y(_13640_));
 sky130_fd_sc_hd__a22oi_2 _35684_ (.A1(_13556_),
    .A2(_13485_),
    .B1(_13563_),
    .B2(_13564_),
    .Y(_13641_));
 sky130_fd_sc_hd__nor3_2 _35685_ (.A(_13557_),
    .B(_13547_),
    .C(_13551_),
    .Y(_13642_));
 sky130_fd_sc_hd__o21bai_2 _35686_ (.A1(_13641_),
    .A2(_13642_),
    .B1_N(_13566_),
    .Y(_13643_));
 sky130_fd_sc_hd__nand3_2 _35687_ (.A(_13552_),
    .B(_13566_),
    .C(_13565_),
    .Y(_13644_));
 sky130_fd_sc_hd__inv_2 _35688_ (.A(_13633_),
    .Y(_13645_));
 sky130_fd_sc_hd__a21oi_2 _35689_ (.A1(_13626_),
    .A2(_13631_),
    .B1(_13627_),
    .Y(_13646_));
 sky130_fd_sc_hd__nor2_2 _35690_ (.A(_13645_),
    .B(_13646_),
    .Y(_13647_));
 sky130_fd_sc_hd__a21oi_2 _35691_ (.A1(_13625_),
    .A2(_13635_),
    .B1(_13633_),
    .Y(_13648_));
 sky130_fd_sc_hd__a21oi_2 _35692_ (.A1(_13647_),
    .A2(_13635_),
    .B1(_13648_),
    .Y(_13649_));
 sky130_fd_sc_hd__nand3_2 _35693_ (.A(_13643_),
    .B(_13644_),
    .C(_13649_),
    .Y(_13650_));
 sky130_fd_sc_hd__nand3_2 _35694_ (.A(_13638_),
    .B(_13640_),
    .C(_13650_),
    .Y(_13651_));
 sky130_fd_sc_hd__a21oi_2 _35695_ (.A1(_13625_),
    .A2(_13635_),
    .B1(_13645_),
    .Y(_13652_));
 sky130_fd_sc_hd__and3_2 _35696_ (.A(_13625_),
    .B(_13645_),
    .C(_13635_),
    .X(_13653_));
 sky130_fd_sc_hd__o22ai_2 _35697_ (.A1(_13652_),
    .A2(_13653_),
    .B1(_13567_),
    .B2(_13569_),
    .Y(_13654_));
 sky130_fd_sc_hd__a21boi_2 _35698_ (.A1(_13262_),
    .A2(_13335_),
    .B1_N(_13268_),
    .Y(_13655_));
 sky130_fd_sc_hd__nand3_2 _35699_ (.A(_13643_),
    .B(_13644_),
    .C(_13637_),
    .Y(_13656_));
 sky130_fd_sc_hd__nand3_2 _35700_ (.A(_13654_),
    .B(_13655_),
    .C(_13656_),
    .Y(_13657_));
 sky130_fd_sc_hd__nand2_2 _35701_ (.A(_13651_),
    .B(_13657_),
    .Y(_13658_));
 sky130_fd_sc_hd__a21oi_2 _35702_ (.A1(_13283_),
    .A2(_13284_),
    .B1(_13282_),
    .Y(_13659_));
 sky130_fd_sc_hd__o21a_2 _35703_ (.A1(_05447_),
    .A2(_19382_),
    .B1(\pcpi_mul.rs1[32] ),
    .X(_13660_));
 sky130_fd_sc_hd__nand3_2 _35704_ (.A(_11759_),
    .B(_19379_),
    .C(_06334_),
    .Y(_13661_));
 sky130_fd_sc_hd__nand2_2 _35705_ (.A(_13660_),
    .B(_13661_),
    .Y(_13662_));
 sky130_fd_sc_hd__nand2_2 _35706_ (.A(_13662_),
    .B(_13050_),
    .Y(_13663_));
 sky130_fd_sc_hd__nand3_2 _35707_ (.A(_13660_),
    .B(_13046_),
    .C(_13661_),
    .Y(_13664_));
 sky130_fd_sc_hd__nand3_2 _35708_ (.A(_13659_),
    .B(_13663_),
    .C(_13664_),
    .Y(_13665_));
 sky130_fd_sc_hd__a21o_2 _35709_ (.A1(_13283_),
    .A2(_13284_),
    .B1(_13282_),
    .X(_13666_));
 sky130_fd_sc_hd__nand2_2 _35710_ (.A(_13662_),
    .B(_13046_),
    .Y(_13667_));
 sky130_fd_sc_hd__nand3_2 _35711_ (.A(_13050_),
    .B(_13660_),
    .C(_13661_),
    .Y(_13668_));
 sky130_fd_sc_hd__buf_1 _35712_ (.A(_13668_),
    .X(_13669_));
 sky130_fd_sc_hd__nand3_2 _35713_ (.A(_13666_),
    .B(_13667_),
    .C(_13669_),
    .Y(_13670_));
 sky130_fd_sc_hd__nor2_2 _35714_ (.A(_13051_),
    .B(_13359_),
    .Y(_13671_));
 sky130_fd_sc_hd__o2bb2ai_2 _35715_ (.A1_N(_13665_),
    .A2_N(_13670_),
    .B1(_13361_),
    .B2(_13671_),
    .Y(_13672_));
 sky130_fd_sc_hd__nor2_2 _35716_ (.A(_13361_),
    .B(_13671_),
    .Y(_13673_));
 sky130_fd_sc_hd__nand3_2 _35717_ (.A(_13670_),
    .B(_13665_),
    .C(_13673_),
    .Y(_13674_));
 sky130_fd_sc_hd__a21oi_2 _35718_ (.A1(_13273_),
    .A2(_13276_),
    .B1(_13280_),
    .Y(_13675_));
 sky130_fd_sc_hd__o21ai_2 _35719_ (.A1(_13288_),
    .A2(_13675_),
    .B1(_13281_),
    .Y(_13676_));
 sky130_fd_sc_hd__a21oi_2 _35720_ (.A1(_13672_),
    .A2(_13674_),
    .B1(_13676_),
    .Y(_13677_));
 sky130_fd_sc_hd__inv_2 _35721_ (.A(_13665_),
    .Y(_13678_));
 sky130_fd_sc_hd__nand2_2 _35722_ (.A(_13670_),
    .B(_13673_),
    .Y(_13679_));
 sky130_fd_sc_hd__o211a_2 _35723_ (.A1(_13678_),
    .A2(_13679_),
    .B1(_13672_),
    .C1(_13676_),
    .X(_13680_));
 sky130_fd_sc_hd__a21bo_2 _35724_ (.A1(_13371_),
    .A2(_13374_),
    .B1_N(_13367_),
    .X(_13681_));
 sky130_fd_sc_hd__o21bai_2 _35725_ (.A1(_13677_),
    .A2(_13680_),
    .B1_N(_13681_),
    .Y(_13682_));
 sky130_fd_sc_hd__a21o_2 _35726_ (.A1(_13672_),
    .A2(_13674_),
    .B1(_13676_),
    .X(_13683_));
 sky130_fd_sc_hd__nand3_2 _35727_ (.A(_13676_),
    .B(_13674_),
    .C(_13672_),
    .Y(_13684_));
 sky130_fd_sc_hd__nand3_2 _35728_ (.A(_13683_),
    .B(_13684_),
    .C(_13681_),
    .Y(_13685_));
 sky130_fd_sc_hd__inv_2 _35729_ (.A(_13386_),
    .Y(_13686_));
 sky130_fd_sc_hd__o21ai_2 _35730_ (.A1(_13686_),
    .A2(_13379_),
    .B1(_13385_),
    .Y(_13687_));
 sky130_fd_sc_hd__a21oi_2 _35731_ (.A1(_13682_),
    .A2(_13685_),
    .B1(_13687_),
    .Y(_13688_));
 sky130_fd_sc_hd__a21oi_2 _35732_ (.A1(_13382_),
    .A2(_13383_),
    .B1(_13686_),
    .Y(_13689_));
 sky130_fd_sc_hd__o211a_2 _35733_ (.A1(_13380_),
    .A2(_13689_),
    .B1(_13685_),
    .C1(_13682_),
    .X(_13690_));
 sky130_fd_sc_hd__o21ai_2 _35734_ (.A1(_13688_),
    .A2(_13690_),
    .B1(_13398_),
    .Y(_13691_));
 sky130_fd_sc_hd__nand2_2 _35735_ (.A(_13333_),
    .B(_13329_),
    .Y(_13692_));
 sky130_fd_sc_hd__nand2_2 _35736_ (.A(_13692_),
    .B(_13332_),
    .Y(_13693_));
 sky130_fd_sc_hd__a21o_2 _35737_ (.A1(_13682_),
    .A2(_13685_),
    .B1(_13687_),
    .X(_13694_));
 sky130_fd_sc_hd__nand3_2 _35738_ (.A(_13682_),
    .B(_13687_),
    .C(_13685_),
    .Y(_13695_));
 sky130_fd_sc_hd__nand3_2 _35739_ (.A(_13694_),
    .B(_13406_),
    .C(_13695_),
    .Y(_13696_));
 sky130_fd_sc_hd__nand3_2 _35740_ (.A(_13691_),
    .B(_13693_),
    .C(_13696_),
    .Y(_13697_));
 sky130_fd_sc_hd__o22ai_2 _35741_ (.A1(_13352_),
    .A2(_13354_),
    .B1(_13688_),
    .B2(_13690_),
    .Y(_13698_));
 sky130_fd_sc_hd__inv_2 _35742_ (.A(_13324_),
    .Y(_13699_));
 sky130_fd_sc_hd__nand2_2 _35743_ (.A(_13319_),
    .B(_13325_),
    .Y(_13700_));
 sky130_fd_sc_hd__o22ai_2 _35744_ (.A1(_13699_),
    .A2(_13700_),
    .B1(_13329_),
    .B2(_13326_),
    .Y(_13701_));
 sky130_fd_sc_hd__buf_1 _35745_ (.A(_13397_),
    .X(_13702_));
 sky130_fd_sc_hd__nand3_2 _35746_ (.A(_13694_),
    .B(_13702_),
    .C(_13695_),
    .Y(_13703_));
 sky130_fd_sc_hd__nand3_2 _35747_ (.A(_13698_),
    .B(_13701_),
    .C(_13703_),
    .Y(_13704_));
 sky130_fd_sc_hd__nand2_2 _35748_ (.A(_13396_),
    .B(_13398_),
    .Y(_13705_));
 sky130_fd_sc_hd__nand2_2 _35749_ (.A(_13705_),
    .B(_13399_),
    .Y(_13706_));
 sky130_fd_sc_hd__a21oi_2 _35750_ (.A1(_13697_),
    .A2(_13704_),
    .B1(_13706_),
    .Y(_13707_));
 sky130_fd_sc_hd__and3_2 _35751_ (.A(_13697_),
    .B(_13704_),
    .C(_13706_),
    .X(_13708_));
 sky130_fd_sc_hd__nor2_2 _35752_ (.A(_13707_),
    .B(_13708_),
    .Y(_13709_));
 sky130_fd_sc_hd__nand2_2 _35753_ (.A(_13658_),
    .B(_13709_),
    .Y(_13710_));
 sky130_fd_sc_hd__nand2_2 _35754_ (.A(_13697_),
    .B(_13704_),
    .Y(_13711_));
 sky130_fd_sc_hd__inv_2 _35755_ (.A(_13706_),
    .Y(_13712_));
 sky130_fd_sc_hd__nand2_2 _35756_ (.A(_13711_),
    .B(_13712_),
    .Y(_13713_));
 sky130_fd_sc_hd__nand3_2 _35757_ (.A(_13697_),
    .B(_13704_),
    .C(_13706_),
    .Y(_13714_));
 sky130_fd_sc_hd__nand2_2 _35758_ (.A(_13713_),
    .B(_13714_),
    .Y(_13715_));
 sky130_fd_sc_hd__nand3_2 _35759_ (.A(_13651_),
    .B(_13657_),
    .C(_13715_),
    .Y(_13716_));
 sky130_fd_sc_hd__a21boi_2 _35760_ (.A1(_13413_),
    .A2(_13342_),
    .B1_N(_13349_),
    .Y(_13717_));
 sky130_fd_sc_hd__nand3_2 _35761_ (.A(_13710_),
    .B(_13716_),
    .C(_13717_),
    .Y(_13718_));
 sky130_fd_sc_hd__nand2_2 _35762_ (.A(_13658_),
    .B(_13715_),
    .Y(_13719_));
 sky130_fd_sc_hd__nand2_2 _35763_ (.A(_13413_),
    .B(_13342_),
    .Y(_13720_));
 sky130_fd_sc_hd__nand2_2 _35764_ (.A(_13720_),
    .B(_13349_),
    .Y(_13721_));
 sky130_fd_sc_hd__nand3_2 _35765_ (.A(_13651_),
    .B(_13657_),
    .C(_13709_),
    .Y(_13722_));
 sky130_fd_sc_hd__nand3_2 _35766_ (.A(_13719_),
    .B(_13721_),
    .C(_13722_),
    .Y(_13723_));
 sky130_fd_sc_hd__nor2_2 _35767_ (.A(_13351_),
    .B(_13354_),
    .Y(_13724_));
 sky130_fd_sc_hd__buf_1 _35768_ (.A(_13724_),
    .X(_13725_));
 sky130_fd_sc_hd__and2b_2 _35769_ (.A_N(_13409_),
    .B(_13401_),
    .X(_13726_));
 sky130_fd_sc_hd__nor2_2 _35770_ (.A(_13725_),
    .B(_13726_),
    .Y(_13727_));
 sky130_fd_sc_hd__and2_2 _35771_ (.A(_13726_),
    .B(_13725_),
    .X(_13728_));
 sky130_fd_sc_hd__o2bb2ai_2 _35772_ (.A1_N(_13718_),
    .A2_N(_13723_),
    .B1(_13727_),
    .B2(_13728_),
    .Y(_13729_));
 sky130_fd_sc_hd__nand2_2 _35773_ (.A(_13418_),
    .B(_13436_),
    .Y(_13730_));
 sky130_fd_sc_hd__nand2_2 _35774_ (.A(_13730_),
    .B(_13425_),
    .Y(_13731_));
 sky130_fd_sc_hd__nor2_2 _35775_ (.A(_13727_),
    .B(_13728_),
    .Y(_13732_));
 sky130_fd_sc_hd__nand3_2 _35776_ (.A(_13723_),
    .B(_13718_),
    .C(_13732_),
    .Y(_13733_));
 sky130_fd_sc_hd__nand3_2 _35777_ (.A(_13729_),
    .B(_13731_),
    .C(_13733_),
    .Y(_13734_));
 sky130_fd_sc_hd__inv_2 _35778_ (.A(_13724_),
    .Y(_13735_));
 sky130_fd_sc_hd__buf_1 _35779_ (.A(_13735_),
    .X(_13736_));
 sky130_fd_sc_hd__buf_1 _35780_ (.A(_13736_),
    .X(_13737_));
 sky130_fd_sc_hd__nor2_2 _35781_ (.A(_13737_),
    .B(_13726_),
    .Y(_13738_));
 sky130_fd_sc_hd__and2_2 _35782_ (.A(_13726_),
    .B(_13736_),
    .X(_13739_));
 sky130_fd_sc_hd__o2bb2ai_2 _35783_ (.A1_N(_13718_),
    .A2_N(_13723_),
    .B1(_13738_),
    .B2(_13739_),
    .Y(_13740_));
 sky130_fd_sc_hd__nand3b_2 _35784_ (.A_N(_13732_),
    .B(_13723_),
    .C(_13718_),
    .Y(_13741_));
 sky130_fd_sc_hd__a21boi_2 _35785_ (.A1(_13418_),
    .A2(_13436_),
    .B1_N(_13425_),
    .Y(_13742_));
 sky130_fd_sc_hd__nand3_2 _35786_ (.A(_13740_),
    .B(_13741_),
    .C(_13742_),
    .Y(_13743_));
 sky130_fd_sc_hd__inv_2 _35787_ (.A(_13429_),
    .Y(_13744_));
 sky130_fd_sc_hd__a21o_2 _35788_ (.A1(_13734_),
    .A2(_13743_),
    .B1(_13744_),
    .X(_13745_));
 sky130_fd_sc_hd__a21boi_2 _35789_ (.A1(_13435_),
    .A2(_13119_),
    .B1_N(_13439_),
    .Y(_13746_));
 sky130_fd_sc_hd__nand3_2 _35790_ (.A(_13734_),
    .B(_13743_),
    .C(_13744_),
    .Y(_13747_));
 sky130_fd_sc_hd__nand3_2 _35791_ (.A(_13745_),
    .B(_13746_),
    .C(_13747_),
    .Y(_13748_));
 sky130_fd_sc_hd__nand2_2 _35792_ (.A(_13435_),
    .B(_13119_),
    .Y(_13749_));
 sky130_fd_sc_hd__nand2_2 _35793_ (.A(_13749_),
    .B(_13439_),
    .Y(_13750_));
 sky130_fd_sc_hd__o2bb2ai_2 _35794_ (.A1_N(_13743_),
    .A2_N(_13734_),
    .B1(_13426_),
    .B2(_13428_),
    .Y(_13751_));
 sky130_fd_sc_hd__nand3_2 _35795_ (.A(_13734_),
    .B(_13743_),
    .C(_13429_),
    .Y(_13752_));
 sky130_fd_sc_hd__nand3_2 _35796_ (.A(_13750_),
    .B(_13751_),
    .C(_13752_),
    .Y(_13753_));
 sky130_fd_sc_hd__nand2_2 _35797_ (.A(_13748_),
    .B(_13753_),
    .Y(_13754_));
 sky130_fd_sc_hd__a21oi_2 _35798_ (.A1(_13117_),
    .A2(_13124_),
    .B1(_13125_),
    .Y(_13755_));
 sky130_fd_sc_hd__o21ai_2 _35799_ (.A1(_12836_),
    .A2(_12837_),
    .B1(_13126_),
    .Y(_13756_));
 sky130_fd_sc_hd__o2111a_2 _35800_ (.A1(_13755_),
    .A2(_13756_),
    .B1(_13133_),
    .C1(_13449_),
    .D1(_13445_),
    .X(_13757_));
 sky130_fd_sc_hd__nand3_2 _35801_ (.A(_13757_),
    .B(_12513_),
    .C(_12833_),
    .Y(_13758_));
 sky130_fd_sc_hd__nand2_2 _35802_ (.A(_11855_),
    .B(_12188_),
    .Y(_13759_));
 sky130_fd_sc_hd__nor2_2 _35803_ (.A(_13758_),
    .B(_13759_),
    .Y(_13760_));
 sky130_fd_sc_hd__o2111ai_2 _35804_ (.A1(_13755_),
    .A2(_13756_),
    .B1(_13449_),
    .C1(_13133_),
    .D1(_13445_),
    .Y(_13761_));
 sky130_fd_sc_hd__a21oi_2 _35805_ (.A1(_13447_),
    .A2(_13448_),
    .B1(_13444_),
    .Y(_13762_));
 sky130_fd_sc_hd__o21a_2 _35806_ (.A1(_13128_),
    .A2(_13762_),
    .B1(_13449_),
    .X(_13763_));
 sky130_fd_sc_hd__o21ai_2 _35807_ (.A1(_13136_),
    .A2(_13761_),
    .B1(_13763_),
    .Y(_13764_));
 sky130_fd_sc_hd__o21bai_2 _35808_ (.A1(_13758_),
    .A2(_12516_),
    .B1_N(_13764_),
    .Y(_13765_));
 sky130_fd_sc_hd__a21oi_2 _35809_ (.A1(_11157_),
    .A2(_13760_),
    .B1(_13765_),
    .Y(_13766_));
 sky130_fd_sc_hd__or2_2 _35810_ (.A(_13754_),
    .B(_13766_),
    .X(_13767_));
 sky130_fd_sc_hd__nand2_2 _35811_ (.A(_13766_),
    .B(_13754_),
    .Y(_13768_));
 sky130_fd_sc_hd__and2_2 _35812_ (.A(_13767_),
    .B(_13768_),
    .X(_02659_));
 sky130_fd_sc_hd__nand2_2 _35813_ (.A(_13714_),
    .B(_13704_),
    .Y(_13769_));
 sky130_fd_sc_hd__inv_2 _35814_ (.A(_13769_),
    .Y(_13770_));
 sky130_fd_sc_hd__nor2_2 _35815_ (.A(_13725_),
    .B(_13770_),
    .Y(_13771_));
 sky130_fd_sc_hd__buf_1 _35816_ (.A(_13771_),
    .X(_13772_));
 sky130_fd_sc_hd__nor2_2 _35817_ (.A(_13736_),
    .B(_13769_),
    .Y(_13773_));
 sky130_fd_sc_hd__o21ai_2 _35818_ (.A1(_13637_),
    .A2(_13567_),
    .B1(_13644_),
    .Y(_13774_));
 sky130_fd_sc_hd__nand2_2 _35819_ (.A(_07898_),
    .B(_08661_),
    .Y(_13775_));
 sky130_fd_sc_hd__nand2_2 _35820_ (.A(_08345_),
    .B(_19564_),
    .Y(_13776_));
 sky130_fd_sc_hd__or2_2 _35821_ (.A(_13775_),
    .B(_13776_),
    .X(_13777_));
 sky130_fd_sc_hd__nor2_2 _35822_ (.A(_08352_),
    .B(_10513_),
    .Y(_13778_));
 sky130_fd_sc_hd__nand2_2 _35823_ (.A(_13775_),
    .B(_13776_),
    .Y(_13779_));
 sky130_fd_sc_hd__nand3_2 _35824_ (.A(_13777_),
    .B(_13778_),
    .C(_13779_),
    .Y(_13780_));
 sky130_fd_sc_hd__a21o_2 _35825_ (.A1(_09009_),
    .A2(_10380_),
    .B1(_13775_),
    .X(_13781_));
 sky130_fd_sc_hd__a21o_2 _35826_ (.A1(_09008_),
    .A2(_08662_),
    .B1(_13776_),
    .X(_13782_));
 sky130_fd_sc_hd__o211ai_2 _35827_ (.A1(_11300_),
    .A2(_10514_),
    .B1(_13781_),
    .C1(_13782_),
    .Y(_13783_));
 sky130_fd_sc_hd__a31o_2 _35828_ (.A1(_13473_),
    .A2(_12069_),
    .A3(_08910_),
    .B1(_13469_),
    .X(_13784_));
 sky130_fd_sc_hd__a21oi_2 _35829_ (.A1(_13780_),
    .A2(_13783_),
    .B1(_13784_),
    .Y(_13785_));
 sky130_fd_sc_hd__a21oi_2 _35830_ (.A1(_13467_),
    .A2(_13468_),
    .B1(_13471_),
    .Y(_13786_));
 sky130_fd_sc_hd__o211a_2 _35831_ (.A1(_13469_),
    .A2(_13786_),
    .B1(_13783_),
    .C1(_13780_),
    .X(_13787_));
 sky130_fd_sc_hd__a31o_2 _35832_ (.A1(_13603_),
    .A2(_19360_),
    .A3(_19566_),
    .B1(_13599_),
    .X(_13788_));
 sky130_fd_sc_hd__o21bai_2 _35833_ (.A1(_13785_),
    .A2(_13787_),
    .B1_N(_13788_),
    .Y(_13789_));
 sky130_fd_sc_hd__a21o_2 _35834_ (.A1(_13780_),
    .A2(_13783_),
    .B1(_13784_),
    .X(_13790_));
 sky130_fd_sc_hd__nand3_2 _35835_ (.A(_13780_),
    .B(_13784_),
    .C(_13783_),
    .Y(_13791_));
 sky130_fd_sc_hd__nand3_2 _35836_ (.A(_13790_),
    .B(_13791_),
    .C(_13788_),
    .Y(_13792_));
 sky130_fd_sc_hd__o21ai_2 _35837_ (.A1(_13608_),
    .A2(_13606_),
    .B1(_13607_),
    .Y(_13793_));
 sky130_fd_sc_hd__a21oi_2 _35838_ (.A1(_13789_),
    .A2(_13792_),
    .B1(_13793_),
    .Y(_13794_));
 sky130_fd_sc_hd__and3_2 _35839_ (.A(_13789_),
    .B(_13793_),
    .C(_13792_),
    .X(_13795_));
 sky130_fd_sc_hd__nand2_2 _35840_ (.A(_19363_),
    .B(_19557_),
    .Y(_13796_));
 sky130_fd_sc_hd__nand2_2 _35841_ (.A(_07020_),
    .B(_19552_),
    .Y(_13797_));
 sky130_fd_sc_hd__nor2_2 _35842_ (.A(_13796_),
    .B(_13797_),
    .Y(_13798_));
 sky130_fd_sc_hd__and2_2 _35843_ (.A(_13796_),
    .B(_13797_),
    .X(_13799_));
 sky130_fd_sc_hd__nor2_2 _35844_ (.A(_06119_),
    .B(_10532_),
    .Y(_13800_));
 sky130_fd_sc_hd__o21bai_2 _35845_ (.A1(_13798_),
    .A2(_13799_),
    .B1_N(_13800_),
    .Y(_13801_));
 sky130_fd_sc_hd__nand2_2 _35846_ (.A(_13796_),
    .B(_13797_),
    .Y(_13802_));
 sky130_fd_sc_hd__nand3b_2 _35847_ (.A_N(_13798_),
    .B(_13800_),
    .C(_13802_),
    .Y(_13803_));
 sky130_fd_sc_hd__nand2_2 _35848_ (.A(_13801_),
    .B(_13803_),
    .Y(_13804_));
 sky130_fd_sc_hd__a21oi_2 _35849_ (.A1(_13574_),
    .A2(_13576_),
    .B1(_13572_),
    .Y(_13805_));
 sky130_fd_sc_hd__nand2_2 _35850_ (.A(_13804_),
    .B(_13805_),
    .Y(_13806_));
 sky130_fd_sc_hd__nand3b_2 _35851_ (.A_N(_13805_),
    .B(_13801_),
    .C(_13803_),
    .Y(_13807_));
 sky130_fd_sc_hd__a22oi_2 _35852_ (.A1(_05801_),
    .A2(_10537_),
    .B1(_08331_),
    .B2(_11427_),
    .Y(_13808_));
 sky130_fd_sc_hd__nand2_2 _35853_ (.A(_11023_),
    .B(_19375_),
    .Y(_13809_));
 sky130_fd_sc_hd__inv_2 _35854_ (.A(_13809_),
    .Y(_13810_));
 sky130_fd_sc_hd__and4_2 _35855_ (.A(_05807_),
    .B(_05808_),
    .C(_11427_),
    .D(_10537_),
    .X(_13811_));
 sky130_fd_sc_hd__nor3_2 _35856_ (.A(_13808_),
    .B(_13810_),
    .C(_13811_),
    .Y(_13812_));
 sky130_fd_sc_hd__o21a_2 _35857_ (.A1(_13808_),
    .A2(_13811_),
    .B1(_13810_),
    .X(_13813_));
 sky130_fd_sc_hd__nor2_2 _35858_ (.A(_13812_),
    .B(_13813_),
    .Y(_13814_));
 sky130_fd_sc_hd__a21o_2 _35859_ (.A1(_13806_),
    .A2(_13807_),
    .B1(_13814_),
    .X(_13815_));
 sky130_fd_sc_hd__nand3_2 _35860_ (.A(_13806_),
    .B(_13807_),
    .C(_13814_),
    .Y(_13816_));
 sky130_fd_sc_hd__nand2_2 _35861_ (.A(_13815_),
    .B(_13816_),
    .Y(_13817_));
 sky130_fd_sc_hd__o21bai_2 _35862_ (.A1(_13794_),
    .A2(_13795_),
    .B1_N(_13817_),
    .Y(_13818_));
 sky130_fd_sc_hd__a21o_2 _35863_ (.A1(_13789_),
    .A2(_13792_),
    .B1(_13793_),
    .X(_13819_));
 sky130_fd_sc_hd__nand3_2 _35864_ (.A(_13789_),
    .B(_13793_),
    .C(_13792_),
    .Y(_13820_));
 sky130_fd_sc_hd__nand3_2 _35865_ (.A(_13819_),
    .B(_13817_),
    .C(_13820_),
    .Y(_13821_));
 sky130_fd_sc_hd__o21ai_2 _35866_ (.A1(_13553_),
    .A2(_13555_),
    .B1(_13481_),
    .Y(_13822_));
 sky130_fd_sc_hd__a21o_2 _35867_ (.A1(_13818_),
    .A2(_13821_),
    .B1(_13822_),
    .X(_13823_));
 sky130_fd_sc_hd__nand3_2 _35868_ (.A(_13818_),
    .B(_13822_),
    .C(_13821_),
    .Y(_13824_));
 sky130_fd_sc_hd__nand2_2 _35869_ (.A(_13630_),
    .B(_13614_),
    .Y(_13825_));
 sky130_fd_sc_hd__nand2_2 _35870_ (.A(_13825_),
    .B(_13618_),
    .Y(_13826_));
 sky130_fd_sc_hd__and3_2 _35871_ (.A(_13823_),
    .B(_13824_),
    .C(_13826_),
    .X(_13827_));
 sky130_fd_sc_hd__a21oi_2 _35872_ (.A1(_13823_),
    .A2(_13824_),
    .B1(_13826_),
    .Y(_13828_));
 sky130_fd_sc_hd__o21a_2 _35873_ (.A1(_13520_),
    .A2(_13508_),
    .B1(_13515_),
    .X(_13829_));
 sky130_fd_sc_hd__nand2_2 _35874_ (.A(_19315_),
    .B(_07939_),
    .Y(_13830_));
 sky130_fd_sc_hd__nand2_2 _35875_ (.A(_09602_),
    .B(_07311_),
    .Y(_13831_));
 sky130_fd_sc_hd__nor2_2 _35876_ (.A(_13830_),
    .B(_13831_),
    .Y(_13832_));
 sky130_fd_sc_hd__inv_2 _35877_ (.A(_13832_),
    .Y(_13833_));
 sky130_fd_sc_hd__nand2_2 _35878_ (.A(_19323_),
    .B(_06388_),
    .Y(_13834_));
 sky130_fd_sc_hd__nand2_2 _35879_ (.A(_13830_),
    .B(_13831_),
    .Y(_13835_));
 sky130_fd_sc_hd__and3_2 _35880_ (.A(_13833_),
    .B(_13834_),
    .C(_13835_),
    .X(_13836_));
 sky130_fd_sc_hd__inv_2 _35881_ (.A(_13835_),
    .Y(_13837_));
 sky130_fd_sc_hd__nor2_2 _35882_ (.A(_13832_),
    .B(_13837_),
    .Y(_13838_));
 sky130_fd_sc_hd__nor2_2 _35883_ (.A(_13834_),
    .B(_13838_),
    .Y(_13839_));
 sky130_fd_sc_hd__nand2_2 _35884_ (.A(_19307_),
    .B(_05598_),
    .Y(_13840_));
 sky130_fd_sc_hd__nand3b_2 _35885_ (.A_N(_13840_),
    .B(_10824_),
    .C(_06494_),
    .Y(_13841_));
 sky130_fd_sc_hd__o21ai_2 _35886_ (.A1(_05737_),
    .A2(_11509_),
    .B1(_13840_),
    .Y(_13842_));
 sky130_fd_sc_hd__o2bb2ai_2 _35887_ (.A1_N(_13841_),
    .A2_N(_13842_),
    .B1(_10151_),
    .B2(_06225_),
    .Y(_13843_));
 sky130_fd_sc_hd__nor2_2 _35888_ (.A(_10150_),
    .B(_06224_),
    .Y(_13844_));
 sky130_fd_sc_hd__nand3_2 _35889_ (.A(_13841_),
    .B(_13842_),
    .C(_13844_),
    .Y(_13845_));
 sky130_fd_sc_hd__a21o_2 _35890_ (.A1(_13505_),
    .A2(_13503_),
    .B1(_13500_),
    .X(_13846_));
 sky130_fd_sc_hd__a21oi_2 _35891_ (.A1(_13843_),
    .A2(_13845_),
    .B1(_13846_),
    .Y(_13847_));
 sky130_fd_sc_hd__buf_1 _35892_ (.A(_11509_),
    .X(_13848_));
 sky130_fd_sc_hd__o21a_2 _35893_ (.A1(_19614_),
    .A2(_13848_),
    .B1(_13840_),
    .X(_13849_));
 sky130_fd_sc_hd__nand2_2 _35894_ (.A(_13841_),
    .B(_13844_),
    .Y(_13850_));
 sky130_fd_sc_hd__o211a_2 _35895_ (.A1(_13849_),
    .A2(_13850_),
    .B1(_13846_),
    .C1(_13843_),
    .X(_13851_));
 sky130_fd_sc_hd__o22ai_2 _35896_ (.A1(_13836_),
    .A2(_13839_),
    .B1(_13847_),
    .B2(_13851_),
    .Y(_13852_));
 sky130_fd_sc_hd__a21o_2 _35897_ (.A1(_13843_),
    .A2(_13845_),
    .B1(_13846_),
    .X(_13853_));
 sky130_fd_sc_hd__nand3_2 _35898_ (.A(_13843_),
    .B(_13846_),
    .C(_13845_),
    .Y(_13854_));
 sky130_fd_sc_hd__inv_2 _35899_ (.A(_13834_),
    .Y(_13855_));
 sky130_fd_sc_hd__nand2_2 _35900_ (.A(_13838_),
    .B(_13855_),
    .Y(_13856_));
 sky130_fd_sc_hd__o21ai_2 _35901_ (.A1(_13832_),
    .A2(_13837_),
    .B1(_13834_),
    .Y(_13857_));
 sky130_fd_sc_hd__nand2_2 _35902_ (.A(_13856_),
    .B(_13857_),
    .Y(_13858_));
 sky130_fd_sc_hd__nand3_2 _35903_ (.A(_13853_),
    .B(_13854_),
    .C(_13858_),
    .Y(_13859_));
 sky130_fd_sc_hd__nand3_2 _35904_ (.A(_13829_),
    .B(_13852_),
    .C(_13859_),
    .Y(_13860_));
 sky130_fd_sc_hd__o2bb2ai_2 _35905_ (.A1_N(_13856_),
    .A2_N(_13857_),
    .B1(_13847_),
    .B2(_13851_),
    .Y(_13861_));
 sky130_fd_sc_hd__o211ai_2 _35906_ (.A1(_13836_),
    .A2(_13839_),
    .B1(_13854_),
    .C1(_13853_),
    .Y(_13862_));
 sky130_fd_sc_hd__o21ai_2 _35907_ (.A1(_13520_),
    .A2(_13508_),
    .B1(_13515_),
    .Y(_13863_));
 sky130_fd_sc_hd__nand3_2 _35908_ (.A(_13861_),
    .B(_13862_),
    .C(_13863_),
    .Y(_13864_));
 sky130_fd_sc_hd__nand2_2 _35909_ (.A(_13860_),
    .B(_13864_),
    .Y(_13865_));
 sky130_fd_sc_hd__a21oi_2 _35910_ (.A1(_13491_),
    .A2(_13496_),
    .B1(_13489_),
    .Y(_13866_));
 sky130_fd_sc_hd__and4_2 _35911_ (.A(_19328_),
    .B(_10156_),
    .C(_06950_),
    .D(_06557_),
    .X(_13867_));
 sky130_fd_sc_hd__inv_2 _35912_ (.A(_09120_),
    .Y(_13868_));
 sky130_fd_sc_hd__nand2_2 _35913_ (.A(_11205_),
    .B(_06954_),
    .Y(_13869_));
 sky130_fd_sc_hd__o21a_2 _35914_ (.A1(_13868_),
    .A2(_10268_),
    .B1(_13869_),
    .X(_13870_));
 sky130_fd_sc_hd__nand2_2 _35915_ (.A(_10862_),
    .B(_07380_),
    .Y(_13871_));
 sky130_fd_sc_hd__o21ai_2 _35916_ (.A1(_13867_),
    .A2(_13870_),
    .B1(_13871_),
    .Y(_13872_));
 sky130_fd_sc_hd__buf_1 _35917_ (.A(_13868_),
    .X(_13873_));
 sky130_fd_sc_hd__o21ai_2 _35918_ (.A1(_13873_),
    .A2(_10279_),
    .B1(_13869_),
    .Y(_13874_));
 sky130_fd_sc_hd__inv_2 _35919_ (.A(_13871_),
    .Y(_13875_));
 sky130_fd_sc_hd__nand3b_2 _35920_ (.A_N(_13867_),
    .B(_13874_),
    .C(_13875_),
    .Y(_13876_));
 sky130_fd_sc_hd__nand3b_2 _35921_ (.A_N(_13866_),
    .B(_13872_),
    .C(_13876_),
    .Y(_13877_));
 sky130_fd_sc_hd__o21ai_2 _35922_ (.A1(_13867_),
    .A2(_13870_),
    .B1(_13875_),
    .Y(_13878_));
 sky130_fd_sc_hd__nand3b_2 _35923_ (.A_N(_13867_),
    .B(_13874_),
    .C(_13871_),
    .Y(_13879_));
 sky130_fd_sc_hd__nand3_2 _35924_ (.A(_13878_),
    .B(_13866_),
    .C(_13879_),
    .Y(_13880_));
 sky130_fd_sc_hd__nand2_2 _35925_ (.A(_13531_),
    .B(_13529_),
    .Y(_13881_));
 sky130_fd_sc_hd__a21oi_2 _35926_ (.A1(_13877_),
    .A2(_13880_),
    .B1(_13881_),
    .Y(_13882_));
 sky130_fd_sc_hd__and3_2 _35927_ (.A(_13877_),
    .B(_13880_),
    .C(_13881_),
    .X(_13883_));
 sky130_fd_sc_hd__nor2_2 _35928_ (.A(_13882_),
    .B(_13883_),
    .Y(_13884_));
 sky130_fd_sc_hd__nand2_2 _35929_ (.A(_13865_),
    .B(_13884_),
    .Y(_13885_));
 sky130_fd_sc_hd__a21boi_2 _35930_ (.A1(_13544_),
    .A2(_13522_),
    .B1_N(_13517_),
    .Y(_13886_));
 sky130_fd_sc_hd__nand3_2 _35931_ (.A(_13877_),
    .B(_13880_),
    .C(_13881_),
    .Y(_13887_));
 sky130_fd_sc_hd__or2b_2 _35932_ (.A(_13882_),
    .B_N(_13887_),
    .X(_13888_));
 sky130_fd_sc_hd__nand3_2 _35933_ (.A(_13888_),
    .B(_13860_),
    .C(_13864_),
    .Y(_13889_));
 sky130_fd_sc_hd__nand3_2 _35934_ (.A(_13885_),
    .B(_13886_),
    .C(_13889_),
    .Y(_13890_));
 sky130_fd_sc_hd__nand2_2 _35935_ (.A(_13865_),
    .B(_13888_),
    .Y(_13891_));
 sky130_fd_sc_hd__inv_2 _35936_ (.A(_13516_),
    .Y(_13892_));
 sky130_fd_sc_hd__nand2_2 _35937_ (.A(_13511_),
    .B(_13512_),
    .Y(_13893_));
 sky130_fd_sc_hd__o2bb2ai_2 _35938_ (.A1_N(_13522_),
    .A2_N(_13544_),
    .B1(_13892_),
    .B2(_13893_),
    .Y(_13894_));
 sky130_fd_sc_hd__nand3_2 _35939_ (.A(_13884_),
    .B(_13860_),
    .C(_13864_),
    .Y(_13895_));
 sky130_fd_sc_hd__nand3_2 _35940_ (.A(_13891_),
    .B(_13894_),
    .C(_13895_),
    .Y(_13896_));
 sky130_fd_sc_hd__nor2_2 _35941_ (.A(_13456_),
    .B(_13460_),
    .Y(_13897_));
 sky130_fd_sc_hd__nand2_2 _35942_ (.A(_08391_),
    .B(_07156_),
    .Y(_13898_));
 sky130_fd_sc_hd__nand2_2 _35943_ (.A(_08386_),
    .B(_07377_),
    .Y(_13899_));
 sky130_fd_sc_hd__nor2_2 _35944_ (.A(_13898_),
    .B(_13899_),
    .Y(_13900_));
 sky130_fd_sc_hd__nand2_2 _35945_ (.A(_13898_),
    .B(_13899_),
    .Y(_13901_));
 sky130_fd_sc_hd__nand2_2 _35946_ (.A(_07976_),
    .B(_07590_),
    .Y(_13902_));
 sky130_fd_sc_hd__inv_2 _35947_ (.A(_13902_),
    .Y(_13903_));
 sky130_fd_sc_hd__nand3b_2 _35948_ (.A_N(_13900_),
    .B(_13901_),
    .C(_13903_),
    .Y(_13904_));
 sky130_fd_sc_hd__and2_2 _35949_ (.A(_13898_),
    .B(_13899_),
    .X(_13905_));
 sky130_fd_sc_hd__o21ai_2 _35950_ (.A1(_13900_),
    .A2(_13905_),
    .B1(_13902_),
    .Y(_13906_));
 sky130_fd_sc_hd__o211ai_2 _35951_ (.A1(_13453_),
    .A2(_13897_),
    .B1(_13904_),
    .C1(_13906_),
    .Y(_13907_));
 sky130_fd_sc_hd__o21ai_2 _35952_ (.A1(_13900_),
    .A2(_13905_),
    .B1(_13903_),
    .Y(_13908_));
 sky130_fd_sc_hd__nand3b_2 _35953_ (.A_N(_13900_),
    .B(_13901_),
    .C(_13902_),
    .Y(_13909_));
 sky130_fd_sc_hd__a21oi_2 _35954_ (.A1(_13455_),
    .A2(_13457_),
    .B1(_13453_),
    .Y(_13910_));
 sky130_fd_sc_hd__nand3_2 _35955_ (.A(_13908_),
    .B(_13909_),
    .C(_13910_),
    .Y(_13911_));
 sky130_fd_sc_hd__nand2_2 _35956_ (.A(_19347_),
    .B(_09250_),
    .Y(_13912_));
 sky130_fd_sc_hd__nand2_2 _35957_ (.A(_08159_),
    .B(_08103_),
    .Y(_13913_));
 sky130_fd_sc_hd__nor2_2 _35958_ (.A(_13912_),
    .B(_13913_),
    .Y(_13914_));
 sky130_fd_sc_hd__nor2_2 _35959_ (.A(_11251_),
    .B(_12088_),
    .Y(_13915_));
 sky130_fd_sc_hd__inv_2 _35960_ (.A(_13915_),
    .Y(_13916_));
 sky130_fd_sc_hd__nand2_2 _35961_ (.A(_13912_),
    .B(_13913_),
    .Y(_13917_));
 sky130_fd_sc_hd__nand3b_2 _35962_ (.A_N(_13914_),
    .B(_13916_),
    .C(_13917_),
    .Y(_13918_));
 sky130_fd_sc_hd__and2_2 _35963_ (.A(_13912_),
    .B(_13913_),
    .X(_13919_));
 sky130_fd_sc_hd__o21ai_2 _35964_ (.A1(_13914_),
    .A2(_13919_),
    .B1(_13915_),
    .Y(_13920_));
 sky130_fd_sc_hd__nand2_2 _35965_ (.A(_13918_),
    .B(_13920_),
    .Y(_13921_));
 sky130_fd_sc_hd__a21oi_2 _35966_ (.A1(_13907_),
    .A2(_13911_),
    .B1(_13921_),
    .Y(_13922_));
 sky130_fd_sc_hd__and3_2 _35967_ (.A(_13921_),
    .B(_13907_),
    .C(_13911_),
    .X(_13923_));
 sky130_fd_sc_hd__o2bb2ai_2 _35968_ (.A1_N(_13533_),
    .A2_N(_13543_),
    .B1(_13922_),
    .B2(_13923_),
    .Y(_13924_));
 sky130_fd_sc_hd__o21ai_2 _35969_ (.A1(_13536_),
    .A2(_13542_),
    .B1(_13534_),
    .Y(_13925_));
 sky130_fd_sc_hd__nand3_2 _35970_ (.A(_13921_),
    .B(_13907_),
    .C(_13911_),
    .Y(_13926_));
 sky130_fd_sc_hd__nand3b_2 _35971_ (.A_N(_13922_),
    .B(_13925_),
    .C(_13926_),
    .Y(_13927_));
 sky130_fd_sc_hd__inv_2 _35972_ (.A(_13462_),
    .Y(_13928_));
 sky130_fd_sc_hd__and2_2 _35973_ (.A(_13466_),
    .B(_13475_),
    .X(_13929_));
 sky130_fd_sc_hd__or2_2 _35974_ (.A(_13928_),
    .B(_13929_),
    .X(_13930_));
 sky130_fd_sc_hd__a21oi_2 _35975_ (.A1(_13924_),
    .A2(_13927_),
    .B1(_13930_),
    .Y(_13931_));
 sky130_fd_sc_hd__o211a_2 _35976_ (.A1(_13928_),
    .A2(_13929_),
    .B1(_13927_),
    .C1(_13924_),
    .X(_13932_));
 sky130_fd_sc_hd__o2bb2ai_2 _35977_ (.A1_N(_13890_),
    .A2_N(_13896_),
    .B1(_13931_),
    .B2(_13932_),
    .Y(_13933_));
 sky130_fd_sc_hd__nor2_2 _35978_ (.A(_13931_),
    .B(_13932_),
    .Y(_13934_));
 sky130_fd_sc_hd__nand3_2 _35979_ (.A(_13934_),
    .B(_13896_),
    .C(_13890_),
    .Y(_13935_));
 sky130_fd_sc_hd__nand2_2 _35980_ (.A(_13546_),
    .B(_13540_),
    .Y(_13936_));
 sky130_fd_sc_hd__o22ai_2 _35981_ (.A1(_13561_),
    .A2(_13936_),
    .B1(_13557_),
    .B2(_13547_),
    .Y(_13937_));
 sky130_fd_sc_hd__a21oi_2 _35982_ (.A1(_13933_),
    .A2(_13935_),
    .B1(_13937_),
    .Y(_13938_));
 sky130_fd_sc_hd__and3_2 _35983_ (.A(_13891_),
    .B(_13894_),
    .C(_13895_),
    .X(_13939_));
 sky130_fd_sc_hd__nand2_2 _35984_ (.A(_13934_),
    .B(_13890_),
    .Y(_13940_));
 sky130_fd_sc_hd__o211a_2 _35985_ (.A1(_13939_),
    .A2(_13940_),
    .B1(_13937_),
    .C1(_13933_),
    .X(_13941_));
 sky130_fd_sc_hd__o22ai_2 _35986_ (.A1(_13827_),
    .A2(_13828_),
    .B1(_13938_),
    .B2(_13941_),
    .Y(_13942_));
 sky130_fd_sc_hd__and2_2 _35987_ (.A(_13825_),
    .B(_13618_),
    .X(_13943_));
 sky130_fd_sc_hd__a21oi_2 _35988_ (.A1(_13818_),
    .A2(_13821_),
    .B1(_13822_),
    .Y(_13944_));
 sky130_fd_sc_hd__nor2_2 _35989_ (.A(_13943_),
    .B(_13944_),
    .Y(_13945_));
 sky130_fd_sc_hd__a21oi_2 _35990_ (.A1(_13824_),
    .A2(_13945_),
    .B1(_13828_),
    .Y(_13946_));
 sky130_fd_sc_hd__nand3_2 _35991_ (.A(_13933_),
    .B(_13937_),
    .C(_13935_),
    .Y(_13947_));
 sky130_fd_sc_hd__a21o_2 _35992_ (.A1(_13933_),
    .A2(_13935_),
    .B1(_13937_),
    .X(_13948_));
 sky130_fd_sc_hd__nand3_2 _35993_ (.A(_13946_),
    .B(_13947_),
    .C(_13948_),
    .Y(_13949_));
 sky130_fd_sc_hd__nand3_2 _35994_ (.A(_13774_),
    .B(_13942_),
    .C(_13949_),
    .Y(_13950_));
 sky130_fd_sc_hd__a21oi_2 _35995_ (.A1(_13643_),
    .A2(_13649_),
    .B1(_13569_),
    .Y(_13951_));
 sky130_fd_sc_hd__o21ai_2 _35996_ (.A1(_13938_),
    .A2(_13941_),
    .B1(_13946_),
    .Y(_13952_));
 sky130_fd_sc_hd__inv_2 _35997_ (.A(_13824_),
    .Y(_13953_));
 sky130_fd_sc_hd__o21ai_2 _35998_ (.A1(_13944_),
    .A2(_13953_),
    .B1(_13943_),
    .Y(_13954_));
 sky130_fd_sc_hd__nand2_2 _35999_ (.A(_13945_),
    .B(_13824_),
    .Y(_13955_));
 sky130_fd_sc_hd__nand2_2 _36000_ (.A(_13954_),
    .B(_13955_),
    .Y(_13956_));
 sky130_fd_sc_hd__nand3_2 _36001_ (.A(_13956_),
    .B(_13948_),
    .C(_13947_),
    .Y(_13957_));
 sky130_fd_sc_hd__nand3_2 _36002_ (.A(_13951_),
    .B(_13952_),
    .C(_13957_),
    .Y(_13958_));
 sky130_fd_sc_hd__a21oi_2 _36003_ (.A1(_13583_),
    .A2(_13584_),
    .B1(_13587_),
    .Y(_13959_));
 sky130_fd_sc_hd__nor2_2 _36004_ (.A(_13585_),
    .B(_13959_),
    .Y(_13960_));
 sky130_fd_sc_hd__nand3_2 _36005_ (.A(_13960_),
    .B(_13663_),
    .C(_13664_),
    .Y(_13961_));
 sky130_fd_sc_hd__o211ai_2 _36006_ (.A1(_13585_),
    .A2(_13959_),
    .B1(_13669_),
    .C1(_13667_),
    .Y(_13962_));
 sky130_fd_sc_hd__nand2_2 _36007_ (.A(_13669_),
    .B(_13661_),
    .Y(_13963_));
 sky130_fd_sc_hd__a21o_2 _36008_ (.A1(_13961_),
    .A2(_13962_),
    .B1(_13963_),
    .X(_13964_));
 sky130_fd_sc_hd__buf_1 _36009_ (.A(_13963_),
    .X(_13965_));
 sky130_fd_sc_hd__nand3_2 _36010_ (.A(_13961_),
    .B(_13962_),
    .C(_13965_),
    .Y(_13966_));
 sky130_fd_sc_hd__nand2_2 _36011_ (.A(_13964_),
    .B(_13966_),
    .Y(_13967_));
 sky130_fd_sc_hd__o21a_2 _36012_ (.A1(_13620_),
    .A2(_13579_),
    .B1(_13595_),
    .X(_13968_));
 sky130_fd_sc_hd__nand2_2 _36013_ (.A(_13967_),
    .B(_13968_),
    .Y(_13969_));
 sky130_fd_sc_hd__o21ai_2 _36014_ (.A1(_13620_),
    .A2(_13579_),
    .B1(_13595_),
    .Y(_13970_));
 sky130_fd_sc_hd__nand3_2 _36015_ (.A(_13970_),
    .B(_13966_),
    .C(_13964_),
    .Y(_13971_));
 sky130_fd_sc_hd__o31ai_2 _36016_ (.A1(_13361_),
    .A2(_13671_),
    .A3(_13678_),
    .B1(_13670_),
    .Y(_13972_));
 sky130_fd_sc_hd__a21oi_2 _36017_ (.A1(_13969_),
    .A2(_13971_),
    .B1(_13972_),
    .Y(_13973_));
 sky130_fd_sc_hd__nand3_2 _36018_ (.A(_13969_),
    .B(_13972_),
    .C(_13971_),
    .Y(_13974_));
 sky130_fd_sc_hd__inv_2 _36019_ (.A(_13974_),
    .Y(_13975_));
 sky130_fd_sc_hd__a21oi_2 _36020_ (.A1(_13683_),
    .A2(_13681_),
    .B1(_13680_),
    .Y(_13976_));
 sky130_fd_sc_hd__o21ai_2 _36021_ (.A1(_13973_),
    .A2(_13975_),
    .B1(_13976_),
    .Y(_13977_));
 sky130_fd_sc_hd__nand2_2 _36022_ (.A(_13685_),
    .B(_13684_),
    .Y(_13978_));
 sky130_fd_sc_hd__a21o_2 _36023_ (.A1(_13969_),
    .A2(_13971_),
    .B1(_13972_),
    .X(_13979_));
 sky130_fd_sc_hd__nand3_2 _36024_ (.A(_13978_),
    .B(_13979_),
    .C(_13974_),
    .Y(_13980_));
 sky130_fd_sc_hd__nand3_2 _36025_ (.A(_13977_),
    .B(_13405_),
    .C(_13980_),
    .Y(_13981_));
 sky130_fd_sc_hd__a21oi_2 _36026_ (.A1(_13979_),
    .A2(_13974_),
    .B1(_13978_),
    .Y(_13982_));
 sky130_fd_sc_hd__nor3_2 _36027_ (.A(_13973_),
    .B(_13976_),
    .C(_13975_),
    .Y(_13983_));
 sky130_fd_sc_hd__o21ai_2 _36028_ (.A1(_13982_),
    .A2(_13983_),
    .B1(_13702_),
    .Y(_13984_));
 sky130_fd_sc_hd__o2111ai_2 _36029_ (.A1(_13646_),
    .A2(_13645_),
    .B1(_13635_),
    .C1(_13981_),
    .D1(_13984_),
    .Y(_13985_));
 sky130_fd_sc_hd__o21ai_2 _36030_ (.A1(_13982_),
    .A2(_13983_),
    .B1(_13406_),
    .Y(_13986_));
 sky130_fd_sc_hd__o21ai_2 _36031_ (.A1(_13645_),
    .A2(_13646_),
    .B1(_13632_),
    .Y(_13987_));
 sky130_fd_sc_hd__nand3_2 _36032_ (.A(_13977_),
    .B(_13397_),
    .C(_13980_),
    .Y(_13988_));
 sky130_fd_sc_hd__nand3_2 _36033_ (.A(_13986_),
    .B(_13987_),
    .C(_13988_),
    .Y(_13989_));
 sky130_fd_sc_hd__nor2_2 _36034_ (.A(_13405_),
    .B(_13688_),
    .Y(_13990_));
 sky130_fd_sc_hd__or2_2 _36035_ (.A(_13690_),
    .B(_13990_),
    .X(_13991_));
 sky130_fd_sc_hd__a21oi_2 _36036_ (.A1(_13985_),
    .A2(_13989_),
    .B1(_13991_),
    .Y(_13992_));
 sky130_fd_sc_hd__o211a_2 _36037_ (.A1(_13690_),
    .A2(_13990_),
    .B1(_13989_),
    .C1(_13985_),
    .X(_13993_));
 sky130_fd_sc_hd__o2bb2ai_2 _36038_ (.A1_N(_13950_),
    .A2_N(_13958_),
    .B1(_13992_),
    .B2(_13993_),
    .Y(_13994_));
 sky130_fd_sc_hd__nor2_2 _36039_ (.A(_13992_),
    .B(_13993_),
    .Y(_13995_));
 sky130_fd_sc_hd__nand3_2 _36040_ (.A(_13995_),
    .B(_13958_),
    .C(_13950_),
    .Y(_13996_));
 sky130_fd_sc_hd__nand2_2 _36041_ (.A(_13657_),
    .B(_13709_),
    .Y(_13997_));
 sky130_fd_sc_hd__nand2_2 _36042_ (.A(_13997_),
    .B(_13651_),
    .Y(_13998_));
 sky130_fd_sc_hd__a21oi_2 _36043_ (.A1(_13994_),
    .A2(_13996_),
    .B1(_13998_),
    .Y(_13999_));
 sky130_fd_sc_hd__and3_2 _36044_ (.A(_13638_),
    .B(_13640_),
    .C(_13650_),
    .X(_14000_));
 sky130_fd_sc_hd__a31oi_2 _36045_ (.A1(_13655_),
    .A2(_13654_),
    .A3(_13656_),
    .B1(_13715_),
    .Y(_14001_));
 sky130_fd_sc_hd__o211a_2 _36046_ (.A1(_14000_),
    .A2(_14001_),
    .B1(_13996_),
    .C1(_13994_),
    .X(_14002_));
 sky130_fd_sc_hd__o22ai_2 _36047_ (.A1(_13772_),
    .A2(_13773_),
    .B1(_13999_),
    .B2(_14002_),
    .Y(_14003_));
 sky130_fd_sc_hd__nand2_2 _36048_ (.A(_13718_),
    .B(_13732_),
    .Y(_14004_));
 sky130_fd_sc_hd__nand2_2 _36049_ (.A(_14004_),
    .B(_13723_),
    .Y(_14005_));
 sky130_fd_sc_hd__a21o_2 _36050_ (.A1(_13994_),
    .A2(_13996_),
    .B1(_13998_),
    .X(_14006_));
 sky130_fd_sc_hd__nand3_2 _36051_ (.A(_13998_),
    .B(_13994_),
    .C(_13996_),
    .Y(_14007_));
 sky130_fd_sc_hd__nor2_2 _36052_ (.A(_13773_),
    .B(_13772_),
    .Y(_14008_));
 sky130_fd_sc_hd__nand3_2 _36053_ (.A(_14006_),
    .B(_14007_),
    .C(_14008_),
    .Y(_14009_));
 sky130_fd_sc_hd__nand3_2 _36054_ (.A(_14003_),
    .B(_14005_),
    .C(_14009_),
    .Y(_14010_));
 sky130_fd_sc_hd__o21ai_2 _36055_ (.A1(_13999_),
    .A2(_14002_),
    .B1(_14008_),
    .Y(_14011_));
 sky130_fd_sc_hd__a21boi_2 _36056_ (.A1(_13718_),
    .A2(_13732_),
    .B1_N(_13723_),
    .Y(_14012_));
 sky130_fd_sc_hd__nor2_2 _36057_ (.A(_13736_),
    .B(_13708_),
    .Y(_14013_));
 sky130_fd_sc_hd__a21o_2 _36058_ (.A1(_13704_),
    .A2(_14013_),
    .B1(_13771_),
    .X(_14014_));
 sky130_fd_sc_hd__nand3_2 _36059_ (.A(_14006_),
    .B(_14007_),
    .C(_14014_),
    .Y(_14015_));
 sky130_fd_sc_hd__nand3_2 _36060_ (.A(_14011_),
    .B(_14012_),
    .C(_14015_),
    .Y(_14016_));
 sky130_fd_sc_hd__buf_1 _36061_ (.A(_13724_),
    .X(_14017_));
 sky130_fd_sc_hd__buf_1 _36062_ (.A(_14017_),
    .X(_14018_));
 sky130_fd_sc_hd__buf_1 _36063_ (.A(_14018_),
    .X(_14019_));
 sky130_fd_sc_hd__o2bb2ai_2 _36064_ (.A1_N(_14010_),
    .A2_N(_14016_),
    .B1(_14019_),
    .B2(_13726_),
    .Y(_14020_));
 sky130_fd_sc_hd__nand3_2 _36065_ (.A(_14016_),
    .B(_14010_),
    .C(_13727_),
    .Y(_14021_));
 sky130_fd_sc_hd__a21oi_2 _36066_ (.A1(_13740_),
    .A2(_13741_),
    .B1(_13742_),
    .Y(_14022_));
 sky130_fd_sc_hd__a21o_2 _36067_ (.A1(_13429_),
    .A2(_13743_),
    .B1(_14022_),
    .X(_14023_));
 sky130_fd_sc_hd__a21oi_2 _36068_ (.A1(_14020_),
    .A2(_14021_),
    .B1(_14023_),
    .Y(_14024_));
 sky130_fd_sc_hd__a21oi_2 _36069_ (.A1(_14016_),
    .A2(_14010_),
    .B1(_13727_),
    .Y(_14025_));
 sky130_fd_sc_hd__a31oi_2 _36070_ (.A1(_13740_),
    .A2(_13742_),
    .A3(_13741_),
    .B1(_13744_),
    .Y(_14026_));
 sky130_fd_sc_hd__o21ai_2 _36071_ (.A1(_14022_),
    .A2(_14026_),
    .B1(_14021_),
    .Y(_14027_));
 sky130_fd_sc_hd__nor2_2 _36072_ (.A(_14025_),
    .B(_14027_),
    .Y(_14028_));
 sky130_fd_sc_hd__nor2_2 _36073_ (.A(_14024_),
    .B(_14028_),
    .Y(_14029_));
 sky130_fd_sc_hd__nand2_2 _36074_ (.A(_13767_),
    .B(_13753_),
    .Y(_14030_));
 sky130_fd_sc_hd__xor2_2 _36075_ (.A(_14029_),
    .B(_14030_),
    .X(_02660_));
 sky130_fd_sc_hd__o21ai_2 _36076_ (.A1(_14014_),
    .A2(_13999_),
    .B1(_14007_),
    .Y(_14031_));
 sky130_fd_sc_hd__and3_2 _36077_ (.A(_11169_),
    .B(_13146_),
    .C(_06540_),
    .X(_14032_));
 sky130_fd_sc_hd__nand2_2 _36078_ (.A(_14032_),
    .B(_09012_),
    .Y(_14033_));
 sky130_fd_sc_hd__a22o_2 _36079_ (.A1(_10700_),
    .A2(_06074_),
    .B1(_09012_),
    .B2(_11122_),
    .X(_14034_));
 sky130_fd_sc_hd__buf_1 _36080_ (.A(_06391_),
    .X(_14035_));
 sky130_fd_sc_hd__o2bb2ai_2 _36081_ (.A1_N(_14033_),
    .A2_N(_14034_),
    .B1(_10151_),
    .B2(_14035_),
    .Y(_14036_));
 sky130_fd_sc_hd__nand2_2 _36082_ (.A(_10827_),
    .B(_19604_),
    .Y(_14037_));
 sky130_fd_sc_hd__nand3b_2 _36083_ (.A_N(_14037_),
    .B(_14034_),
    .C(_14033_),
    .Y(_14038_));
 sky130_fd_sc_hd__nand2_2 _36084_ (.A(_13845_),
    .B(_13841_),
    .Y(_14039_));
 sky130_fd_sc_hd__a21oi_2 _36085_ (.A1(_14036_),
    .A2(_14038_),
    .B1(_14039_),
    .Y(_14040_));
 sky130_fd_sc_hd__and3_2 _36086_ (.A(_14036_),
    .B(_14039_),
    .C(_14038_),
    .X(_14041_));
 sky130_fd_sc_hd__buf_1 _36087_ (.A(_10136_),
    .X(_14042_));
 sky130_fd_sc_hd__and4_2 _36088_ (.A(_10139_),
    .B(_14042_),
    .C(_19598_),
    .D(_19601_),
    .X(_14043_));
 sky130_fd_sc_hd__a22o_2 _36089_ (.A1(_19316_),
    .A2(_06059_),
    .B1(_09838_),
    .B2(_19597_),
    .X(_14044_));
 sky130_fd_sc_hd__inv_2 _36090_ (.A(_14044_),
    .Y(_14045_));
 sky130_fd_sc_hd__nor2_2 _36091_ (.A(_14043_),
    .B(_14045_),
    .Y(_14046_));
 sky130_fd_sc_hd__nor2_2 _36092_ (.A(_09358_),
    .B(_06959_),
    .Y(_14047_));
 sky130_fd_sc_hd__nand2_2 _36093_ (.A(_14046_),
    .B(_14047_),
    .Y(_14048_));
 sky130_fd_sc_hd__inv_2 _36094_ (.A(_14047_),
    .Y(_14049_));
 sky130_fd_sc_hd__o21ai_2 _36095_ (.A1(_14043_),
    .A2(_14045_),
    .B1(_14049_),
    .Y(_14050_));
 sky130_fd_sc_hd__nand2_2 _36096_ (.A(_14048_),
    .B(_14050_),
    .Y(_14051_));
 sky130_fd_sc_hd__o21ai_2 _36097_ (.A1(_14040_),
    .A2(_14041_),
    .B1(_14051_),
    .Y(_14052_));
 sky130_fd_sc_hd__o21ai_2 _36098_ (.A1(_13847_),
    .A2(_13858_),
    .B1(_13854_),
    .Y(_14053_));
 sky130_fd_sc_hd__inv_2 _36099_ (.A(_14039_),
    .Y(_14054_));
 sky130_fd_sc_hd__nand2_2 _36100_ (.A(_14036_),
    .B(_14038_),
    .Y(_14055_));
 sky130_fd_sc_hd__nand2_2 _36101_ (.A(_14054_),
    .B(_14055_),
    .Y(_14056_));
 sky130_fd_sc_hd__nand3_2 _36102_ (.A(_14036_),
    .B(_14039_),
    .C(_14038_),
    .Y(_14057_));
 sky130_fd_sc_hd__nand2_2 _36103_ (.A(_14046_),
    .B(_14049_),
    .Y(_14058_));
 sky130_fd_sc_hd__o21ai_2 _36104_ (.A1(_14043_),
    .A2(_14045_),
    .B1(_14047_),
    .Y(_14059_));
 sky130_fd_sc_hd__nand2_2 _36105_ (.A(_14058_),
    .B(_14059_),
    .Y(_14060_));
 sky130_fd_sc_hd__nand3_2 _36106_ (.A(_14056_),
    .B(_14057_),
    .C(_14060_),
    .Y(_14061_));
 sky130_fd_sc_hd__nand3_2 _36107_ (.A(_14052_),
    .B(_14053_),
    .C(_14061_),
    .Y(_14062_));
 sky130_fd_sc_hd__o21ai_2 _36108_ (.A1(_14040_),
    .A2(_14041_),
    .B1(_14060_),
    .Y(_14063_));
 sky130_fd_sc_hd__o21a_2 _36109_ (.A1(_13847_),
    .A2(_13858_),
    .B1(_13854_),
    .X(_14064_));
 sky130_fd_sc_hd__nand3_2 _36110_ (.A(_14056_),
    .B(_14057_),
    .C(_14051_),
    .Y(_14065_));
 sky130_fd_sc_hd__nand3_2 _36111_ (.A(_14063_),
    .B(_14064_),
    .C(_14065_),
    .Y(_14066_));
 sky130_fd_sc_hd__nand2_2 _36112_ (.A(_11205_),
    .B(_19591_),
    .Y(_14067_));
 sky130_fd_sc_hd__buf_1 _36113_ (.A(_10156_),
    .X(_14068_));
 sky130_fd_sc_hd__nand2_2 _36114_ (.A(_14068_),
    .B(_19589_),
    .Y(_14069_));
 sky130_fd_sc_hd__nand2_2 _36115_ (.A(_14067_),
    .B(_14069_),
    .Y(_14070_));
 sky130_fd_sc_hd__or2_2 _36116_ (.A(_14067_),
    .B(_14069_),
    .X(_14071_));
 sky130_fd_sc_hd__o2bb2ai_2 _36117_ (.A1_N(_14070_),
    .A2_N(_14071_),
    .B1(_08424_),
    .B2(_08611_),
    .Y(_14072_));
 sky130_fd_sc_hd__nor2_2 _36118_ (.A(_08424_),
    .B(_08611_),
    .Y(_14073_));
 sky130_fd_sc_hd__nand3_2 _36119_ (.A(_14071_),
    .B(_14073_),
    .C(_14070_),
    .Y(_14074_));
 sky130_fd_sc_hd__a21o_2 _36120_ (.A1(_13855_),
    .A2(_13835_),
    .B1(_13832_),
    .X(_14075_));
 sky130_fd_sc_hd__a21o_2 _36121_ (.A1(_14072_),
    .A2(_14074_),
    .B1(_14075_),
    .X(_14076_));
 sky130_fd_sc_hd__nand3_2 _36122_ (.A(_14072_),
    .B(_14075_),
    .C(_14074_),
    .Y(_14077_));
 sky130_fd_sc_hd__a21oi_2 _36123_ (.A1(_13874_),
    .A2(_13875_),
    .B1(_13867_),
    .Y(_14078_));
 sky130_fd_sc_hd__a21boi_2 _36124_ (.A1(_14076_),
    .A2(_14077_),
    .B1_N(_14078_),
    .Y(_14079_));
 sky130_fd_sc_hd__nand2_2 _36125_ (.A(_14076_),
    .B(_14077_),
    .Y(_14080_));
 sky130_fd_sc_hd__nor2_2 _36126_ (.A(_14078_),
    .B(_14080_),
    .Y(_14081_));
 sky130_fd_sc_hd__o2bb2ai_2 _36127_ (.A1_N(_14062_),
    .A2_N(_14066_),
    .B1(_14079_),
    .B2(_14081_),
    .Y(_14082_));
 sky130_fd_sc_hd__nand2_2 _36128_ (.A(_13884_),
    .B(_13860_),
    .Y(_14083_));
 sky130_fd_sc_hd__nand2_2 _36129_ (.A(_14083_),
    .B(_13864_),
    .Y(_14084_));
 sky130_fd_sc_hd__a21oi_2 _36130_ (.A1(_14072_),
    .A2(_14074_),
    .B1(_14075_),
    .Y(_14085_));
 sky130_fd_sc_hd__nor2_2 _36131_ (.A(_14078_),
    .B(_14085_),
    .Y(_14086_));
 sky130_fd_sc_hd__a21oi_2 _36132_ (.A1(_14077_),
    .A2(_14086_),
    .B1(_14079_),
    .Y(_14087_));
 sky130_fd_sc_hd__nand3_2 _36133_ (.A(_14087_),
    .B(_14066_),
    .C(_14062_),
    .Y(_14088_));
 sky130_fd_sc_hd__nand3_2 _36134_ (.A(_14082_),
    .B(_14084_),
    .C(_14088_),
    .Y(_14089_));
 sky130_fd_sc_hd__nand2_2 _36135_ (.A(_14066_),
    .B(_14062_),
    .Y(_14090_));
 sky130_fd_sc_hd__nand2_2 _36136_ (.A(_14090_),
    .B(_14087_),
    .Y(_14091_));
 sky130_fd_sc_hd__a21boi_2 _36137_ (.A1(_13884_),
    .A2(_13860_),
    .B1_N(_13864_),
    .Y(_14092_));
 sky130_fd_sc_hd__o211ai_2 _36138_ (.A1(_14079_),
    .A2(_14081_),
    .B1(_14066_),
    .C1(_14062_),
    .Y(_14093_));
 sky130_fd_sc_hd__nand3_2 _36139_ (.A(_14091_),
    .B(_14092_),
    .C(_14093_),
    .Y(_14094_));
 sky130_fd_sc_hd__buf_1 _36140_ (.A(_19337_),
    .X(_14095_));
 sky130_fd_sc_hd__and4_2 _36141_ (.A(_14095_),
    .B(_10656_),
    .C(_19581_),
    .D(_07852_),
    .X(_14096_));
 sky130_fd_sc_hd__inv_2 _36142_ (.A(_19340_),
    .Y(_14097_));
 sky130_fd_sc_hd__nand2_2 _36143_ (.A(_14095_),
    .B(_07852_),
    .Y(_14098_));
 sky130_fd_sc_hd__o21a_2 _36144_ (.A1(_14097_),
    .A2(_09263_),
    .B1(_14098_),
    .X(_14099_));
 sky130_fd_sc_hd__nand2_2 _36145_ (.A(_19343_),
    .B(_19578_),
    .Y(_14100_));
 sky130_fd_sc_hd__o21ai_2 _36146_ (.A1(_14096_),
    .A2(_14099_),
    .B1(_14100_),
    .Y(_14101_));
 sky130_fd_sc_hd__a21o_2 _36147_ (.A1(_13903_),
    .A2(_13901_),
    .B1(_13900_),
    .X(_14102_));
 sky130_fd_sc_hd__o21ai_2 _36148_ (.A1(_14097_),
    .A2(_09263_),
    .B1(_14098_),
    .Y(_14103_));
 sky130_fd_sc_hd__inv_2 _36149_ (.A(_14100_),
    .Y(_14104_));
 sky130_fd_sc_hd__nand3b_2 _36150_ (.A_N(_14096_),
    .B(_14103_),
    .C(_14104_),
    .Y(_14105_));
 sky130_fd_sc_hd__nand3_2 _36151_ (.A(_14101_),
    .B(_14102_),
    .C(_14105_),
    .Y(_14106_));
 sky130_fd_sc_hd__o21ai_2 _36152_ (.A1(_14096_),
    .A2(_14099_),
    .B1(_14104_),
    .Y(_14107_));
 sky130_fd_sc_hd__a21oi_2 _36153_ (.A1(_13903_),
    .A2(_13901_),
    .B1(_13900_),
    .Y(_14108_));
 sky130_fd_sc_hd__nand3b_2 _36154_ (.A_N(_14096_),
    .B(_14103_),
    .C(_14100_),
    .Y(_14109_));
 sky130_fd_sc_hd__nand3_2 _36155_ (.A(_14107_),
    .B(_14108_),
    .C(_14109_),
    .Y(_14110_));
 sky130_fd_sc_hd__and4_2 _36156_ (.A(_08808_),
    .B(_08185_),
    .C(_08496_),
    .D(_19574_),
    .X(_14111_));
 sky130_fd_sc_hd__buf_1 _36157_ (.A(_19570_),
    .X(_14112_));
 sky130_fd_sc_hd__a22o_2 _36158_ (.A1(_07481_),
    .A2(_09994_),
    .B1(_07907_),
    .B2(_14112_),
    .X(_14113_));
 sky130_fd_sc_hd__inv_2 _36159_ (.A(_14113_),
    .Y(_14114_));
 sky130_fd_sc_hd__nand2_2 _36160_ (.A(_19353_),
    .B(_19569_),
    .Y(_14115_));
 sky130_fd_sc_hd__o21bai_2 _36161_ (.A1(_14111_),
    .A2(_14114_),
    .B1_N(_14115_),
    .Y(_14116_));
 sky130_fd_sc_hd__nand3b_2 _36162_ (.A_N(_14111_),
    .B(_14115_),
    .C(_14113_),
    .Y(_14117_));
 sky130_fd_sc_hd__nand2_2 _36163_ (.A(_14116_),
    .B(_14117_),
    .Y(_14118_));
 sky130_fd_sc_hd__a21o_2 _36164_ (.A1(_14106_),
    .A2(_14110_),
    .B1(_14118_),
    .X(_14119_));
 sky130_fd_sc_hd__nand3_2 _36165_ (.A(_14118_),
    .B(_14106_),
    .C(_14110_),
    .Y(_14120_));
 sky130_fd_sc_hd__nand2_2 _36166_ (.A(_13887_),
    .B(_13877_),
    .Y(_14121_));
 sky130_fd_sc_hd__a21o_2 _36167_ (.A1(_14119_),
    .A2(_14120_),
    .B1(_14121_),
    .X(_14122_));
 sky130_fd_sc_hd__nand3_2 _36168_ (.A(_14121_),
    .B(_14119_),
    .C(_14120_),
    .Y(_14123_));
 sky130_fd_sc_hd__or2b_2 _36169_ (.A(_13921_),
    .B_N(_13907_),
    .X(_14124_));
 sky130_fd_sc_hd__and2_2 _36170_ (.A(_14124_),
    .B(_13911_),
    .X(_14125_));
 sky130_fd_sc_hd__a21oi_2 _36171_ (.A1(_14122_),
    .A2(_14123_),
    .B1(_14125_),
    .Y(_14126_));
 sky130_fd_sc_hd__inv_2 _36172_ (.A(_14123_),
    .Y(_14127_));
 sky130_fd_sc_hd__nand2_2 _36173_ (.A(_14122_),
    .B(_14125_),
    .Y(_14128_));
 sky130_fd_sc_hd__nor2_2 _36174_ (.A(_14127_),
    .B(_14128_),
    .Y(_14129_));
 sky130_fd_sc_hd__o2bb2ai_2 _36175_ (.A1_N(_14089_),
    .A2_N(_14094_),
    .B1(_14126_),
    .B2(_14129_),
    .Y(_14130_));
 sky130_fd_sc_hd__nand2_2 _36176_ (.A(_14124_),
    .B(_13911_),
    .Y(_14131_));
 sky130_fd_sc_hd__a21oi_2 _36177_ (.A1(_14119_),
    .A2(_14120_),
    .B1(_14121_),
    .Y(_14132_));
 sky130_fd_sc_hd__nor2_2 _36178_ (.A(_14131_),
    .B(_14132_),
    .Y(_14133_));
 sky130_fd_sc_hd__a21oi_2 _36179_ (.A1(_14123_),
    .A2(_14133_),
    .B1(_14126_),
    .Y(_14134_));
 sky130_fd_sc_hd__nand3_2 _36180_ (.A(_14134_),
    .B(_14094_),
    .C(_14089_),
    .Y(_14135_));
 sky130_fd_sc_hd__nand2_2 _36181_ (.A(_13940_),
    .B(_13896_),
    .Y(_14136_));
 sky130_fd_sc_hd__a21oi_2 _36182_ (.A1(_14130_),
    .A2(_14135_),
    .B1(_14136_),
    .Y(_14137_));
 sky130_fd_sc_hd__and3_2 _36183_ (.A(_14082_),
    .B(_14084_),
    .C(_14088_),
    .X(_14138_));
 sky130_fd_sc_hd__nand2_2 _36184_ (.A(_14134_),
    .B(_14094_),
    .Y(_14139_));
 sky130_fd_sc_hd__o211a_2 _36185_ (.A1(_14138_),
    .A2(_14139_),
    .B1(_14136_),
    .C1(_14130_),
    .X(_14140_));
 sky130_fd_sc_hd__nand2_2 _36186_ (.A(_06271_),
    .B(_19553_),
    .Y(_14141_));
 sky130_fd_sc_hd__nand2_2 _36187_ (.A(_06115_),
    .B(_11765_),
    .Y(_14142_));
 sky130_fd_sc_hd__nor2_2 _36188_ (.A(_14141_),
    .B(_14142_),
    .Y(_14143_));
 sky130_fd_sc_hd__and2_2 _36189_ (.A(_14141_),
    .B(_14142_),
    .X(_14144_));
 sky130_fd_sc_hd__nor2_2 _36190_ (.A(_06121_),
    .B(_10535_),
    .Y(_14145_));
 sky130_fd_sc_hd__o21bai_2 _36191_ (.A1(_14143_),
    .A2(_14144_),
    .B1_N(_14145_),
    .Y(_14146_));
 sky130_fd_sc_hd__nand2_2 _36192_ (.A(_14141_),
    .B(_14142_),
    .Y(_14147_));
 sky130_fd_sc_hd__nand3b_2 _36193_ (.A_N(_14143_),
    .B(_14145_),
    .C(_14147_),
    .Y(_14148_));
 sky130_fd_sc_hd__a31o_2 _36194_ (.A1(_13802_),
    .A2(_19369_),
    .A3(_19550_),
    .B1(_13798_),
    .X(_14149_));
 sky130_fd_sc_hd__a21o_2 _36195_ (.A1(_14146_),
    .A2(_14148_),
    .B1(_14149_),
    .X(_14150_));
 sky130_fd_sc_hd__nand3_2 _36196_ (.A(_14146_),
    .B(_14149_),
    .C(_14148_),
    .Y(_14151_));
 sky130_fd_sc_hd__a22oi_2 _36197_ (.A1(_18157_),
    .A2(_19374_),
    .B1(_19371_),
    .B2(_19541_),
    .Y(_14152_));
 sky130_fd_sc_hd__buf_1 _36198_ (.A(_11759_),
    .X(_14153_));
 sky130_fd_sc_hd__and4_2 _36199_ (.A(_14153_),
    .B(_05801_),
    .C(_05803_),
    .D(_11901_),
    .X(_14154_));
 sky130_fd_sc_hd__nor2_2 _36200_ (.A(_14152_),
    .B(_14154_),
    .Y(_14155_));
 sky130_fd_sc_hd__xor2_2 _36201_ (.A(_13810_),
    .B(_14155_),
    .X(_14156_));
 sky130_fd_sc_hd__a21oi_2 _36202_ (.A1(_14150_),
    .A2(_14151_),
    .B1(_14156_),
    .Y(_14157_));
 sky130_fd_sc_hd__nand3_2 _36203_ (.A(_14156_),
    .B(_14150_),
    .C(_14151_),
    .Y(_14158_));
 sky130_fd_sc_hd__inv_2 _36204_ (.A(_14158_),
    .Y(_14159_));
 sky130_fd_sc_hd__nand2_2 _36205_ (.A(_06822_),
    .B(_19564_),
    .Y(_14160_));
 sky130_fd_sc_hd__nand2_2 _36206_ (.A(_06828_),
    .B(_08905_),
    .Y(_14161_));
 sky130_fd_sc_hd__and2_2 _36207_ (.A(_14160_),
    .B(_14161_),
    .X(_14162_));
 sky130_fd_sc_hd__nor2_2 _36208_ (.A(_11300_),
    .B(_13274_),
    .Y(_14163_));
 sky130_fd_sc_hd__or2_2 _36209_ (.A(_14160_),
    .B(_14161_),
    .X(_14164_));
 sky130_fd_sc_hd__nand3b_2 _36210_ (.A_N(_14162_),
    .B(_14163_),
    .C(_14164_),
    .Y(_14165_));
 sky130_fd_sc_hd__nor2_2 _36211_ (.A(_14160_),
    .B(_14161_),
    .Y(_14166_));
 sky130_fd_sc_hd__o21bai_2 _36212_ (.A1(_14166_),
    .A2(_14162_),
    .B1_N(_14163_),
    .Y(_14167_));
 sky130_fd_sc_hd__nand2_2 _36213_ (.A(_14165_),
    .B(_14167_),
    .Y(_14168_));
 sky130_fd_sc_hd__a31o_2 _36214_ (.A1(_13917_),
    .A2(_12069_),
    .A3(_19571_),
    .B1(_13914_),
    .X(_14169_));
 sky130_fd_sc_hd__inv_2 _36215_ (.A(_14169_),
    .Y(_14170_));
 sky130_fd_sc_hd__nand2_2 _36216_ (.A(_14168_),
    .B(_14170_),
    .Y(_14171_));
 sky130_fd_sc_hd__nand3_2 _36217_ (.A(_14165_),
    .B(_14167_),
    .C(_14169_),
    .Y(_14172_));
 sky130_fd_sc_hd__nand2_2 _36218_ (.A(_14171_),
    .B(_14172_),
    .Y(_14173_));
 sky130_fd_sc_hd__and2_2 _36219_ (.A(_13780_),
    .B(_13777_),
    .X(_14174_));
 sky130_fd_sc_hd__nand2_2 _36220_ (.A(_14173_),
    .B(_14174_),
    .Y(_14175_));
 sky130_fd_sc_hd__nand3b_2 _36221_ (.A_N(_14174_),
    .B(_14171_),
    .C(_14172_),
    .Y(_14176_));
 sky130_fd_sc_hd__nand2_2 _36222_ (.A(_13792_),
    .B(_13791_),
    .Y(_14177_));
 sky130_fd_sc_hd__a21oi_2 _36223_ (.A1(_14175_),
    .A2(_14176_),
    .B1(_14177_),
    .Y(_14178_));
 sky130_fd_sc_hd__and3_2 _36224_ (.A(_14175_),
    .B(_14177_),
    .C(_14176_),
    .X(_14179_));
 sky130_fd_sc_hd__o22ai_2 _36225_ (.A1(_14157_),
    .A2(_14159_),
    .B1(_14178_),
    .B2(_14179_),
    .Y(_14180_));
 sky130_fd_sc_hd__a21o_2 _36226_ (.A1(_14175_),
    .A2(_14176_),
    .B1(_14177_),
    .X(_14181_));
 sky130_fd_sc_hd__nand3_2 _36227_ (.A(_14175_),
    .B(_14177_),
    .C(_14176_),
    .Y(_14182_));
 sky130_fd_sc_hd__nor2_2 _36228_ (.A(_14157_),
    .B(_14159_),
    .Y(_14183_));
 sky130_fd_sc_hd__nand3_2 _36229_ (.A(_14181_),
    .B(_14182_),
    .C(_14183_),
    .Y(_14184_));
 sky130_fd_sc_hd__a21bo_2 _36230_ (.A1(_13924_),
    .A2(_13930_),
    .B1_N(_13927_),
    .X(_14185_));
 sky130_fd_sc_hd__nand3_2 _36231_ (.A(_14180_),
    .B(_14184_),
    .C(_14185_),
    .Y(_14186_));
 sky130_fd_sc_hd__o21ai_2 _36232_ (.A1(_14178_),
    .A2(_14179_),
    .B1(_14183_),
    .Y(_14187_));
 sky130_fd_sc_hd__a21boi_2 _36233_ (.A1(_13930_),
    .A2(_13924_),
    .B1_N(_13927_),
    .Y(_14188_));
 sky130_fd_sc_hd__or2b_2 _36234_ (.A(_14157_),
    .B_N(_14158_),
    .X(_14189_));
 sky130_fd_sc_hd__nand3_2 _36235_ (.A(_14181_),
    .B(_14182_),
    .C(_14189_),
    .Y(_14190_));
 sky130_fd_sc_hd__nand2_2 _36236_ (.A(_13819_),
    .B(_13817_),
    .Y(_14191_));
 sky130_fd_sc_hd__and2_2 _36237_ (.A(_14191_),
    .B(_13820_),
    .X(_14192_));
 sky130_fd_sc_hd__a31oi_2 _36238_ (.A1(_14187_),
    .A2(_14188_),
    .A3(_14190_),
    .B1(_14192_),
    .Y(_14193_));
 sky130_fd_sc_hd__nand3_2 _36239_ (.A(_14187_),
    .B(_14188_),
    .C(_14190_),
    .Y(_14194_));
 sky130_fd_sc_hd__nand2_2 _36240_ (.A(_14191_),
    .B(_13820_),
    .Y(_14195_));
 sky130_fd_sc_hd__a21oi_2 _36241_ (.A1(_14194_),
    .A2(_14186_),
    .B1(_14195_),
    .Y(_14196_));
 sky130_fd_sc_hd__a21oi_2 _36242_ (.A1(_14186_),
    .A2(_14193_),
    .B1(_14196_),
    .Y(_14197_));
 sky130_fd_sc_hd__o21ai_2 _36243_ (.A1(_14137_),
    .A2(_14140_),
    .B1(_14197_),
    .Y(_14198_));
 sky130_fd_sc_hd__a21oi_2 _36244_ (.A1(_13946_),
    .A2(_13948_),
    .B1(_13941_),
    .Y(_14199_));
 sky130_fd_sc_hd__a21o_2 _36245_ (.A1(_14130_),
    .A2(_14135_),
    .B1(_14136_),
    .X(_14200_));
 sky130_fd_sc_hd__nand3_2 _36246_ (.A(_14130_),
    .B(_14136_),
    .C(_14135_),
    .Y(_14201_));
 sky130_fd_sc_hd__a21o_2 _36247_ (.A1(_14194_),
    .A2(_14186_),
    .B1(_14195_),
    .X(_14202_));
 sky130_fd_sc_hd__nand2_2 _36248_ (.A(_14193_),
    .B(_14186_),
    .Y(_14203_));
 sky130_fd_sc_hd__nand2_2 _36249_ (.A(_14202_),
    .B(_14203_),
    .Y(_14204_));
 sky130_fd_sc_hd__nand3_2 _36250_ (.A(_14200_),
    .B(_14201_),
    .C(_14204_),
    .Y(_14205_));
 sky130_fd_sc_hd__nand3_2 _36251_ (.A(_14198_),
    .B(_14199_),
    .C(_14205_),
    .Y(_14206_));
 sky130_fd_sc_hd__o21ai_2 _36252_ (.A1(_14137_),
    .A2(_14140_),
    .B1(_14204_),
    .Y(_14207_));
 sky130_fd_sc_hd__o21ai_2 _36253_ (.A1(_13938_),
    .A2(_13956_),
    .B1(_13947_),
    .Y(_14208_));
 sky130_fd_sc_hd__nand3_2 _36254_ (.A(_14200_),
    .B(_14197_),
    .C(_14201_),
    .Y(_14209_));
 sky130_fd_sc_hd__nand3_2 _36255_ (.A(_14207_),
    .B(_14208_),
    .C(_14209_),
    .Y(_14210_));
 sky130_fd_sc_hd__nand2_2 _36256_ (.A(_14206_),
    .B(_14210_),
    .Y(_14211_));
 sky130_fd_sc_hd__nand2_2 _36257_ (.A(_13667_),
    .B(_13668_),
    .Y(_14212_));
 sky130_fd_sc_hd__nor2_2 _36258_ (.A(_13809_),
    .B(_13808_),
    .Y(_14213_));
 sky130_fd_sc_hd__nor2_2 _36259_ (.A(_13811_),
    .B(_14213_),
    .Y(_14214_));
 sky130_fd_sc_hd__nand2_2 _36260_ (.A(_14212_),
    .B(_14214_),
    .Y(_14215_));
 sky130_fd_sc_hd__o211ai_2 _36261_ (.A1(_13811_),
    .A2(_14213_),
    .B1(_13669_),
    .C1(_13667_),
    .Y(_14216_));
 sky130_fd_sc_hd__buf_1 _36262_ (.A(_13963_),
    .X(_14217_));
 sky130_fd_sc_hd__a21o_2 _36263_ (.A1(_14215_),
    .A2(_14216_),
    .B1(_14217_),
    .X(_14218_));
 sky130_fd_sc_hd__nand3_2 _36264_ (.A(_14215_),
    .B(_14216_),
    .C(_13965_),
    .Y(_14219_));
 sky130_fd_sc_hd__o21ai_2 _36265_ (.A1(_13813_),
    .A2(_13812_),
    .B1(_13806_),
    .Y(_14220_));
 sky130_fd_sc_hd__nand2_2 _36266_ (.A(_14220_),
    .B(_13807_),
    .Y(_14221_));
 sky130_fd_sc_hd__a21oi_2 _36267_ (.A1(_14218_),
    .A2(_14219_),
    .B1(_14221_),
    .Y(_14222_));
 sky130_fd_sc_hd__inv_2 _36268_ (.A(_13814_),
    .Y(_14223_));
 sky130_fd_sc_hd__a21boi_2 _36269_ (.A1(_14223_),
    .A2(_13806_),
    .B1_N(_13807_),
    .Y(_14224_));
 sky130_fd_sc_hd__nand2_2 _36270_ (.A(_14218_),
    .B(_14219_),
    .Y(_14225_));
 sky130_fd_sc_hd__nor2_2 _36271_ (.A(_14224_),
    .B(_14225_),
    .Y(_14226_));
 sky130_fd_sc_hd__inv_2 _36272_ (.A(_13962_),
    .Y(_14227_));
 sky130_fd_sc_hd__and2_2 _36273_ (.A(_13961_),
    .B(_13965_),
    .X(_14228_));
 sky130_fd_sc_hd__nor2_2 _36274_ (.A(_14227_),
    .B(_14228_),
    .Y(_14229_));
 sky130_fd_sc_hd__o21ai_2 _36275_ (.A1(_14222_),
    .A2(_14226_),
    .B1(_14229_),
    .Y(_14230_));
 sky130_fd_sc_hd__a21oi_2 _36276_ (.A1(_14215_),
    .A2(_14216_),
    .B1(_14217_),
    .Y(_14231_));
 sky130_fd_sc_hd__inv_2 _36277_ (.A(_14219_),
    .Y(_14232_));
 sky130_fd_sc_hd__o21ai_2 _36278_ (.A1(_14231_),
    .A2(_14232_),
    .B1(_14224_),
    .Y(_14233_));
 sky130_fd_sc_hd__nand3_2 _36279_ (.A(_14221_),
    .B(_14219_),
    .C(_14218_),
    .Y(_14234_));
 sky130_fd_sc_hd__inv_2 _36280_ (.A(_14229_),
    .Y(_14235_));
 sky130_fd_sc_hd__nand3_2 _36281_ (.A(_14233_),
    .B(_14234_),
    .C(_14235_),
    .Y(_14236_));
 sky130_fd_sc_hd__nand2_2 _36282_ (.A(_13974_),
    .B(_13971_),
    .Y(_14237_));
 sky130_fd_sc_hd__nand3_2 _36283_ (.A(_14230_),
    .B(_14236_),
    .C(_14237_),
    .Y(_14238_));
 sky130_fd_sc_hd__inv_2 _36284_ (.A(_14238_),
    .Y(_14239_));
 sky130_fd_sc_hd__a21oi_2 _36285_ (.A1(_14233_),
    .A2(_14234_),
    .B1(_14235_),
    .Y(_14240_));
 sky130_fd_sc_hd__o211a_2 _36286_ (.A1(_14227_),
    .A2(_14228_),
    .B1(_14234_),
    .C1(_14233_),
    .X(_14241_));
 sky130_fd_sc_hd__o21bai_2 _36287_ (.A1(_14240_),
    .A2(_14241_),
    .B1_N(_14237_),
    .Y(_14242_));
 sky130_fd_sc_hd__buf_1 _36288_ (.A(_14242_),
    .X(_14243_));
 sky130_fd_sc_hd__nand2_2 _36289_ (.A(_14243_),
    .B(_13398_),
    .Y(_14244_));
 sky130_fd_sc_hd__o21ai_2 _36290_ (.A1(_13943_),
    .A2(_13944_),
    .B1(_13824_),
    .Y(_14245_));
 sky130_fd_sc_hd__o2bb2ai_2 _36291_ (.A1_N(_14238_),
    .A2_N(_14243_),
    .B1(_13352_),
    .B2(_13354_),
    .Y(_14246_));
 sky130_fd_sc_hd__o211a_2 _36292_ (.A1(_14239_),
    .A2(_14244_),
    .B1(_14245_),
    .C1(_14246_),
    .X(_14247_));
 sky130_fd_sc_hd__buf_1 _36293_ (.A(_13702_),
    .X(_14248_));
 sky130_fd_sc_hd__a21oi_2 _36294_ (.A1(_14243_),
    .A2(_14238_),
    .B1(_14248_),
    .Y(_14249_));
 sky130_fd_sc_hd__and3_2 _36295_ (.A(_14242_),
    .B(_13398_),
    .C(_14238_),
    .X(_14250_));
 sky130_fd_sc_hd__o21bai_2 _36296_ (.A1(_14249_),
    .A2(_14250_),
    .B1_N(_14245_),
    .Y(_14251_));
 sky130_fd_sc_hd__nand2_2 _36297_ (.A(_13988_),
    .B(_13980_),
    .Y(_14252_));
 sky130_fd_sc_hd__nand2_2 _36298_ (.A(_14251_),
    .B(_14252_),
    .Y(_14253_));
 sky130_fd_sc_hd__nand3_2 _36299_ (.A(_14243_),
    .B(_13402_),
    .C(_14238_),
    .Y(_14254_));
 sky130_fd_sc_hd__a21oi_2 _36300_ (.A1(_14246_),
    .A2(_14254_),
    .B1(_14245_),
    .Y(_14255_));
 sky130_fd_sc_hd__o21bai_2 _36301_ (.A1(_14255_),
    .A2(_14247_),
    .B1_N(_14252_),
    .Y(_14256_));
 sky130_fd_sc_hd__o21ai_2 _36302_ (.A1(_14247_),
    .A2(_14253_),
    .B1(_14256_),
    .Y(_14257_));
 sky130_fd_sc_hd__nand2_2 _36303_ (.A(_14211_),
    .B(_14257_),
    .Y(_14258_));
 sky130_fd_sc_hd__nand2_2 _36304_ (.A(_13995_),
    .B(_13958_),
    .Y(_14259_));
 sky130_fd_sc_hd__nand2_2 _36305_ (.A(_14259_),
    .B(_13950_),
    .Y(_14260_));
 sky130_fd_sc_hd__o21a_2 _36306_ (.A1(_14247_),
    .A2(_14253_),
    .B1(_14256_),
    .X(_14261_));
 sky130_fd_sc_hd__nand3_2 _36307_ (.A(_14261_),
    .B(_14210_),
    .C(_14206_),
    .Y(_14262_));
 sky130_fd_sc_hd__nand3_2 _36308_ (.A(_14258_),
    .B(_14260_),
    .C(_14262_),
    .Y(_14263_));
 sky130_fd_sc_hd__nand2_2 _36309_ (.A(_14211_),
    .B(_14261_),
    .Y(_14264_));
 sky130_fd_sc_hd__a21boi_2 _36310_ (.A1(_13995_),
    .A2(_13958_),
    .B1_N(_13950_),
    .Y(_14265_));
 sky130_fd_sc_hd__nand3_2 _36311_ (.A(_14257_),
    .B(_14206_),
    .C(_14210_),
    .Y(_14266_));
 sky130_fd_sc_hd__nand3_2 _36312_ (.A(_14264_),
    .B(_14265_),
    .C(_14266_),
    .Y(_14267_));
 sky130_fd_sc_hd__nand2_2 _36313_ (.A(_14263_),
    .B(_14267_),
    .Y(_14268_));
 sky130_fd_sc_hd__nand3_2 _36314_ (.A(_13985_),
    .B(_13991_),
    .C(_13989_),
    .Y(_14269_));
 sky130_fd_sc_hd__nand2_2 _36315_ (.A(_14269_),
    .B(_13989_),
    .Y(_14270_));
 sky130_fd_sc_hd__nor2_2 _36316_ (.A(_13735_),
    .B(_14270_),
    .Y(_14271_));
 sky130_fd_sc_hd__inv_2 _36317_ (.A(_14270_),
    .Y(_14272_));
 sky130_fd_sc_hd__nor2_2 _36318_ (.A(_13725_),
    .B(_14272_),
    .Y(_14273_));
 sky130_fd_sc_hd__nor2_2 _36319_ (.A(_14271_),
    .B(_14273_),
    .Y(_14274_));
 sky130_fd_sc_hd__nand2_2 _36320_ (.A(_14268_),
    .B(_14274_),
    .Y(_14275_));
 sky130_fd_sc_hd__inv_2 _36321_ (.A(_14274_),
    .Y(_14276_));
 sky130_fd_sc_hd__nand3_2 _36322_ (.A(_14276_),
    .B(_14263_),
    .C(_14267_),
    .Y(_14277_));
 sky130_fd_sc_hd__nand3b_2 _36323_ (.A_N(_14031_),
    .B(_14275_),
    .C(_14277_),
    .Y(_14278_));
 sky130_fd_sc_hd__nand2_2 _36324_ (.A(_14268_),
    .B(_14276_),
    .Y(_14279_));
 sky130_fd_sc_hd__nand3_2 _36325_ (.A(_14263_),
    .B(_14267_),
    .C(_14274_),
    .Y(_14280_));
 sky130_fd_sc_hd__nand3_2 _36326_ (.A(_14279_),
    .B(_14280_),
    .C(_14031_),
    .Y(_14281_));
 sky130_fd_sc_hd__nand3_2 _36327_ (.A(_14278_),
    .B(_13772_),
    .C(_14281_),
    .Y(_14282_));
 sky130_fd_sc_hd__inv_2 _36328_ (.A(_14282_),
    .Y(_14283_));
 sky130_fd_sc_hd__inv_2 _36329_ (.A(_13772_),
    .Y(_14284_));
 sky130_fd_sc_hd__nand2_2 _36330_ (.A(_14278_),
    .B(_14281_),
    .Y(_14285_));
 sky130_fd_sc_hd__nand2_2 _36331_ (.A(_14003_),
    .B(_14009_),
    .Y(_14286_));
 sky130_fd_sc_hd__nor2_2 _36332_ (.A(_14012_),
    .B(_14286_),
    .Y(_14287_));
 sky130_fd_sc_hd__a21boi_2 _36333_ (.A1(_14286_),
    .A2(_14012_),
    .B1_N(_13727_),
    .Y(_14288_));
 sky130_fd_sc_hd__o2bb2ai_2 _36334_ (.A1_N(_14284_),
    .A2_N(_14285_),
    .B1(_14287_),
    .B2(_14288_),
    .Y(_14289_));
 sky130_fd_sc_hd__nand2_2 _36335_ (.A(_14285_),
    .B(_13772_),
    .Y(_14290_));
 sky130_fd_sc_hd__a21oi_2 _36336_ (.A1(_13727_),
    .A2(_14016_),
    .B1(_14287_),
    .Y(_14291_));
 sky130_fd_sc_hd__nand3_2 _36337_ (.A(_14278_),
    .B(_14284_),
    .C(_14281_),
    .Y(_14292_));
 sky130_fd_sc_hd__nand3_2 _36338_ (.A(_14290_),
    .B(_14291_),
    .C(_14292_),
    .Y(_14293_));
 sky130_fd_sc_hd__o21a_2 _36339_ (.A1(_14283_),
    .A2(_14289_),
    .B1(_14293_),
    .X(_14294_));
 sky130_fd_sc_hd__nor3_2 _36340_ (.A(_14024_),
    .B(_14028_),
    .C(_13754_),
    .Y(_14295_));
 sky130_fd_sc_hd__or2b_2 _36341_ (.A(_13766_),
    .B_N(_14295_),
    .X(_14296_));
 sky130_fd_sc_hd__nand3_2 _36342_ (.A(_14023_),
    .B(_14020_),
    .C(_14021_),
    .Y(_14297_));
 sky130_fd_sc_hd__a21o_2 _36343_ (.A1(_14297_),
    .A2(_13753_),
    .B1(_14024_),
    .X(_14298_));
 sky130_fd_sc_hd__nand2_2 _36344_ (.A(_14296_),
    .B(_14298_),
    .Y(_14299_));
 sky130_fd_sc_hd__nor2_2 _36345_ (.A(_14294_),
    .B(_14299_),
    .Y(_14300_));
 sky130_fd_sc_hd__and2_2 _36346_ (.A(_14299_),
    .B(_14294_),
    .X(_14301_));
 sky130_fd_sc_hd__nor2_2 _36347_ (.A(_14300_),
    .B(_14301_),
    .Y(_02661_));
 sky130_fd_sc_hd__nand2_2 _36348_ (.A(_14285_),
    .B(_14284_),
    .Y(_14302_));
 sky130_fd_sc_hd__nand3b_2 _36349_ (.A_N(_14291_),
    .B(_14282_),
    .C(_14302_),
    .Y(_14303_));
 sky130_fd_sc_hd__a21oi_2 _36350_ (.A1(_14103_),
    .A2(_14104_),
    .B1(_14096_),
    .Y(_14304_));
 sky130_fd_sc_hd__and4_2 _36351_ (.A(_14095_),
    .B(_10656_),
    .C(_07845_),
    .D(_07848_),
    .X(_14305_));
 sky130_fd_sc_hd__a22o_2 _36352_ (.A1(_10655_),
    .A2(_07848_),
    .B1(_13454_),
    .B2(_19578_),
    .X(_14306_));
 sky130_fd_sc_hd__inv_2 _36353_ (.A(_14306_),
    .Y(_14307_));
 sky130_fd_sc_hd__nand2_2 _36354_ (.A(_19343_),
    .B(_12349_),
    .Y(_14308_));
 sky130_fd_sc_hd__o21ai_2 _36355_ (.A1(_14305_),
    .A2(_14307_),
    .B1(_14308_),
    .Y(_14309_));
 sky130_fd_sc_hd__inv_2 _36356_ (.A(_14308_),
    .Y(_14310_));
 sky130_fd_sc_hd__nand3b_2 _36357_ (.A_N(_14305_),
    .B(_14306_),
    .C(_14310_),
    .Y(_14311_));
 sky130_fd_sc_hd__nand3b_2 _36358_ (.A_N(_14304_),
    .B(_14309_),
    .C(_14311_),
    .Y(_14312_));
 sky130_fd_sc_hd__o21ai_2 _36359_ (.A1(_14305_),
    .A2(_14307_),
    .B1(_14310_),
    .Y(_14313_));
 sky130_fd_sc_hd__nand3b_2 _36360_ (.A_N(_14305_),
    .B(_14306_),
    .C(_14308_),
    .Y(_14314_));
 sky130_fd_sc_hd__nand3_2 _36361_ (.A(_14313_),
    .B(_14304_),
    .C(_14314_),
    .Y(_14315_));
 sky130_fd_sc_hd__and4_2 _36362_ (.A(_08808_),
    .B(_08185_),
    .C(_08664_),
    .D(_08496_),
    .X(_14316_));
 sky130_fd_sc_hd__o22a_2 _36363_ (.A1(_12596_),
    .A2(_12090_),
    .B1(_12597_),
    .B2(_09226_),
    .X(_14317_));
 sky130_fd_sc_hd__nor2_2 _36364_ (.A(_11251_),
    .B(_11671_),
    .Y(_14318_));
 sky130_fd_sc_hd__o21ai_2 _36365_ (.A1(_14316_),
    .A2(_14317_),
    .B1(_14318_),
    .Y(_14319_));
 sky130_fd_sc_hd__inv_2 _36366_ (.A(_14318_),
    .Y(_14320_));
 sky130_fd_sc_hd__a22o_2 _36367_ (.A1(_10210_),
    .A2(_14112_),
    .B1(_07907_),
    .B2(_08922_),
    .X(_14321_));
 sky130_fd_sc_hd__nand3b_2 _36368_ (.A_N(_14316_),
    .B(_14320_),
    .C(_14321_),
    .Y(_14322_));
 sky130_fd_sc_hd__nand2_2 _36369_ (.A(_14319_),
    .B(_14322_),
    .Y(_14323_));
 sky130_fd_sc_hd__a21o_2 _36370_ (.A1(_14312_),
    .A2(_14315_),
    .B1(_14323_),
    .X(_14324_));
 sky130_fd_sc_hd__nand3_2 _36371_ (.A(_14312_),
    .B(_14315_),
    .C(_14323_),
    .Y(_14325_));
 sky130_fd_sc_hd__o21ai_2 _36372_ (.A1(_14078_),
    .A2(_14085_),
    .B1(_14077_),
    .Y(_14326_));
 sky130_fd_sc_hd__a21o_2 _36373_ (.A1(_14324_),
    .A2(_14325_),
    .B1(_14326_),
    .X(_14327_));
 sky130_fd_sc_hd__nand3_2 _36374_ (.A(_14324_),
    .B(_14326_),
    .C(_14325_),
    .Y(_14328_));
 sky130_fd_sc_hd__inv_2 _36375_ (.A(_14106_),
    .Y(_14329_));
 sky130_fd_sc_hd__and2_2 _36376_ (.A(_14118_),
    .B(_14110_),
    .X(_14330_));
 sky130_fd_sc_hd__or2_2 _36377_ (.A(_14329_),
    .B(_14330_),
    .X(_14331_));
 sky130_fd_sc_hd__a21oi_2 _36378_ (.A1(_14327_),
    .A2(_14328_),
    .B1(_14331_),
    .Y(_14332_));
 sky130_fd_sc_hd__and3_2 _36379_ (.A(_14327_),
    .B(_14328_),
    .C(_14331_),
    .X(_14333_));
 sky130_fd_sc_hd__nand2_2 _36380_ (.A(_19329_),
    .B(_19589_),
    .Y(_14334_));
 sky130_fd_sc_hd__a21o_2 _36381_ (.A1(_19332_),
    .A2(_19586_),
    .B1(_14334_),
    .X(_14335_));
 sky130_fd_sc_hd__nand2_2 _36382_ (.A(_14068_),
    .B(_08959_),
    .Y(_14336_));
 sky130_fd_sc_hd__a21o_2 _36383_ (.A1(_19329_),
    .A2(_19589_),
    .B1(_14336_),
    .X(_14337_));
 sky130_fd_sc_hd__nand2_2 _36384_ (.A(_14335_),
    .B(_14337_),
    .Y(_14338_));
 sky130_fd_sc_hd__buf_1 _36385_ (.A(_08423_),
    .X(_14339_));
 sky130_fd_sc_hd__nor2_2 _36386_ (.A(_14339_),
    .B(_08957_),
    .Y(_14340_));
 sky130_fd_sc_hd__nand2_2 _36387_ (.A(_14338_),
    .B(_14340_),
    .Y(_14341_));
 sky130_fd_sc_hd__nand3b_2 _36388_ (.A_N(_14340_),
    .B(_14335_),
    .C(_14337_),
    .Y(_14342_));
 sky130_fd_sc_hd__a21o_2 _36389_ (.A1(_14047_),
    .A2(_14044_),
    .B1(_14043_),
    .X(_14343_));
 sky130_fd_sc_hd__a21o_2 _36390_ (.A1(_14341_),
    .A2(_14342_),
    .B1(_14343_),
    .X(_14344_));
 sky130_fd_sc_hd__nand3_2 _36391_ (.A(_14341_),
    .B(_14343_),
    .C(_14342_),
    .Y(_14345_));
 sky130_fd_sc_hd__nand2_2 _36392_ (.A(_14074_),
    .B(_14071_),
    .Y(_14346_));
 sky130_fd_sc_hd__and3_2 _36393_ (.A(_14344_),
    .B(_14345_),
    .C(_14346_),
    .X(_14347_));
 sky130_fd_sc_hd__a21oi_2 _36394_ (.A1(_14344_),
    .A2(_14345_),
    .B1(_14346_),
    .Y(_14348_));
 sky130_fd_sc_hd__buf_1 _36395_ (.A(_07313_),
    .X(_14349_));
 sky130_fd_sc_hd__buf_1 _36396_ (.A(_10824_),
    .X(_14350_));
 sky130_fd_sc_hd__buf_1 _36397_ (.A(_10823_),
    .X(_14351_));
 sky130_fd_sc_hd__and4_2 _36398_ (.A(_06225_),
    .B(_14350_),
    .C(_14351_),
    .D(_19604_),
    .X(_14352_));
 sky130_fd_sc_hd__buf_1 _36399_ (.A(_11164_),
    .X(_14353_));
 sky130_fd_sc_hd__o22a_2 _36400_ (.A1(_19607_),
    .A2(_18183_),
    .B1(_14353_),
    .B2(_14035_),
    .X(_14354_));
 sky130_fd_sc_hd__o22ai_2 _36401_ (.A1(_10152_),
    .A2(_14349_),
    .B1(_14352_),
    .B2(_14354_),
    .Y(_14355_));
 sky130_fd_sc_hd__buf_1 _36402_ (.A(_11514_),
    .X(_14356_));
 sky130_fd_sc_hd__a22o_2 _36403_ (.A1(_10700_),
    .A2(_06073_),
    .B1(_06688_),
    .B2(_14356_),
    .X(_14357_));
 sky130_fd_sc_hd__and3_2 _36404_ (.A(_10818_),
    .B(_10699_),
    .C(_05897_),
    .X(_14358_));
 sky130_fd_sc_hd__nand2_2 _36405_ (.A(_14358_),
    .B(_06688_),
    .Y(_14359_));
 sky130_fd_sc_hd__nor2_2 _36406_ (.A(_10151_),
    .B(_14349_),
    .Y(_14360_));
 sky130_fd_sc_hd__nand3_2 _36407_ (.A(_14357_),
    .B(_14359_),
    .C(_14360_),
    .Y(_14361_));
 sky130_fd_sc_hd__o22a_2 _36408_ (.A1(_19610_),
    .A2(_13848_),
    .B1(_14353_),
    .B2(_06225_),
    .X(_14362_));
 sky130_fd_sc_hd__o21ai_2 _36409_ (.A1(_14037_),
    .A2(_14362_),
    .B1(_14033_),
    .Y(_14363_));
 sky130_fd_sc_hd__a21oi_2 _36410_ (.A1(_14355_),
    .A2(_14361_),
    .B1(_14363_),
    .Y(_14364_));
 sky130_fd_sc_hd__nand2_2 _36411_ (.A(_14359_),
    .B(_14360_),
    .Y(_14365_));
 sky130_fd_sc_hd__o211a_2 _36412_ (.A1(_14354_),
    .A2(_14365_),
    .B1(_14363_),
    .C1(_14355_),
    .X(_14366_));
 sky130_fd_sc_hd__nor2_2 _36413_ (.A(_09358_),
    .B(_10279_),
    .Y(_14367_));
 sky130_fd_sc_hd__nand3_2 _36414_ (.A(_10139_),
    .B(_19320_),
    .C(_06954_),
    .Y(_14368_));
 sky130_fd_sc_hd__nor2_2 _36415_ (.A(_06397_),
    .B(_14368_),
    .Y(_14369_));
 sky130_fd_sc_hd__inv_2 _36416_ (.A(_19315_),
    .Y(_14370_));
 sky130_fd_sc_hd__buf_1 _36417_ (.A(_14370_),
    .X(_14371_));
 sky130_fd_sc_hd__nand2_2 _36418_ (.A(_14042_),
    .B(_19595_),
    .Y(_14372_));
 sky130_fd_sc_hd__o21a_2 _36419_ (.A1(_14371_),
    .A2(_06397_),
    .B1(_14372_),
    .X(_14373_));
 sky130_fd_sc_hd__nor3_2 _36420_ (.A(_14367_),
    .B(_14369_),
    .C(_14373_),
    .Y(_14374_));
 sky130_fd_sc_hd__o21a_2 _36421_ (.A1(_14369_),
    .A2(_14373_),
    .B1(_14367_),
    .X(_14375_));
 sky130_fd_sc_hd__nor2_2 _36422_ (.A(_14374_),
    .B(_14375_),
    .Y(_14376_));
 sky130_fd_sc_hd__o21ai_2 _36423_ (.A1(_14364_),
    .A2(_14366_),
    .B1(_14376_),
    .Y(_14377_));
 sky130_fd_sc_hd__a21o_2 _36424_ (.A1(_14355_),
    .A2(_14361_),
    .B1(_14363_),
    .X(_14378_));
 sky130_fd_sc_hd__nand3_2 _36425_ (.A(_14355_),
    .B(_14363_),
    .C(_14361_),
    .Y(_14379_));
 sky130_fd_sc_hd__nand3b_2 _36426_ (.A_N(_14376_),
    .B(_14378_),
    .C(_14379_),
    .Y(_14380_));
 sky130_fd_sc_hd__o21ai_2 _36427_ (.A1(_14040_),
    .A2(_14051_),
    .B1(_14057_),
    .Y(_14381_));
 sky130_fd_sc_hd__a21oi_2 _36428_ (.A1(_14377_),
    .A2(_14380_),
    .B1(_14381_),
    .Y(_14382_));
 sky130_fd_sc_hd__a22oi_2 _36429_ (.A1(_14058_),
    .A2(_14059_),
    .B1(_14054_),
    .B2(_14055_),
    .Y(_14383_));
 sky130_fd_sc_hd__o211a_2 _36430_ (.A1(_14041_),
    .A2(_14383_),
    .B1(_14380_),
    .C1(_14377_),
    .X(_14384_));
 sky130_fd_sc_hd__o22ai_2 _36431_ (.A1(_14347_),
    .A2(_14348_),
    .B1(_14382_),
    .B2(_14384_),
    .Y(_14385_));
 sky130_fd_sc_hd__nor2_2 _36432_ (.A(_14060_),
    .B(_14041_),
    .Y(_14386_));
 sky130_fd_sc_hd__o2bb2ai_2 _36433_ (.A1_N(_14377_),
    .A2_N(_14380_),
    .B1(_14040_),
    .B2(_14386_),
    .Y(_14387_));
 sky130_fd_sc_hd__nand3_2 _36434_ (.A(_14381_),
    .B(_14377_),
    .C(_14380_),
    .Y(_14388_));
 sky130_fd_sc_hd__nor2_2 _36435_ (.A(_14348_),
    .B(_14347_),
    .Y(_14389_));
 sky130_fd_sc_hd__nand3_2 _36436_ (.A(_14387_),
    .B(_14388_),
    .C(_14389_),
    .Y(_14390_));
 sky130_fd_sc_hd__inv_2 _36437_ (.A(_14061_),
    .Y(_14391_));
 sky130_fd_sc_hd__nand2_2 _36438_ (.A(_14052_),
    .B(_14053_),
    .Y(_14392_));
 sky130_fd_sc_hd__o2bb2ai_2 _36439_ (.A1_N(_14066_),
    .A2_N(_14087_),
    .B1(_14391_),
    .B2(_14392_),
    .Y(_14393_));
 sky130_fd_sc_hd__a21oi_2 _36440_ (.A1(_14385_),
    .A2(_14390_),
    .B1(_14393_),
    .Y(_14394_));
 sky130_fd_sc_hd__nand2_2 _36441_ (.A(_14389_),
    .B(_14388_),
    .Y(_14395_));
 sky130_fd_sc_hd__o211a_2 _36442_ (.A1(_14382_),
    .A2(_14395_),
    .B1(_14393_),
    .C1(_14385_),
    .X(_14396_));
 sky130_fd_sc_hd__o22ai_2 _36443_ (.A1(_14332_),
    .A2(_14333_),
    .B1(_14394_),
    .B2(_14396_),
    .Y(_14397_));
 sky130_fd_sc_hd__nand2_2 _36444_ (.A(_14139_),
    .B(_14089_),
    .Y(_14398_));
 sky130_fd_sc_hd__a21o_2 _36445_ (.A1(_14385_),
    .A2(_14390_),
    .B1(_14393_),
    .X(_14399_));
 sky130_fd_sc_hd__nor2_2 _36446_ (.A(_14332_),
    .B(_14333_),
    .Y(_14400_));
 sky130_fd_sc_hd__nand3_2 _36447_ (.A(_14385_),
    .B(_14393_),
    .C(_14390_),
    .Y(_14401_));
 sky130_fd_sc_hd__nand3_2 _36448_ (.A(_14399_),
    .B(_14400_),
    .C(_14401_),
    .Y(_14402_));
 sky130_fd_sc_hd__nand3_2 _36449_ (.A(_14397_),
    .B(_14398_),
    .C(_14402_),
    .Y(_14403_));
 sky130_fd_sc_hd__o21ai_2 _36450_ (.A1(_14394_),
    .A2(_14396_),
    .B1(_14400_),
    .Y(_14404_));
 sky130_fd_sc_hd__a21oi_2 _36451_ (.A1(_14134_),
    .A2(_14094_),
    .B1(_14138_),
    .Y(_14405_));
 sky130_fd_sc_hd__nand2_2 _36452_ (.A(_14327_),
    .B(_14328_),
    .Y(_14406_));
 sky130_fd_sc_hd__nor2_2 _36453_ (.A(_14329_),
    .B(_14330_),
    .Y(_14407_));
 sky130_fd_sc_hd__nand2_2 _36454_ (.A(_14406_),
    .B(_14407_),
    .Y(_14408_));
 sky130_fd_sc_hd__nand3_2 _36455_ (.A(_14327_),
    .B(_14328_),
    .C(_14331_),
    .Y(_14409_));
 sky130_fd_sc_hd__nand2_2 _36456_ (.A(_14408_),
    .B(_14409_),
    .Y(_14410_));
 sky130_fd_sc_hd__nand3_2 _36457_ (.A(_14399_),
    .B(_14410_),
    .C(_14401_),
    .Y(_14411_));
 sky130_fd_sc_hd__nand3_2 _36458_ (.A(_14404_),
    .B(_14405_),
    .C(_14411_),
    .Y(_14412_));
 sky130_fd_sc_hd__nor2_2 _36459_ (.A(_06119_),
    .B(_10519_),
    .Y(_14413_));
 sky130_fd_sc_hd__nand2_2 _36460_ (.A(_06790_),
    .B(_11765_),
    .Y(_14414_));
 sky130_fd_sc_hd__a21o_2 _36461_ (.A1(_19366_),
    .A2(_11038_),
    .B1(_14414_),
    .X(_14415_));
 sky130_fd_sc_hd__nand2_2 _36462_ (.A(_08320_),
    .B(_10537_),
    .Y(_14416_));
 sky130_fd_sc_hd__a21o_2 _36463_ (.A1(_19364_),
    .A2(_10371_),
    .B1(_14416_),
    .X(_14417_));
 sky130_fd_sc_hd__nand3b_2 _36464_ (.A_N(_14413_),
    .B(_14415_),
    .C(_14417_),
    .Y(_14418_));
 sky130_fd_sc_hd__nor2_2 _36465_ (.A(_14414_),
    .B(_14416_),
    .Y(_14419_));
 sky130_fd_sc_hd__nand2_2 _36466_ (.A(_14414_),
    .B(_14416_),
    .Y(_14420_));
 sky130_fd_sc_hd__nand3b_2 _36467_ (.A_N(_14419_),
    .B(_14413_),
    .C(_14420_),
    .Y(_14421_));
 sky130_fd_sc_hd__a31o_2 _36468_ (.A1(_14147_),
    .A2(_19369_),
    .A3(_19546_),
    .B1(_14143_),
    .X(_14422_));
 sky130_fd_sc_hd__a21o_2 _36469_ (.A1(_14418_),
    .A2(_14421_),
    .B1(_14422_),
    .X(_14423_));
 sky130_fd_sc_hd__nand3_2 _36470_ (.A(_14422_),
    .B(_14418_),
    .C(_14421_),
    .Y(_14424_));
 sky130_fd_sc_hd__o21a_2 _36471_ (.A1(_06430_),
    .A2(_06432_),
    .B1(_11759_),
    .X(_14425_));
 sky130_fd_sc_hd__nand3_2 _36472_ (.A(_11023_),
    .B(_05800_),
    .C(_05802_),
    .Y(_14426_));
 sky130_fd_sc_hd__nand2_2 _36473_ (.A(_14425_),
    .B(_14426_),
    .Y(_14427_));
 sky130_fd_sc_hd__nand2_2 _36474_ (.A(_14427_),
    .B(_13809_),
    .Y(_14428_));
 sky130_fd_sc_hd__o21a_2 _36475_ (.A1(_05498_),
    .A2(_14427_),
    .B1(_14428_),
    .X(_14429_));
 sky130_fd_sc_hd__buf_1 _36476_ (.A(_14429_),
    .X(_14430_));
 sky130_fd_sc_hd__a21oi_2 _36477_ (.A1(_14423_),
    .A2(_14424_),
    .B1(_14430_),
    .Y(_14431_));
 sky130_fd_sc_hd__and3_2 _36478_ (.A(_14423_),
    .B(_14424_),
    .C(_14430_),
    .X(_14432_));
 sky130_fd_sc_hd__nand2_2 _36479_ (.A(_07898_),
    .B(_19561_),
    .Y(_14433_));
 sky130_fd_sc_hd__nand2_2 _36480_ (.A(_08345_),
    .B(_09203_),
    .Y(_14434_));
 sky130_fd_sc_hd__nor2_2 _36481_ (.A(_14433_),
    .B(_14434_),
    .Y(_14435_));
 sky130_fd_sc_hd__and2_2 _36482_ (.A(_14433_),
    .B(_14434_),
    .X(_14436_));
 sky130_fd_sc_hd__nor2_2 _36483_ (.A(_08352_),
    .B(_10542_),
    .Y(_14437_));
 sky130_fd_sc_hd__o21bai_2 _36484_ (.A1(_14435_),
    .A2(_14436_),
    .B1_N(_14437_),
    .Y(_14438_));
 sky130_fd_sc_hd__or2_2 _36485_ (.A(_14433_),
    .B(_14434_),
    .X(_14439_));
 sky130_fd_sc_hd__nand2_2 _36486_ (.A(_14433_),
    .B(_14434_),
    .Y(_14440_));
 sky130_fd_sc_hd__nand3_2 _36487_ (.A(_14439_),
    .B(_14437_),
    .C(_14440_),
    .Y(_14441_));
 sky130_fd_sc_hd__a31o_2 _36488_ (.A1(_14113_),
    .A2(_19353_),
    .A3(_09223_),
    .B1(_14111_),
    .X(_14442_));
 sky130_fd_sc_hd__a21oi_2 _36489_ (.A1(_14438_),
    .A2(_14441_),
    .B1(_14442_),
    .Y(_14443_));
 sky130_fd_sc_hd__and3_2 _36490_ (.A(_14442_),
    .B(_14438_),
    .C(_14441_),
    .X(_14444_));
 sky130_fd_sc_hd__nand2_2 _36491_ (.A(_14165_),
    .B(_14164_),
    .Y(_14445_));
 sky130_fd_sc_hd__o21bai_2 _36492_ (.A1(_14443_),
    .A2(_14444_),
    .B1_N(_14445_),
    .Y(_14446_));
 sky130_fd_sc_hd__a21o_2 _36493_ (.A1(_14438_),
    .A2(_14441_),
    .B1(_14442_),
    .X(_14447_));
 sky130_fd_sc_hd__nand3_2 _36494_ (.A(_14442_),
    .B(_14438_),
    .C(_14441_),
    .Y(_14448_));
 sky130_fd_sc_hd__nand3_2 _36495_ (.A(_14447_),
    .B(_14448_),
    .C(_14445_),
    .Y(_14449_));
 sky130_fd_sc_hd__a21oi_2 _36496_ (.A1(_14165_),
    .A2(_14167_),
    .B1(_14169_),
    .Y(_14450_));
 sky130_fd_sc_hd__o21ai_2 _36497_ (.A1(_14174_),
    .A2(_14450_),
    .B1(_14172_),
    .Y(_14451_));
 sky130_fd_sc_hd__a21oi_2 _36498_ (.A1(_14446_),
    .A2(_14449_),
    .B1(_14451_),
    .Y(_14452_));
 sky130_fd_sc_hd__nand2_2 _36499_ (.A(_14447_),
    .B(_14445_),
    .Y(_14453_));
 sky130_fd_sc_hd__o211a_2 _36500_ (.A1(_14444_),
    .A2(_14453_),
    .B1(_14451_),
    .C1(_14446_),
    .X(_14454_));
 sky130_fd_sc_hd__o22ai_2 _36501_ (.A1(_14431_),
    .A2(_14432_),
    .B1(_14452_),
    .B2(_14454_),
    .Y(_14455_));
 sky130_fd_sc_hd__a21o_2 _36502_ (.A1(_14446_),
    .A2(_14449_),
    .B1(_14451_),
    .X(_14456_));
 sky130_fd_sc_hd__nor2_2 _36503_ (.A(_14431_),
    .B(_14432_),
    .Y(_14457_));
 sky130_fd_sc_hd__nand3_2 _36504_ (.A(_14446_),
    .B(_14451_),
    .C(_14449_),
    .Y(_14458_));
 sky130_fd_sc_hd__nand3_2 _36505_ (.A(_14456_),
    .B(_14457_),
    .C(_14458_),
    .Y(_14459_));
 sky130_fd_sc_hd__nand2_2 _36506_ (.A(_14128_),
    .B(_14123_),
    .Y(_14460_));
 sky130_fd_sc_hd__a21o_2 _36507_ (.A1(_14455_),
    .A2(_14459_),
    .B1(_14460_),
    .X(_14461_));
 sky130_fd_sc_hd__nand3_2 _36508_ (.A(_14460_),
    .B(_14455_),
    .C(_14459_),
    .Y(_14462_));
 sky130_fd_sc_hd__a21oi_2 _36509_ (.A1(_14181_),
    .A2(_14183_),
    .B1(_14179_),
    .Y(_14463_));
 sky130_fd_sc_hd__inv_2 _36510_ (.A(_14463_),
    .Y(_14464_));
 sky130_fd_sc_hd__nand3_2 _36511_ (.A(_14461_),
    .B(_14462_),
    .C(_14464_),
    .Y(_14465_));
 sky130_fd_sc_hd__inv_2 _36512_ (.A(_14465_),
    .Y(_14466_));
 sky130_fd_sc_hd__a21oi_2 _36513_ (.A1(_14461_),
    .A2(_14462_),
    .B1(_14464_),
    .Y(_14467_));
 sky130_fd_sc_hd__o2bb2ai_2 _36514_ (.A1_N(_14403_),
    .A2_N(_14412_),
    .B1(_14466_),
    .B2(_14467_),
    .Y(_14468_));
 sky130_fd_sc_hd__o21ai_2 _36515_ (.A1(_14137_),
    .A2(_14204_),
    .B1(_14201_),
    .Y(_14469_));
 sky130_fd_sc_hd__a21oi_2 _36516_ (.A1(_14455_),
    .A2(_14459_),
    .B1(_14460_),
    .Y(_14470_));
 sky130_fd_sc_hd__nor2_2 _36517_ (.A(_14463_),
    .B(_14470_),
    .Y(_14471_));
 sky130_fd_sc_hd__a21oi_2 _36518_ (.A1(_14462_),
    .A2(_14471_),
    .B1(_14467_),
    .Y(_14472_));
 sky130_fd_sc_hd__nand3_2 _36519_ (.A(_14472_),
    .B(_14412_),
    .C(_14403_),
    .Y(_14473_));
 sky130_fd_sc_hd__nand3_2 _36520_ (.A(_14468_),
    .B(_14469_),
    .C(_14473_),
    .Y(_14474_));
 sky130_fd_sc_hd__o211a_2 _36521_ (.A1(_14127_),
    .A2(_14133_),
    .B1(_14459_),
    .C1(_14455_),
    .X(_14475_));
 sky130_fd_sc_hd__o21ai_2 _36522_ (.A1(_14470_),
    .A2(_14475_),
    .B1(_14463_),
    .Y(_14476_));
 sky130_fd_sc_hd__nand2_2 _36523_ (.A(_14476_),
    .B(_14465_),
    .Y(_14477_));
 sky130_fd_sc_hd__a21o_2 _36524_ (.A1(_14412_),
    .A2(_14403_),
    .B1(_14477_),
    .X(_14478_));
 sky130_fd_sc_hd__a21oi_2 _36525_ (.A1(_14200_),
    .A2(_14197_),
    .B1(_14140_),
    .Y(_14479_));
 sky130_fd_sc_hd__nand3_2 _36526_ (.A(_14412_),
    .B(_14403_),
    .C(_14477_),
    .Y(_14480_));
 sky130_fd_sc_hd__nand3_2 _36527_ (.A(_14478_),
    .B(_14479_),
    .C(_14480_),
    .Y(_14481_));
 sky130_fd_sc_hd__buf_1 _36528_ (.A(_13406_),
    .X(_14482_));
 sky130_fd_sc_hd__nand2_2 _36529_ (.A(_14238_),
    .B(_14482_),
    .Y(_14483_));
 sky130_fd_sc_hd__a22o_2 _36530_ (.A1(_11429_),
    .A2(_05808_),
    .B1(_19371_),
    .B2(_11427_),
    .X(_14484_));
 sky130_fd_sc_hd__a21oi_2 _36531_ (.A1(_14484_),
    .A2(_13810_),
    .B1(_14154_),
    .Y(_14485_));
 sky130_fd_sc_hd__nand2_2 _36532_ (.A(_14212_),
    .B(_14485_),
    .Y(_14486_));
 sky130_fd_sc_hd__nand3b_2 _36533_ (.A_N(_14485_),
    .B(_13667_),
    .C(_13669_),
    .Y(_14487_));
 sky130_fd_sc_hd__buf_1 _36534_ (.A(_14217_),
    .X(_14488_));
 sky130_fd_sc_hd__a21oi_2 _36535_ (.A1(_14486_),
    .A2(_14487_),
    .B1(_14488_),
    .Y(_14489_));
 sky130_fd_sc_hd__and3_2 _36536_ (.A(_14486_),
    .B(_14487_),
    .C(_14488_),
    .X(_14490_));
 sky130_fd_sc_hd__a21boi_2 _36537_ (.A1(_14156_),
    .A2(_14150_),
    .B1_N(_14151_),
    .Y(_14491_));
 sky130_fd_sc_hd__o21ai_2 _36538_ (.A1(_14489_),
    .A2(_14490_),
    .B1(_14491_),
    .Y(_14492_));
 sky130_fd_sc_hd__a21oi_2 _36539_ (.A1(_14146_),
    .A2(_14148_),
    .B1(_14149_),
    .Y(_14493_));
 sky130_fd_sc_hd__xor2_2 _36540_ (.A(_13809_),
    .B(_14155_),
    .X(_14494_));
 sky130_fd_sc_hd__o21ai_2 _36541_ (.A1(_14493_),
    .A2(_14494_),
    .B1(_14151_),
    .Y(_14495_));
 sky130_fd_sc_hd__nand3_2 _36542_ (.A(_14486_),
    .B(_14487_),
    .C(_14488_),
    .Y(_14496_));
 sky130_fd_sc_hd__a21o_2 _36543_ (.A1(_14486_),
    .A2(_14487_),
    .B1(_14488_),
    .X(_14497_));
 sky130_fd_sc_hd__nand3_2 _36544_ (.A(_14495_),
    .B(_14496_),
    .C(_14497_),
    .Y(_14498_));
 sky130_fd_sc_hd__inv_2 _36545_ (.A(_14216_),
    .Y(_14499_));
 sky130_fd_sc_hd__and2_2 _36546_ (.A(_14215_),
    .B(_14488_),
    .X(_14500_));
 sky130_fd_sc_hd__or2_2 _36547_ (.A(_14499_),
    .B(_14500_),
    .X(_14501_));
 sky130_fd_sc_hd__a21oi_2 _36548_ (.A1(_14492_),
    .A2(_14498_),
    .B1(_14501_),
    .Y(_14502_));
 sky130_fd_sc_hd__o211a_2 _36549_ (.A1(_14499_),
    .A2(_14500_),
    .B1(_14498_),
    .C1(_14492_),
    .X(_14503_));
 sky130_fd_sc_hd__a21oi_2 _36550_ (.A1(_14233_),
    .A2(_14235_),
    .B1(_14226_),
    .Y(_14504_));
 sky130_fd_sc_hd__o21ai_2 _36551_ (.A1(_14502_),
    .A2(_14503_),
    .B1(_14504_),
    .Y(_14505_));
 sky130_fd_sc_hd__a21o_2 _36552_ (.A1(_14492_),
    .A2(_14498_),
    .B1(_14501_),
    .X(_14506_));
 sky130_fd_sc_hd__nand3_2 _36553_ (.A(_14501_),
    .B(_14492_),
    .C(_14498_),
    .Y(_14507_));
 sky130_fd_sc_hd__o21ai_2 _36554_ (.A1(_14229_),
    .A2(_14222_),
    .B1(_14234_),
    .Y(_14508_));
 sky130_fd_sc_hd__nand3_2 _36555_ (.A(_14506_),
    .B(_14507_),
    .C(_14508_),
    .Y(_14509_));
 sky130_fd_sc_hd__a21oi_2 _36556_ (.A1(_14505_),
    .A2(_14509_),
    .B1(_14248_),
    .Y(_14510_));
 sky130_fd_sc_hd__nand2_2 _36557_ (.A(_14506_),
    .B(_14508_),
    .Y(_14511_));
 sky130_fd_sc_hd__o211a_2 _36558_ (.A1(_14503_),
    .A2(_14511_),
    .B1(_13402_),
    .C1(_14505_),
    .X(_14512_));
 sky130_fd_sc_hd__and3_2 _36559_ (.A(_14180_),
    .B(_14184_),
    .C(_14185_),
    .X(_14513_));
 sky130_fd_sc_hd__nor2_2 _36560_ (.A(_14513_),
    .B(_14193_),
    .Y(_14514_));
 sky130_fd_sc_hd__o21ai_2 _36561_ (.A1(_14510_),
    .A2(_14512_),
    .B1(_14514_),
    .Y(_14515_));
 sky130_fd_sc_hd__inv_2 _36562_ (.A(_14184_),
    .Y(_14516_));
 sky130_fd_sc_hd__nand2_2 _36563_ (.A(_14180_),
    .B(_14185_),
    .Y(_14517_));
 sky130_fd_sc_hd__o2bb2ai_2 _36564_ (.A1_N(_14194_),
    .A2_N(_14195_),
    .B1(_14516_),
    .B2(_14517_),
    .Y(_14518_));
 sky130_fd_sc_hd__nand3_2 _36565_ (.A(_14505_),
    .B(_13402_),
    .C(_14509_),
    .Y(_14519_));
 sky130_fd_sc_hd__o2bb2ai_2 _36566_ (.A1_N(_14509_),
    .A2_N(_14505_),
    .B1(_13352_),
    .B2(_13354_),
    .Y(_14520_));
 sky130_fd_sc_hd__nand3_2 _36567_ (.A(_14518_),
    .B(_14519_),
    .C(_14520_),
    .Y(_14521_));
 sky130_fd_sc_hd__a22oi_2 _36568_ (.A1(_14243_),
    .A2(_14483_),
    .B1(_14515_),
    .B2(_14521_),
    .Y(_14522_));
 sky130_fd_sc_hd__inv_2 _36569_ (.A(_14244_),
    .Y(_14523_));
 sky130_fd_sc_hd__o211a_2 _36570_ (.A1(_14239_),
    .A2(_14523_),
    .B1(_14521_),
    .C1(_14515_),
    .X(_14524_));
 sky130_fd_sc_hd__o2bb2ai_2 _36571_ (.A1_N(_14474_),
    .A2_N(_14481_),
    .B1(_14522_),
    .B2(_14524_),
    .Y(_14525_));
 sky130_fd_sc_hd__nor2_2 _36572_ (.A(_14522_),
    .B(_14524_),
    .Y(_14526_));
 sky130_fd_sc_hd__nand3_2 _36573_ (.A(_14526_),
    .B(_14481_),
    .C(_14474_),
    .Y(_14527_));
 sky130_fd_sc_hd__inv_2 _36574_ (.A(_14209_),
    .Y(_14528_));
 sky130_fd_sc_hd__nand2_2 _36575_ (.A(_14207_),
    .B(_14208_),
    .Y(_14529_));
 sky130_fd_sc_hd__a21oi_2 _36576_ (.A1(_14207_),
    .A2(_14209_),
    .B1(_14208_),
    .Y(_14530_));
 sky130_fd_sc_hd__o22ai_2 _36577_ (.A1(_14528_),
    .A2(_14529_),
    .B1(_14257_),
    .B2(_14530_),
    .Y(_14531_));
 sky130_fd_sc_hd__a21oi_2 _36578_ (.A1(_14525_),
    .A2(_14527_),
    .B1(_14531_),
    .Y(_14532_));
 sky130_fd_sc_hd__and3_2 _36579_ (.A(_14468_),
    .B(_14469_),
    .C(_14473_),
    .X(_14533_));
 sky130_fd_sc_hd__nand2_2 _36580_ (.A(_14526_),
    .B(_14481_),
    .Y(_14534_));
 sky130_fd_sc_hd__o211a_2 _36581_ (.A1(_14533_),
    .A2(_14534_),
    .B1(_14531_),
    .C1(_14525_),
    .X(_14535_));
 sky130_fd_sc_hd__nand2_2 _36582_ (.A(_14245_),
    .B(_14254_),
    .Y(_14536_));
 sky130_fd_sc_hd__o21ai_2 _36583_ (.A1(_14249_),
    .A2(_14536_),
    .B1(_14253_),
    .Y(_14537_));
 sky130_fd_sc_hd__nor2_2 _36584_ (.A(_13736_),
    .B(_14537_),
    .Y(_14538_));
 sky130_fd_sc_hd__nand2_2 _36585_ (.A(_14537_),
    .B(_13735_),
    .Y(_14539_));
 sky130_fd_sc_hd__inv_2 _36586_ (.A(_14539_),
    .Y(_14540_));
 sky130_fd_sc_hd__nor2_2 _36587_ (.A(_14538_),
    .B(_14540_),
    .Y(_14541_));
 sky130_fd_sc_hd__o21ai_2 _36588_ (.A1(_14532_),
    .A2(_14535_),
    .B1(_14541_),
    .Y(_14542_));
 sky130_fd_sc_hd__a21boi_2 _36589_ (.A1(_14267_),
    .A2(_14274_),
    .B1_N(_14263_),
    .Y(_14543_));
 sky130_fd_sc_hd__a21o_2 _36590_ (.A1(_14525_),
    .A2(_14527_),
    .B1(_14531_),
    .X(_14544_));
 sky130_fd_sc_hd__nand3_2 _36591_ (.A(_14525_),
    .B(_14531_),
    .C(_14527_),
    .Y(_14545_));
 sky130_fd_sc_hd__or2b_2 _36592_ (.A(_14538_),
    .B_N(_14539_),
    .X(_14546_));
 sky130_fd_sc_hd__nand3_2 _36593_ (.A(_14544_),
    .B(_14545_),
    .C(_14546_),
    .Y(_14547_));
 sky130_fd_sc_hd__nand3_2 _36594_ (.A(_14542_),
    .B(_14543_),
    .C(_14547_),
    .Y(_14548_));
 sky130_fd_sc_hd__buf_1 _36595_ (.A(_14540_),
    .X(_14549_));
 sky130_fd_sc_hd__o22ai_2 _36596_ (.A1(_14549_),
    .A2(_14538_),
    .B1(_14532_),
    .B2(_14535_),
    .Y(_14550_));
 sky130_fd_sc_hd__nand2_2 _36597_ (.A(_14267_),
    .B(_14274_),
    .Y(_14551_));
 sky130_fd_sc_hd__nand2_2 _36598_ (.A(_14551_),
    .B(_14263_),
    .Y(_14552_));
 sky130_fd_sc_hd__nand3_2 _36599_ (.A(_14544_),
    .B(_14541_),
    .C(_14545_),
    .Y(_14553_));
 sky130_fd_sc_hd__nand3_2 _36600_ (.A(_14550_),
    .B(_14552_),
    .C(_14553_),
    .Y(_14554_));
 sky130_fd_sc_hd__nand3_2 _36601_ (.A(_14548_),
    .B(_14554_),
    .C(_14273_),
    .Y(_14555_));
 sky130_fd_sc_hd__nand2_2 _36602_ (.A(_14278_),
    .B(_13772_),
    .Y(_14556_));
 sky130_fd_sc_hd__inv_2 _36603_ (.A(_14273_),
    .Y(_14557_));
 sky130_fd_sc_hd__nand2_2 _36604_ (.A(_14548_),
    .B(_14554_),
    .Y(_14558_));
 sky130_fd_sc_hd__a22oi_2 _36605_ (.A1(_14556_),
    .A2(_14281_),
    .B1(_14557_),
    .B2(_14558_),
    .Y(_14559_));
 sky130_fd_sc_hd__o2bb2ai_2 _36606_ (.A1_N(_14554_),
    .A2_N(_14548_),
    .B1(_14019_),
    .B2(_14272_),
    .Y(_14560_));
 sky130_fd_sc_hd__nand2_2 _36607_ (.A(_14556_),
    .B(_14281_),
    .Y(_14561_));
 sky130_fd_sc_hd__a21oi_2 _36608_ (.A1(_14560_),
    .A2(_14555_),
    .B1(_14561_),
    .Y(_14562_));
 sky130_fd_sc_hd__a21oi_2 _36609_ (.A1(_14555_),
    .A2(_14559_),
    .B1(_14562_),
    .Y(_14563_));
 sky130_fd_sc_hd__nand3b_2 _36610_ (.A_N(_14301_),
    .B(_14303_),
    .C(_14563_),
    .Y(_14564_));
 sky130_fd_sc_hd__nand2_2 _36611_ (.A(_14299_),
    .B(_14294_),
    .Y(_14565_));
 sky130_fd_sc_hd__a21o_2 _36612_ (.A1(_14565_),
    .A2(_14303_),
    .B1(_14563_),
    .X(_14566_));
 sky130_fd_sc_hd__nand2_2 _36613_ (.A(_14564_),
    .B(_14566_),
    .Y(_02662_));
 sky130_fd_sc_hd__o21ai_2 _36614_ (.A1(_14371_),
    .A2(_06397_),
    .B1(_14372_),
    .Y(_14567_));
 sky130_fd_sc_hd__a21oi_2 _36615_ (.A1(_14567_),
    .A2(_14367_),
    .B1(_14369_),
    .Y(_14568_));
 sky130_fd_sc_hd__buf_1 _36616_ (.A(_10166_),
    .X(_14569_));
 sky130_fd_sc_hd__and4_2 _36617_ (.A(_14569_),
    .B(_10867_),
    .C(_07852_),
    .D(_08959_),
    .X(_14570_));
 sky130_fd_sc_hd__inv_2 _36618_ (.A(_10166_),
    .Y(_14571_));
 sky130_fd_sc_hd__o22a_2 _36619_ (.A1(_14571_),
    .A2(_08611_),
    .B1(_13873_),
    .B2(_08957_),
    .X(_14572_));
 sky130_fd_sc_hd__nor2_2 _36620_ (.A(_14570_),
    .B(_14572_),
    .Y(_14573_));
 sky130_fd_sc_hd__nor2_2 _36621_ (.A(_14339_),
    .B(_09246_),
    .Y(_14574_));
 sky130_fd_sc_hd__nand2_2 _36622_ (.A(_14573_),
    .B(_14574_),
    .Y(_14575_));
 sky130_fd_sc_hd__inv_2 _36623_ (.A(_14574_),
    .Y(_14576_));
 sky130_fd_sc_hd__o21ai_2 _36624_ (.A1(_14570_),
    .A2(_14572_),
    .B1(_14576_),
    .Y(_14577_));
 sky130_fd_sc_hd__nand3b_2 _36625_ (.A_N(_14568_),
    .B(_14575_),
    .C(_14577_),
    .Y(_14578_));
 sky130_fd_sc_hd__nand2_2 _36626_ (.A(_14573_),
    .B(_14576_),
    .Y(_14579_));
 sky130_fd_sc_hd__o21ai_2 _36627_ (.A1(_14570_),
    .A2(_14572_),
    .B1(_14574_),
    .Y(_14580_));
 sky130_fd_sc_hd__nand3_2 _36628_ (.A(_14579_),
    .B(_14568_),
    .C(_14580_),
    .Y(_14581_));
 sky130_fd_sc_hd__nor2_2 _36629_ (.A(_14334_),
    .B(_14336_),
    .Y(_14582_));
 sky130_fd_sc_hd__a21oi_2 _36630_ (.A1(_14338_),
    .A2(_14340_),
    .B1(_14582_),
    .Y(_14583_));
 sky130_fd_sc_hd__inv_2 _36631_ (.A(_14583_),
    .Y(_14584_));
 sky130_fd_sc_hd__nand3_2 _36632_ (.A(_14578_),
    .B(_14581_),
    .C(_14584_),
    .Y(_14585_));
 sky130_fd_sc_hd__inv_2 _36633_ (.A(_14585_),
    .Y(_14586_));
 sky130_fd_sc_hd__a21oi_2 _36634_ (.A1(_14578_),
    .A2(_14581_),
    .B1(_14584_),
    .Y(_14587_));
 sky130_fd_sc_hd__o22a_2 _36635_ (.A1(_19604_),
    .A2(_13848_),
    .B1(_14353_),
    .B2(_14349_),
    .X(_14588_));
 sky130_fd_sc_hd__nand2_2 _36636_ (.A(_19312_),
    .B(_19598_),
    .Y(_14589_));
 sky130_fd_sc_hd__a41o_2 _36637_ (.A1(_14035_),
    .A2(_11123_),
    .A3(_19309_),
    .A4(_19601_),
    .B1(_14589_),
    .X(_14590_));
 sky130_fd_sc_hd__nor2_2 _36638_ (.A(_14588_),
    .B(_14590_),
    .Y(_14591_));
 sky130_fd_sc_hd__a22o_2 _36639_ (.A1(_19309_),
    .A2(_19601_),
    .B1(_14035_),
    .B2(_14350_),
    .X(_14592_));
 sky130_fd_sc_hd__and3_2 _36640_ (.A(_14356_),
    .B(_19308_),
    .C(_06222_),
    .X(_14593_));
 sky130_fd_sc_hd__nand2_2 _36641_ (.A(_14593_),
    .B(_14035_),
    .Y(_14594_));
 sky130_fd_sc_hd__inv_2 _36642_ (.A(_14589_),
    .Y(_14595_));
 sky130_fd_sc_hd__a21oi_2 _36643_ (.A1(_14592_),
    .A2(_14594_),
    .B1(_14595_),
    .Y(_14596_));
 sky130_fd_sc_hd__a21oi_2 _36644_ (.A1(_14357_),
    .A2(_14360_),
    .B1(_14352_),
    .Y(_14597_));
 sky130_fd_sc_hd__o21ai_2 _36645_ (.A1(_14591_),
    .A2(_14596_),
    .B1(_14597_),
    .Y(_14598_));
 sky130_fd_sc_hd__nand2_2 _36646_ (.A(_14361_),
    .B(_14359_),
    .Y(_14599_));
 sky130_fd_sc_hd__and4_2 _36647_ (.A(_14035_),
    .B(_11122_),
    .C(_10700_),
    .D(_19601_),
    .X(_14600_));
 sky130_fd_sc_hd__o21ai_2 _36648_ (.A1(_14600_),
    .A2(_14588_),
    .B1(_14589_),
    .Y(_14601_));
 sky130_fd_sc_hd__nand3_2 _36649_ (.A(_14592_),
    .B(_14594_),
    .C(_14595_),
    .Y(_14602_));
 sky130_fd_sc_hd__nand3_2 _36650_ (.A(_14599_),
    .B(_14601_),
    .C(_14602_),
    .Y(_14603_));
 sky130_fd_sc_hd__nand2_2 _36651_ (.A(_14598_),
    .B(_14603_),
    .Y(_14604_));
 sky130_fd_sc_hd__a22oi_2 _36652_ (.A1(_19317_),
    .A2(_19595_),
    .B1(_14042_),
    .B2(_19591_),
    .Y(_14605_));
 sky130_fd_sc_hd__nand2_2 _36653_ (.A(_19323_),
    .B(_07380_),
    .Y(_14606_));
 sky130_fd_sc_hd__inv_2 _36654_ (.A(_14606_),
    .Y(_14607_));
 sky130_fd_sc_hd__nor2_2 _36655_ (.A(_10279_),
    .B(_14368_),
    .Y(_14608_));
 sky130_fd_sc_hd__nor3_2 _36656_ (.A(_14605_),
    .B(_14607_),
    .C(_14608_),
    .Y(_14609_));
 sky130_fd_sc_hd__nor2_2 _36657_ (.A(_14605_),
    .B(_14608_),
    .Y(_14610_));
 sky130_fd_sc_hd__nor2_2 _36658_ (.A(_14606_),
    .B(_14610_),
    .Y(_14611_));
 sky130_fd_sc_hd__nor2_2 _36659_ (.A(_14609_),
    .B(_14611_),
    .Y(_14612_));
 sky130_fd_sc_hd__nand2_2 _36660_ (.A(_14604_),
    .B(_14612_),
    .Y(_14613_));
 sky130_fd_sc_hd__nand2_2 _36661_ (.A(_14610_),
    .B(_14606_),
    .Y(_14614_));
 sky130_fd_sc_hd__or2b_2 _36662_ (.A(_14611_),
    .B_N(_14614_),
    .X(_14615_));
 sky130_fd_sc_hd__nand3_2 _36663_ (.A(_14615_),
    .B(_14598_),
    .C(_14603_),
    .Y(_14616_));
 sky130_fd_sc_hd__o21ai_2 _36664_ (.A1(_14376_),
    .A2(_14364_),
    .B1(_14379_),
    .Y(_14617_));
 sky130_fd_sc_hd__a21oi_2 _36665_ (.A1(_14613_),
    .A2(_14616_),
    .B1(_14617_),
    .Y(_14618_));
 sky130_fd_sc_hd__and3_2 _36666_ (.A(_14613_),
    .B(_14617_),
    .C(_14616_),
    .X(_14619_));
 sky130_fd_sc_hd__o22ai_2 _36667_ (.A1(_14586_),
    .A2(_14587_),
    .B1(_14618_),
    .B2(_14619_),
    .Y(_14620_));
 sky130_fd_sc_hd__a21oi_2 _36668_ (.A1(_14598_),
    .A2(_14603_),
    .B1(_14615_),
    .Y(_14621_));
 sky130_fd_sc_hd__nor2_2 _36669_ (.A(_14612_),
    .B(_14604_),
    .Y(_14622_));
 sky130_fd_sc_hd__o21bai_2 _36670_ (.A1(_14621_),
    .A2(_14622_),
    .B1_N(_14617_),
    .Y(_14623_));
 sky130_fd_sc_hd__and2_2 _36671_ (.A(_14581_),
    .B(_14584_),
    .X(_14624_));
 sky130_fd_sc_hd__a21oi_2 _36672_ (.A1(_14624_),
    .A2(_14578_),
    .B1(_14587_),
    .Y(_14625_));
 sky130_fd_sc_hd__nand3_2 _36673_ (.A(_14613_),
    .B(_14616_),
    .C(_14617_),
    .Y(_14626_));
 sky130_fd_sc_hd__nand3_2 _36674_ (.A(_14623_),
    .B(_14625_),
    .C(_14626_),
    .Y(_14627_));
 sky130_fd_sc_hd__a21oi_2 _36675_ (.A1(_14341_),
    .A2(_14342_),
    .B1(_14343_),
    .Y(_14628_));
 sky130_fd_sc_hd__inv_2 _36676_ (.A(_14345_),
    .Y(_14629_));
 sky130_fd_sc_hd__and2_2 _36677_ (.A(_14074_),
    .B(_14071_),
    .X(_14630_));
 sky130_fd_sc_hd__o21ai_2 _36678_ (.A1(_14628_),
    .A2(_14629_),
    .B1(_14630_),
    .Y(_14631_));
 sky130_fd_sc_hd__nor2_2 _36679_ (.A(_14630_),
    .B(_14628_),
    .Y(_14632_));
 sky130_fd_sc_hd__nand2_2 _36680_ (.A(_14632_),
    .B(_14345_),
    .Y(_14633_));
 sky130_fd_sc_hd__nand2_2 _36681_ (.A(_14631_),
    .B(_14633_),
    .Y(_14634_));
 sky130_fd_sc_hd__o21ai_2 _36682_ (.A1(_14634_),
    .A2(_14382_),
    .B1(_14388_),
    .Y(_14635_));
 sky130_fd_sc_hd__nand3_2 _36683_ (.A(_14620_),
    .B(_14627_),
    .C(_14635_),
    .Y(_14636_));
 sky130_fd_sc_hd__o21ai_2 _36684_ (.A1(_14618_),
    .A2(_14619_),
    .B1(_14625_),
    .Y(_14637_));
 sky130_fd_sc_hd__a21oi_2 _36685_ (.A1(_14387_),
    .A2(_14389_),
    .B1(_14384_),
    .Y(_14638_));
 sky130_fd_sc_hd__a21o_2 _36686_ (.A1(_14578_),
    .A2(_14581_),
    .B1(_14584_),
    .X(_14639_));
 sky130_fd_sc_hd__nand2_2 _36687_ (.A(_14639_),
    .B(_14585_),
    .Y(_14640_));
 sky130_fd_sc_hd__nand3_2 _36688_ (.A(_14623_),
    .B(_14626_),
    .C(_14640_),
    .Y(_14641_));
 sky130_fd_sc_hd__nand3_2 _36689_ (.A(_14637_),
    .B(_14638_),
    .C(_14641_),
    .Y(_14642_));
 sky130_fd_sc_hd__a21o_2 _36690_ (.A1(_14306_),
    .A2(_14310_),
    .B1(_14305_),
    .X(_14643_));
 sky130_fd_sc_hd__and4_2 _36691_ (.A(_19338_),
    .B(_10656_),
    .C(_08910_),
    .D(_19579_),
    .X(_14644_));
 sky130_fd_sc_hd__inv_2 _36692_ (.A(_19337_),
    .Y(_14645_));
 sky130_fd_sc_hd__buf_1 _36693_ (.A(_08667_),
    .X(_14646_));
 sky130_fd_sc_hd__o22a_2 _36694_ (.A1(_14645_),
    .A2(_09679_),
    .B1(_14097_),
    .B2(_14646_),
    .X(_14647_));
 sky130_fd_sc_hd__nor2_2 _36695_ (.A(_07718_),
    .B(_12089_),
    .Y(_14648_));
 sky130_fd_sc_hd__o21ai_2 _36696_ (.A1(_14644_),
    .A2(_14647_),
    .B1(_14648_),
    .Y(_14649_));
 sky130_fd_sc_hd__inv_2 _36697_ (.A(_14648_),
    .Y(_14650_));
 sky130_fd_sc_hd__a22o_2 _36698_ (.A1(_19338_),
    .A2(_19579_),
    .B1(_19341_),
    .B2(_19575_),
    .X(_14651_));
 sky130_fd_sc_hd__nand3b_2 _36699_ (.A_N(_14644_),
    .B(_14650_),
    .C(_14651_),
    .Y(_14652_));
 sky130_fd_sc_hd__nand3b_2 _36700_ (.A_N(_14643_),
    .B(_14649_),
    .C(_14652_),
    .Y(_14653_));
 sky130_fd_sc_hd__o21ai_2 _36701_ (.A1(_14644_),
    .A2(_14647_),
    .B1(_14650_),
    .Y(_14654_));
 sky130_fd_sc_hd__nand3b_2 _36702_ (.A_N(_14644_),
    .B(_14651_),
    .C(_14648_),
    .Y(_14655_));
 sky130_fd_sc_hd__nand3_2 _36703_ (.A(_14654_),
    .B(_14655_),
    .C(_14643_),
    .Y(_14656_));
 sky130_fd_sc_hd__nand2_2 _36704_ (.A(_14653_),
    .B(_14656_),
    .Y(_14657_));
 sky130_fd_sc_hd__nor2_2 _36705_ (.A(_07053_),
    .B(_10514_),
    .Y(_14658_));
 sky130_fd_sc_hd__and4_2 _36706_ (.A(_19348_),
    .B(_19351_),
    .C(_09219_),
    .D(_19568_),
    .X(_14659_));
 sky130_fd_sc_hd__a22o_2 _36707_ (.A1(_10210_),
    .A2(_08922_),
    .B1(_08816_),
    .B2(_09219_),
    .X(_14660_));
 sky130_fd_sc_hd__inv_2 _36708_ (.A(_14660_),
    .Y(_14661_));
 sky130_fd_sc_hd__nor3_2 _36709_ (.A(_14658_),
    .B(_14659_),
    .C(_14661_),
    .Y(_14662_));
 sky130_fd_sc_hd__o21ai_2 _36710_ (.A1(_14659_),
    .A2(_14661_),
    .B1(_14658_),
    .Y(_14663_));
 sky130_fd_sc_hd__and2b_2 _36711_ (.A_N(_14662_),
    .B(_14663_),
    .X(_14664_));
 sky130_fd_sc_hd__nand2_2 _36712_ (.A(_14657_),
    .B(_14664_),
    .Y(_14665_));
 sky130_fd_sc_hd__a211o_2 _36713_ (.A1(_19353_),
    .A2(_19563_),
    .B1(_14659_),
    .C1(_14661_),
    .X(_14666_));
 sky130_fd_sc_hd__nand2_2 _36714_ (.A(_14666_),
    .B(_14663_),
    .Y(_14667_));
 sky130_fd_sc_hd__nand3_2 _36715_ (.A(_14667_),
    .B(_14653_),
    .C(_14656_),
    .Y(_14668_));
 sky130_fd_sc_hd__o21ai_2 _36716_ (.A1(_14630_),
    .A2(_14628_),
    .B1(_14345_),
    .Y(_14669_));
 sky130_fd_sc_hd__a21o_2 _36717_ (.A1(_14665_),
    .A2(_14668_),
    .B1(_14669_),
    .X(_14670_));
 sky130_fd_sc_hd__nand3_2 _36718_ (.A(_14665_),
    .B(_14669_),
    .C(_14668_),
    .Y(_14671_));
 sky130_fd_sc_hd__nand2_2 _36719_ (.A(_14315_),
    .B(_14323_),
    .Y(_14672_));
 sky130_fd_sc_hd__nand2_2 _36720_ (.A(_14672_),
    .B(_14312_),
    .Y(_14673_));
 sky130_fd_sc_hd__a21oi_2 _36721_ (.A1(_14670_),
    .A2(_14671_),
    .B1(_14673_),
    .Y(_14674_));
 sky130_fd_sc_hd__nand3_2 _36722_ (.A(_14670_),
    .B(_14671_),
    .C(_14673_),
    .Y(_14675_));
 sky130_fd_sc_hd__inv_2 _36723_ (.A(_14675_),
    .Y(_14676_));
 sky130_fd_sc_hd__o2bb2ai_2 _36724_ (.A1_N(_14636_),
    .A2_N(_14642_),
    .B1(_14674_),
    .B2(_14676_),
    .Y(_14677_));
 sky130_fd_sc_hd__inv_2 _36725_ (.A(_14673_),
    .Y(_14678_));
 sky130_fd_sc_hd__a21oi_2 _36726_ (.A1(_14665_),
    .A2(_14668_),
    .B1(_14669_),
    .Y(_14679_));
 sky130_fd_sc_hd__nor2_2 _36727_ (.A(_14678_),
    .B(_14679_),
    .Y(_14680_));
 sky130_fd_sc_hd__a21oi_2 _36728_ (.A1(_14680_),
    .A2(_14671_),
    .B1(_14674_),
    .Y(_14681_));
 sky130_fd_sc_hd__nand3_2 _36729_ (.A(_14681_),
    .B(_14642_),
    .C(_14636_),
    .Y(_14682_));
 sky130_fd_sc_hd__o21ai_2 _36730_ (.A1(_14410_),
    .A2(_14394_),
    .B1(_14401_),
    .Y(_14683_));
 sky130_fd_sc_hd__a21oi_2 _36731_ (.A1(_14677_),
    .A2(_14682_),
    .B1(_14683_),
    .Y(_14684_));
 sky130_fd_sc_hd__and3_2 _36732_ (.A(_14620_),
    .B(_14627_),
    .C(_14635_),
    .X(_14685_));
 sky130_fd_sc_hd__nand2_2 _36733_ (.A(_14681_),
    .B(_14642_),
    .Y(_14686_));
 sky130_fd_sc_hd__o211a_2 _36734_ (.A1(_14685_),
    .A2(_14686_),
    .B1(_14677_),
    .C1(_14683_),
    .X(_14687_));
 sky130_fd_sc_hd__nand2_2 _36735_ (.A(_14453_),
    .B(_14448_),
    .Y(_14688_));
 sky130_fd_sc_hd__nand2_2 _36736_ (.A(_07886_),
    .B(_09203_),
    .Y(_14689_));
 sky130_fd_sc_hd__nand2_2 _36737_ (.A(_08345_),
    .B(_11410_),
    .Y(_14690_));
 sky130_fd_sc_hd__and2_2 _36738_ (.A(_14689_),
    .B(_14690_),
    .X(_14691_));
 sky130_fd_sc_hd__nor2_2 _36739_ (.A(_08352_),
    .B(_10533_),
    .Y(_14692_));
 sky130_fd_sc_hd__or2_2 _36740_ (.A(_14689_),
    .B(_14690_),
    .X(_14693_));
 sky130_fd_sc_hd__nand3b_2 _36741_ (.A_N(_14691_),
    .B(_14692_),
    .C(_14693_),
    .Y(_14694_));
 sky130_fd_sc_hd__nor2_2 _36742_ (.A(_14689_),
    .B(_14690_),
    .Y(_14695_));
 sky130_fd_sc_hd__o21bai_2 _36743_ (.A1(_14695_),
    .A2(_14691_),
    .B1_N(_14692_),
    .Y(_14696_));
 sky130_fd_sc_hd__a21o_2 _36744_ (.A1(_14318_),
    .A2(_14321_),
    .B1(_14316_),
    .X(_14697_));
 sky130_fd_sc_hd__a21oi_2 _36745_ (.A1(_14694_),
    .A2(_14696_),
    .B1(_14697_),
    .Y(_14698_));
 sky130_fd_sc_hd__and3_2 _36746_ (.A(_14694_),
    .B(_14697_),
    .C(_14696_),
    .X(_14699_));
 sky130_fd_sc_hd__and2_2 _36747_ (.A(_14441_),
    .B(_14439_),
    .X(_14700_));
 sky130_fd_sc_hd__o21ai_2 _36748_ (.A1(_14698_),
    .A2(_14699_),
    .B1(_14700_),
    .Y(_14701_));
 sky130_fd_sc_hd__nand3_2 _36749_ (.A(_14694_),
    .B(_14697_),
    .C(_14696_),
    .Y(_14702_));
 sky130_fd_sc_hd__nand2_2 _36750_ (.A(_14441_),
    .B(_14439_),
    .Y(_14703_));
 sky130_fd_sc_hd__nand3b_2 _36751_ (.A_N(_14698_),
    .B(_14702_),
    .C(_14703_),
    .Y(_14704_));
 sky130_fd_sc_hd__and3_2 _36752_ (.A(_14688_),
    .B(_14701_),
    .C(_14704_),
    .X(_14705_));
 sky130_fd_sc_hd__a21o_2 _36753_ (.A1(_14701_),
    .A2(_14704_),
    .B1(_14688_),
    .X(_14706_));
 sky130_fd_sc_hd__nand2_2 _36754_ (.A(_06278_),
    .B(_19544_),
    .Y(_14707_));
 sky130_fd_sc_hd__nand2_2 _36755_ (.A(_07450_),
    .B(_19540_),
    .Y(_14708_));
 sky130_fd_sc_hd__nor2_2 _36756_ (.A(_14707_),
    .B(_14708_),
    .Y(_14709_));
 sky130_fd_sc_hd__nand2_2 _36757_ (.A(_14707_),
    .B(_14708_),
    .Y(_14710_));
 sky130_fd_sc_hd__inv_2 _36758_ (.A(_14710_),
    .Y(_14711_));
 sky130_fd_sc_hd__nand2_2 _36759_ (.A(_14153_),
    .B(_19368_),
    .Y(_14712_));
 sky130_fd_sc_hd__o21ai_2 _36760_ (.A1(_14709_),
    .A2(_14711_),
    .B1(_14712_),
    .Y(_14713_));
 sky130_fd_sc_hd__inv_2 _36761_ (.A(_14709_),
    .Y(_14714_));
 sky130_fd_sc_hd__inv_2 _36762_ (.A(_14712_),
    .Y(_14715_));
 sky130_fd_sc_hd__nand3_2 _36763_ (.A(_14714_),
    .B(_14715_),
    .C(_14710_),
    .Y(_14716_));
 sky130_fd_sc_hd__a31o_2 _36764_ (.A1(_14420_),
    .A2(_19369_),
    .A3(_19542_),
    .B1(_14419_),
    .X(_14717_));
 sky130_fd_sc_hd__a21o_2 _36765_ (.A1(_14713_),
    .A2(_14716_),
    .B1(_14717_),
    .X(_14718_));
 sky130_fd_sc_hd__nand3_2 _36766_ (.A(_14713_),
    .B(_14716_),
    .C(_14717_),
    .Y(_14719_));
 sky130_fd_sc_hd__a21oi_2 _36767_ (.A1(_14718_),
    .A2(_14719_),
    .B1(_14430_),
    .Y(_14720_));
 sky130_fd_sc_hd__and3_2 _36768_ (.A(_14718_),
    .B(_14429_),
    .C(_14719_),
    .X(_14721_));
 sky130_fd_sc_hd__nor2_2 _36769_ (.A(_14720_),
    .B(_14721_),
    .Y(_14722_));
 sky130_fd_sc_hd__nand2_2 _36770_ (.A(_14706_),
    .B(_14722_),
    .Y(_14723_));
 sky130_fd_sc_hd__a21oi_2 _36771_ (.A1(_14324_),
    .A2(_14325_),
    .B1(_14326_),
    .Y(_14724_));
 sky130_fd_sc_hd__o21ai_2 _36772_ (.A1(_14407_),
    .A2(_14724_),
    .B1(_14328_),
    .Y(_14725_));
 sky130_fd_sc_hd__a21oi_2 _36773_ (.A1(_14701_),
    .A2(_14704_),
    .B1(_14688_),
    .Y(_14726_));
 sky130_fd_sc_hd__or2_2 _36774_ (.A(_14720_),
    .B(_14721_),
    .X(_14727_));
 sky130_fd_sc_hd__o21ai_2 _36775_ (.A1(_14726_),
    .A2(_14705_),
    .B1(_14727_),
    .Y(_14728_));
 sky130_fd_sc_hd__o211a_2 _36776_ (.A1(_14705_),
    .A2(_14723_),
    .B1(_14725_),
    .C1(_14728_),
    .X(_14729_));
 sky130_fd_sc_hd__nand3_2 _36777_ (.A(_14688_),
    .B(_14701_),
    .C(_14704_),
    .Y(_14730_));
 sky130_fd_sc_hd__nand3_2 _36778_ (.A(_14706_),
    .B(_14730_),
    .C(_14722_),
    .Y(_14731_));
 sky130_fd_sc_hd__a21o_2 _36779_ (.A1(_14728_),
    .A2(_14731_),
    .B1(_14725_),
    .X(_14732_));
 sky130_fd_sc_hd__nand2_2 _36780_ (.A(_14456_),
    .B(_14457_),
    .Y(_14733_));
 sky130_fd_sc_hd__nand2_2 _36781_ (.A(_14733_),
    .B(_14458_),
    .Y(_14734_));
 sky130_fd_sc_hd__nand2_2 _36782_ (.A(_14732_),
    .B(_14734_),
    .Y(_14735_));
 sky130_fd_sc_hd__nor2_2 _36783_ (.A(_14457_),
    .B(_14454_),
    .Y(_14736_));
 sky130_fd_sc_hd__a21oi_2 _36784_ (.A1(_14728_),
    .A2(_14731_),
    .B1(_14725_),
    .Y(_14737_));
 sky130_fd_sc_hd__o22ai_2 _36785_ (.A1(_14452_),
    .A2(_14736_),
    .B1(_14737_),
    .B2(_14729_),
    .Y(_14738_));
 sky130_fd_sc_hd__o21a_2 _36786_ (.A1(_14729_),
    .A2(_14735_),
    .B1(_14738_),
    .X(_14739_));
 sky130_fd_sc_hd__o21ai_2 _36787_ (.A1(_14684_),
    .A2(_14687_),
    .B1(_14739_),
    .Y(_14740_));
 sky130_fd_sc_hd__a21oi_2 _36788_ (.A1(_14404_),
    .A2(_14411_),
    .B1(_14405_),
    .Y(_14741_));
 sky130_fd_sc_hd__a21oi_2 _36789_ (.A1(_14472_),
    .A2(_14412_),
    .B1(_14741_),
    .Y(_14742_));
 sky130_fd_sc_hd__a21o_2 _36790_ (.A1(_14677_),
    .A2(_14682_),
    .B1(_14683_),
    .X(_14743_));
 sky130_fd_sc_hd__nand3_2 _36791_ (.A(_14683_),
    .B(_14677_),
    .C(_14682_),
    .Y(_14744_));
 sky130_fd_sc_hd__nand3_2 _36792_ (.A(_14728_),
    .B(_14725_),
    .C(_14731_),
    .Y(_14745_));
 sky130_fd_sc_hd__nand3_2 _36793_ (.A(_14732_),
    .B(_14745_),
    .C(_14734_),
    .Y(_14746_));
 sky130_fd_sc_hd__nand2_2 _36794_ (.A(_14738_),
    .B(_14746_),
    .Y(_14747_));
 sky130_fd_sc_hd__nand3_2 _36795_ (.A(_14743_),
    .B(_14744_),
    .C(_14747_),
    .Y(_14748_));
 sky130_fd_sc_hd__nand3_2 _36796_ (.A(_14740_),
    .B(_14742_),
    .C(_14748_),
    .Y(_14749_));
 sky130_fd_sc_hd__a31oi_2 _36797_ (.A1(_14405_),
    .A2(_14404_),
    .A3(_14411_),
    .B1(_14477_),
    .Y(_14750_));
 sky130_fd_sc_hd__nand3_2 _36798_ (.A(_14739_),
    .B(_14743_),
    .C(_14744_),
    .Y(_14751_));
 sky130_fd_sc_hd__o21ai_2 _36799_ (.A1(_14684_),
    .A2(_14687_),
    .B1(_14747_),
    .Y(_14752_));
 sky130_fd_sc_hd__o211ai_2 _36800_ (.A1(_14741_),
    .A2(_14750_),
    .B1(_14751_),
    .C1(_14752_),
    .Y(_14753_));
 sky130_fd_sc_hd__a21boi_2 _36801_ (.A1(_14425_),
    .A2(_06020_),
    .B1_N(_14426_),
    .Y(_14754_));
 sky130_fd_sc_hd__nand2_2 _36802_ (.A(_14212_),
    .B(_14754_),
    .Y(_14755_));
 sky130_fd_sc_hd__nand3b_2 _36803_ (.A_N(_14754_),
    .B(_13667_),
    .C(_13669_),
    .Y(_14756_));
 sky130_fd_sc_hd__a21oi_2 _36804_ (.A1(_14755_),
    .A2(_14756_),
    .B1(_14217_),
    .Y(_14757_));
 sky130_fd_sc_hd__and3_2 _36805_ (.A(_14755_),
    .B(_13965_),
    .C(_14756_),
    .X(_14758_));
 sky130_fd_sc_hd__o21ai_2 _36806_ (.A1(_05498_),
    .A2(_14427_),
    .B1(_14428_),
    .Y(_14759_));
 sky130_fd_sc_hd__a21oi_2 _36807_ (.A1(_14418_),
    .A2(_14421_),
    .B1(_14422_),
    .Y(_14760_));
 sky130_fd_sc_hd__o21a_2 _36808_ (.A1(_14759_),
    .A2(_14760_),
    .B1(_14424_),
    .X(_14761_));
 sky130_fd_sc_hd__o21ai_2 _36809_ (.A1(_14757_),
    .A2(_14758_),
    .B1(_14761_),
    .Y(_14762_));
 sky130_fd_sc_hd__and3_2 _36810_ (.A(_13663_),
    .B(_14754_),
    .C(_13664_),
    .X(_14763_));
 sky130_fd_sc_hd__nor2_2 _36811_ (.A(_14754_),
    .B(_14212_),
    .Y(_14764_));
 sky130_fd_sc_hd__inv_2 _36812_ (.A(_13963_),
    .Y(_14765_));
 sky130_fd_sc_hd__o21ai_2 _36813_ (.A1(_14763_),
    .A2(_14764_),
    .B1(_14765_),
    .Y(_14766_));
 sky130_fd_sc_hd__o21ai_2 _36814_ (.A1(_14759_),
    .A2(_14760_),
    .B1(_14424_),
    .Y(_14767_));
 sky130_fd_sc_hd__nand3_2 _36815_ (.A(_14755_),
    .B(_13965_),
    .C(_14756_),
    .Y(_14768_));
 sky130_fd_sc_hd__nand3_2 _36816_ (.A(_14766_),
    .B(_14767_),
    .C(_14768_),
    .Y(_14769_));
 sky130_fd_sc_hd__inv_2 _36817_ (.A(_14487_),
    .Y(_14770_));
 sky130_fd_sc_hd__a21o_2 _36818_ (.A1(_14486_),
    .A2(_14217_),
    .B1(_14770_),
    .X(_14771_));
 sky130_fd_sc_hd__a21oi_2 _36819_ (.A1(_14762_),
    .A2(_14769_),
    .B1(_14771_),
    .Y(_14772_));
 sky130_fd_sc_hd__nand2_2 _36820_ (.A(_14766_),
    .B(_14767_),
    .Y(_14773_));
 sky130_fd_sc_hd__o211a_2 _36821_ (.A1(_14758_),
    .A2(_14773_),
    .B1(_14771_),
    .C1(_14762_),
    .X(_14774_));
 sky130_fd_sc_hd__nor2_2 _36822_ (.A(_14499_),
    .B(_14500_),
    .Y(_14775_));
 sky130_fd_sc_hd__a21oi_2 _36823_ (.A1(_14497_),
    .A2(_14496_),
    .B1(_14495_),
    .Y(_14776_));
 sky130_fd_sc_hd__o21a_2 _36824_ (.A1(_14775_),
    .A2(_14776_),
    .B1(_14498_),
    .X(_14777_));
 sky130_fd_sc_hd__o21ai_2 _36825_ (.A1(_14772_),
    .A2(_14774_),
    .B1(_14777_),
    .Y(_14778_));
 sky130_fd_sc_hd__nand2_2 _36826_ (.A(_14762_),
    .B(_14769_),
    .Y(_14779_));
 sky130_fd_sc_hd__inv_2 _36827_ (.A(_14771_),
    .Y(_14780_));
 sky130_fd_sc_hd__nand2_2 _36828_ (.A(_14779_),
    .B(_14780_),
    .Y(_14781_));
 sky130_fd_sc_hd__o21ai_2 _36829_ (.A1(_14775_),
    .A2(_14776_),
    .B1(_14498_),
    .Y(_14782_));
 sky130_fd_sc_hd__nand3_2 _36830_ (.A(_14762_),
    .B(_14769_),
    .C(_14771_),
    .Y(_14783_));
 sky130_fd_sc_hd__nand3_2 _36831_ (.A(_14781_),
    .B(_14782_),
    .C(_14783_),
    .Y(_14784_));
 sky130_fd_sc_hd__a21oi_2 _36832_ (.A1(_14778_),
    .A2(_14784_),
    .B1(_14248_),
    .Y(_14785_));
 sky130_fd_sc_hd__nand2_2 _36833_ (.A(_14781_),
    .B(_14782_),
    .Y(_14786_));
 sky130_fd_sc_hd__o211a_2 _36834_ (.A1(_14774_),
    .A2(_14786_),
    .B1(_13402_),
    .C1(_14778_),
    .X(_14787_));
 sky130_fd_sc_hd__o21a_2 _36835_ (.A1(_14463_),
    .A2(_14470_),
    .B1(_14462_),
    .X(_14788_));
 sky130_fd_sc_hd__o21ai_2 _36836_ (.A1(_14785_),
    .A2(_14787_),
    .B1(_14788_),
    .Y(_14789_));
 sky130_fd_sc_hd__a21o_2 _36837_ (.A1(_14778_),
    .A2(_14784_),
    .B1(_13402_),
    .X(_14790_));
 sky130_fd_sc_hd__o21ai_2 _36838_ (.A1(_14463_),
    .A2(_14470_),
    .B1(_14462_),
    .Y(_14791_));
 sky130_fd_sc_hd__nand3_2 _36839_ (.A(_14778_),
    .B(_14248_),
    .C(_14784_),
    .Y(_14792_));
 sky130_fd_sc_hd__nand3_2 _36840_ (.A(_14790_),
    .B(_14791_),
    .C(_14792_),
    .Y(_14793_));
 sky130_fd_sc_hd__buf_1 _36841_ (.A(_13398_),
    .X(_14794_));
 sky130_fd_sc_hd__inv_2 _36842_ (.A(_14509_),
    .Y(_14795_));
 sky130_fd_sc_hd__a21o_2 _36843_ (.A1(_14794_),
    .A2(_14505_),
    .B1(_14795_),
    .X(_14796_));
 sky130_fd_sc_hd__a21oi_2 _36844_ (.A1(_14789_),
    .A2(_14793_),
    .B1(_14796_),
    .Y(_14797_));
 sky130_fd_sc_hd__and2_2 _36845_ (.A(_14505_),
    .B(_14248_),
    .X(_14798_));
 sky130_fd_sc_hd__o211a_2 _36846_ (.A1(_14795_),
    .A2(_14798_),
    .B1(_14793_),
    .C1(_14789_),
    .X(_14799_));
 sky130_fd_sc_hd__o2bb2ai_2 _36847_ (.A1_N(_14749_),
    .A2_N(_14753_),
    .B1(_14797_),
    .B2(_14799_),
    .Y(_14800_));
 sky130_fd_sc_hd__nor2_2 _36848_ (.A(_14797_),
    .B(_14799_),
    .Y(_14801_));
 sky130_fd_sc_hd__nand3_2 _36849_ (.A(_14753_),
    .B(_14749_),
    .C(_14801_),
    .Y(_14802_));
 sky130_fd_sc_hd__nand2_2 _36850_ (.A(_14534_),
    .B(_14474_),
    .Y(_14803_));
 sky130_fd_sc_hd__a21oi_2 _36851_ (.A1(_14800_),
    .A2(_14802_),
    .B1(_14803_),
    .Y(_14804_));
 sky130_fd_sc_hd__inv_2 _36852_ (.A(_14243_),
    .Y(_14805_));
 sky130_fd_sc_hd__inv_2 _36853_ (.A(_14483_),
    .Y(_14806_));
 sky130_fd_sc_hd__a21oi_2 _36854_ (.A1(_14520_),
    .A2(_14519_),
    .B1(_14518_),
    .Y(_14807_));
 sky130_fd_sc_hd__o211a_2 _36855_ (.A1(_14513_),
    .A2(_14193_),
    .B1(_14519_),
    .C1(_14520_),
    .X(_14808_));
 sky130_fd_sc_hd__o22ai_2 _36856_ (.A1(_14805_),
    .A2(_14806_),
    .B1(_14807_),
    .B2(_14808_),
    .Y(_14809_));
 sky130_fd_sc_hd__o211ai_2 _36857_ (.A1(_14239_),
    .A2(_14523_),
    .B1(_14521_),
    .C1(_14515_),
    .Y(_14810_));
 sky130_fd_sc_hd__nand2_2 _36858_ (.A(_14809_),
    .B(_14810_),
    .Y(_14811_));
 sky130_fd_sc_hd__a31oi_2 _36859_ (.A1(_14479_),
    .A2(_14480_),
    .A3(_14478_),
    .B1(_14811_),
    .Y(_14812_));
 sky130_fd_sc_hd__o211a_2 _36860_ (.A1(_14533_),
    .A2(_14812_),
    .B1(_14802_),
    .C1(_14800_),
    .X(_14813_));
 sky130_fd_sc_hd__nand2_2 _36861_ (.A(_14810_),
    .B(_14521_),
    .Y(_14814_));
 sky130_fd_sc_hd__xor2_2 _36862_ (.A(_14017_),
    .B(_14814_),
    .X(_14815_));
 sky130_fd_sc_hd__inv_2 _36863_ (.A(_14815_),
    .Y(_14816_));
 sky130_fd_sc_hd__o21ai_2 _36864_ (.A1(_14804_),
    .A2(_14813_),
    .B1(_14816_),
    .Y(_14817_));
 sky130_fd_sc_hd__a21oi_2 _36865_ (.A1(_14544_),
    .A2(_14541_),
    .B1(_14535_),
    .Y(_14818_));
 sky130_fd_sc_hd__a21o_2 _36866_ (.A1(_14800_),
    .A2(_14802_),
    .B1(_14803_),
    .X(_14819_));
 sky130_fd_sc_hd__nand3_2 _36867_ (.A(_14803_),
    .B(_14800_),
    .C(_14802_),
    .Y(_14820_));
 sky130_fd_sc_hd__nand3_2 _36868_ (.A(_14819_),
    .B(_14820_),
    .C(_14815_),
    .Y(_14821_));
 sky130_fd_sc_hd__nand3_2 _36869_ (.A(_14817_),
    .B(_14818_),
    .C(_14821_),
    .Y(_14822_));
 sky130_fd_sc_hd__buf_1 _36870_ (.A(_13725_),
    .X(_14823_));
 sky130_fd_sc_hd__inv_2 _36871_ (.A(_14814_),
    .Y(_14824_));
 sky130_fd_sc_hd__nor2_2 _36872_ (.A(_14823_),
    .B(_14824_),
    .Y(_14825_));
 sky130_fd_sc_hd__nor2_2 _36873_ (.A(_13737_),
    .B(_14814_),
    .Y(_14826_));
 sky130_fd_sc_hd__o22ai_2 _36874_ (.A1(_14825_),
    .A2(_14826_),
    .B1(_14804_),
    .B2(_14813_),
    .Y(_14827_));
 sky130_fd_sc_hd__nand3_2 _36875_ (.A(_14819_),
    .B(_14820_),
    .C(_14816_),
    .Y(_14828_));
 sky130_fd_sc_hd__o21ai_2 _36876_ (.A1(_14546_),
    .A2(_14532_),
    .B1(_14545_),
    .Y(_14829_));
 sky130_fd_sc_hd__nand3_2 _36877_ (.A(_14827_),
    .B(_14828_),
    .C(_14829_),
    .Y(_14830_));
 sky130_fd_sc_hd__a21o_2 _36878_ (.A1(_14822_),
    .A2(_14830_),
    .B1(_14549_),
    .X(_14831_));
 sky130_fd_sc_hd__nand2_2 _36879_ (.A(_14548_),
    .B(_14273_),
    .Y(_14832_));
 sky130_fd_sc_hd__nand2_2 _36880_ (.A(_14832_),
    .B(_14554_),
    .Y(_14833_));
 sky130_fd_sc_hd__nand3_2 _36881_ (.A(_14822_),
    .B(_14830_),
    .C(_14549_),
    .Y(_14834_));
 sky130_fd_sc_hd__nand3_2 _36882_ (.A(_14831_),
    .B(_14833_),
    .C(_14834_),
    .Y(_14835_));
 sky130_fd_sc_hd__inv_2 _36883_ (.A(_14835_),
    .Y(_14836_));
 sky130_fd_sc_hd__a21oi_2 _36884_ (.A1(_14822_),
    .A2(_14830_),
    .B1(_14549_),
    .Y(_14837_));
 sky130_fd_sc_hd__and3_2 _36885_ (.A(_14822_),
    .B(_14830_),
    .C(_14549_),
    .X(_14838_));
 sky130_fd_sc_hd__o21bai_2 _36886_ (.A1(_14837_),
    .A2(_14838_),
    .B1_N(_14833_),
    .Y(_14839_));
 sky130_fd_sc_hd__inv_2 _36887_ (.A(_14839_),
    .Y(_14840_));
 sky130_fd_sc_hd__nor2_2 _36888_ (.A(_14836_),
    .B(_14840_),
    .Y(_14841_));
 sky130_fd_sc_hd__nand3_2 _36889_ (.A(_14295_),
    .B(_14563_),
    .C(_14294_),
    .Y(_14842_));
 sky130_fd_sc_hd__inv_2 _36890_ (.A(_14555_),
    .Y(_14843_));
 sky130_fd_sc_hd__nand2_2 _36891_ (.A(_14561_),
    .B(_14560_),
    .Y(_14844_));
 sky130_fd_sc_hd__a21o_2 _36892_ (.A1(_14560_),
    .A2(_14555_),
    .B1(_14561_),
    .X(_14845_));
 sky130_fd_sc_hd__o2111ai_2 _36893_ (.A1(_14843_),
    .A2(_14844_),
    .B1(_14293_),
    .C1(_14303_),
    .D1(_14845_),
    .Y(_14846_));
 sky130_fd_sc_hd__nand2_2 _36894_ (.A(_14559_),
    .B(_14555_),
    .Y(_14847_));
 sky130_fd_sc_hd__o21a_2 _36895_ (.A1(_14562_),
    .A2(_14303_),
    .B1(_14847_),
    .X(_14848_));
 sky130_fd_sc_hd__o21ai_2 _36896_ (.A1(_14298_),
    .A2(_14846_),
    .B1(_14848_),
    .Y(_14849_));
 sky130_fd_sc_hd__o21bai_2 _36897_ (.A1(_14842_),
    .A2(_13766_),
    .B1_N(_14849_),
    .Y(_14850_));
 sky130_fd_sc_hd__xor2_2 _36898_ (.A(_14841_),
    .B(_14850_),
    .X(_02663_));
 sky130_fd_sc_hd__nand2_2 _36899_ (.A(_14749_),
    .B(_14801_),
    .Y(_14851_));
 sky130_fd_sc_hd__nand2_2 _36900_ (.A(_14851_),
    .B(_14753_),
    .Y(_14852_));
 sky130_fd_sc_hd__o21ai_2 _36901_ (.A1(_14640_),
    .A2(_14618_),
    .B1(_14626_),
    .Y(_14853_));
 sky130_fd_sc_hd__and4_2 _36902_ (.A(_14349_),
    .B(_11122_),
    .C(_14351_),
    .D(_19598_),
    .X(_14854_));
 sky130_fd_sc_hd__buf_1 _36903_ (.A(_11164_),
    .X(_14855_));
 sky130_fd_sc_hd__o22a_2 _36904_ (.A1(_06222_),
    .A2(_18182_),
    .B1(_14855_),
    .B2(_06401_),
    .X(_14856_));
 sky130_fd_sc_hd__nand2_2 _36905_ (.A(_19312_),
    .B(_06954_),
    .Y(_14857_));
 sky130_fd_sc_hd__o21ai_2 _36906_ (.A1(_14854_),
    .A2(_14856_),
    .B1(_14857_),
    .Y(_14858_));
 sky130_fd_sc_hd__a22o_2 _36907_ (.A1(_14351_),
    .A2(_19598_),
    .B1(_14349_),
    .B2(_14350_),
    .X(_14859_));
 sky130_fd_sc_hd__and3_2 _36908_ (.A(_11169_),
    .B(_13146_),
    .C(_19597_),
    .X(_14860_));
 sky130_fd_sc_hd__nand2_2 _36909_ (.A(_14860_),
    .B(_14349_),
    .Y(_14861_));
 sky130_fd_sc_hd__inv_2 _36910_ (.A(_14857_),
    .Y(_14862_));
 sky130_fd_sc_hd__nand3_2 _36911_ (.A(_14859_),
    .B(_14861_),
    .C(_14862_),
    .Y(_14863_));
 sky130_fd_sc_hd__o21ai_2 _36912_ (.A1(_14589_),
    .A2(_14588_),
    .B1(_14594_),
    .Y(_14864_));
 sky130_fd_sc_hd__a21oi_2 _36913_ (.A1(_14858_),
    .A2(_14863_),
    .B1(_14864_),
    .Y(_14865_));
 sky130_fd_sc_hd__and3_2 _36914_ (.A(_14858_),
    .B(_14864_),
    .C(_14863_),
    .X(_14866_));
 sky130_fd_sc_hd__and4_2 _36915_ (.A(_10139_),
    .B(_14042_),
    .C(_19589_),
    .D(_19591_),
    .X(_14867_));
 sky130_fd_sc_hd__inv_2 _36916_ (.A(_19319_),
    .Y(_14868_));
 sky130_fd_sc_hd__buf_1 _36917_ (.A(_14868_),
    .X(_14869_));
 sky130_fd_sc_hd__o22a_2 _36918_ (.A1(_14371_),
    .A2(_10279_),
    .B1(_14869_),
    .B2(_07833_),
    .X(_14870_));
 sky130_fd_sc_hd__nor2_2 _36919_ (.A(_14867_),
    .B(_14870_),
    .Y(_14871_));
 sky130_fd_sc_hd__nor2_2 _36920_ (.A(_09358_),
    .B(_08611_),
    .Y(_14872_));
 sky130_fd_sc_hd__nand2_2 _36921_ (.A(_14871_),
    .B(_14872_),
    .Y(_14873_));
 sky130_fd_sc_hd__inv_2 _36922_ (.A(_14872_),
    .Y(_14874_));
 sky130_fd_sc_hd__o21ai_2 _36923_ (.A1(_14867_),
    .A2(_14870_),
    .B1(_14874_),
    .Y(_14875_));
 sky130_fd_sc_hd__nand2_2 _36924_ (.A(_14873_),
    .B(_14875_),
    .Y(_14876_));
 sky130_fd_sc_hd__o21ai_2 _36925_ (.A1(_14865_),
    .A2(_14866_),
    .B1(_14876_),
    .Y(_14877_));
 sky130_fd_sc_hd__a21oi_2 _36926_ (.A1(_14601_),
    .A2(_14602_),
    .B1(_14599_),
    .Y(_14878_));
 sky130_fd_sc_hd__o21ai_2 _36927_ (.A1(_14612_),
    .A2(_14878_),
    .B1(_14603_),
    .Y(_14879_));
 sky130_fd_sc_hd__a21o_2 _36928_ (.A1(_14858_),
    .A2(_14863_),
    .B1(_14864_),
    .X(_14880_));
 sky130_fd_sc_hd__nand3_2 _36929_ (.A(_14858_),
    .B(_14864_),
    .C(_14863_),
    .Y(_14881_));
 sky130_fd_sc_hd__nand2_2 _36930_ (.A(_14871_),
    .B(_14874_),
    .Y(_14882_));
 sky130_fd_sc_hd__o21ai_2 _36931_ (.A1(_14867_),
    .A2(_14870_),
    .B1(_14872_),
    .Y(_14883_));
 sky130_fd_sc_hd__nand2_2 _36932_ (.A(_14882_),
    .B(_14883_),
    .Y(_14884_));
 sky130_fd_sc_hd__nand3_2 _36933_ (.A(_14880_),
    .B(_14881_),
    .C(_14884_),
    .Y(_14885_));
 sky130_fd_sc_hd__nand3_2 _36934_ (.A(_14877_),
    .B(_14879_),
    .C(_14885_),
    .Y(_14886_));
 sky130_fd_sc_hd__o21a_2 _36935_ (.A1(_14612_),
    .A2(_14878_),
    .B1(_14603_),
    .X(_14887_));
 sky130_fd_sc_hd__o21bai_2 _36936_ (.A1(_14865_),
    .A2(_14866_),
    .B1_N(_14876_),
    .Y(_14888_));
 sky130_fd_sc_hd__nand3_2 _36937_ (.A(_14880_),
    .B(_14881_),
    .C(_14876_),
    .Y(_14889_));
 sky130_fd_sc_hd__nand3_2 _36938_ (.A(_14887_),
    .B(_14888_),
    .C(_14889_),
    .Y(_14890_));
 sky130_fd_sc_hd__nand2_2 _36939_ (.A(_11205_),
    .B(_09933_),
    .Y(_14891_));
 sky130_fd_sc_hd__nand2_2 _36940_ (.A(_10867_),
    .B(_08108_),
    .Y(_14892_));
 sky130_fd_sc_hd__nand2_2 _36941_ (.A(_14891_),
    .B(_14892_),
    .Y(_14893_));
 sky130_fd_sc_hd__or2_2 _36942_ (.A(_14891_),
    .B(_14892_),
    .X(_14894_));
 sky130_fd_sc_hd__o2bb2ai_2 _36943_ (.A1_N(_14893_),
    .A2_N(_14894_),
    .B1(_08424_),
    .B2(_09679_),
    .Y(_14895_));
 sky130_fd_sc_hd__nor2_2 _36944_ (.A(_14339_),
    .B(_09679_),
    .Y(_14896_));
 sky130_fd_sc_hd__nand3_2 _36945_ (.A(_14894_),
    .B(_14896_),
    .C(_14893_),
    .Y(_14897_));
 sky130_fd_sc_hd__nor2_2 _36946_ (.A(_14607_),
    .B(_14608_),
    .Y(_14898_));
 sky130_fd_sc_hd__nor2_2 _36947_ (.A(_14605_),
    .B(_14898_),
    .Y(_14899_));
 sky130_fd_sc_hd__a21o_2 _36948_ (.A1(_14895_),
    .A2(_14897_),
    .B1(_14899_),
    .X(_14900_));
 sky130_fd_sc_hd__nand3_2 _36949_ (.A(_14895_),
    .B(_14899_),
    .C(_14897_),
    .Y(_14901_));
 sky130_fd_sc_hd__nor2_2 _36950_ (.A(_14574_),
    .B(_14570_),
    .Y(_14902_));
 sky130_fd_sc_hd__nor2_2 _36951_ (.A(_14572_),
    .B(_14902_),
    .Y(_14903_));
 sky130_fd_sc_hd__a21oi_2 _36952_ (.A1(_14900_),
    .A2(_14901_),
    .B1(_14903_),
    .Y(_14904_));
 sky130_fd_sc_hd__nand3_2 _36953_ (.A(_14900_),
    .B(_14901_),
    .C(_14903_),
    .Y(_14905_));
 sky130_fd_sc_hd__inv_2 _36954_ (.A(_14905_),
    .Y(_14906_));
 sky130_fd_sc_hd__o2bb2ai_2 _36955_ (.A1_N(_14886_),
    .A2_N(_14890_),
    .B1(_14904_),
    .B2(_14906_),
    .Y(_14907_));
 sky130_fd_sc_hd__inv_2 _36956_ (.A(_14903_),
    .Y(_14908_));
 sky130_fd_sc_hd__a21oi_2 _36957_ (.A1(_14895_),
    .A2(_14897_),
    .B1(_14899_),
    .Y(_14909_));
 sky130_fd_sc_hd__nor2_2 _36958_ (.A(_14908_),
    .B(_14909_),
    .Y(_14910_));
 sky130_fd_sc_hd__a21oi_2 _36959_ (.A1(_14901_),
    .A2(_14910_),
    .B1(_14904_),
    .Y(_14911_));
 sky130_fd_sc_hd__nand3_2 _36960_ (.A(_14911_),
    .B(_14890_),
    .C(_14886_),
    .Y(_14912_));
 sky130_fd_sc_hd__nand3_2 _36961_ (.A(_14853_),
    .B(_14907_),
    .C(_14912_),
    .Y(_14913_));
 sky130_fd_sc_hd__a21oi_2 _36962_ (.A1(_14623_),
    .A2(_14625_),
    .B1(_14619_),
    .Y(_14914_));
 sky130_fd_sc_hd__nand2_2 _36963_ (.A(_14890_),
    .B(_14886_),
    .Y(_14915_));
 sky130_fd_sc_hd__nand2_2 _36964_ (.A(_14915_),
    .B(_14911_),
    .Y(_14916_));
 sky130_fd_sc_hd__and3_2 _36965_ (.A(_14895_),
    .B(_14899_),
    .C(_14897_),
    .X(_14917_));
 sky130_fd_sc_hd__o21ai_2 _36966_ (.A1(_14909_),
    .A2(_14917_),
    .B1(_14908_),
    .Y(_14918_));
 sky130_fd_sc_hd__nand2_2 _36967_ (.A(_14918_),
    .B(_14905_),
    .Y(_14919_));
 sky130_fd_sc_hd__nand3_2 _36968_ (.A(_14890_),
    .B(_14886_),
    .C(_14919_),
    .Y(_14920_));
 sky130_fd_sc_hd__nand3_2 _36969_ (.A(_14914_),
    .B(_14916_),
    .C(_14920_),
    .Y(_14921_));
 sky130_fd_sc_hd__a21o_2 _36970_ (.A1(_14648_),
    .A2(_14651_),
    .B1(_14644_),
    .X(_14922_));
 sky130_fd_sc_hd__and4_2 _36971_ (.A(_14095_),
    .B(_10656_),
    .C(_10966_),
    .D(_08910_),
    .X(_14923_));
 sky130_fd_sc_hd__a22o_2 _36972_ (.A1(_10655_),
    .A2(_09994_),
    .B1(_13454_),
    .B2(_14112_),
    .X(_14924_));
 sky130_fd_sc_hd__inv_2 _36973_ (.A(_14924_),
    .Y(_14925_));
 sky130_fd_sc_hd__nor2_2 _36974_ (.A(_14923_),
    .B(_14925_),
    .Y(_14926_));
 sky130_fd_sc_hd__nor2_2 _36975_ (.A(_07718_),
    .B(_10485_),
    .Y(_14927_));
 sky130_fd_sc_hd__inv_2 _36976_ (.A(_14927_),
    .Y(_14928_));
 sky130_fd_sc_hd__nand2_2 _36977_ (.A(_14926_),
    .B(_14928_),
    .Y(_14929_));
 sky130_fd_sc_hd__o21ai_2 _36978_ (.A1(_14923_),
    .A2(_14925_),
    .B1(_14927_),
    .Y(_14930_));
 sky130_fd_sc_hd__nand3b_2 _36979_ (.A_N(_14922_),
    .B(_14929_),
    .C(_14930_),
    .Y(_14931_));
 sky130_fd_sc_hd__nand2_2 _36980_ (.A(_14926_),
    .B(_14927_),
    .Y(_14932_));
 sky130_fd_sc_hd__o21ai_2 _36981_ (.A1(_14923_),
    .A2(_14925_),
    .B1(_14928_),
    .Y(_14933_));
 sky130_fd_sc_hd__nand3_2 _36982_ (.A(_14932_),
    .B(_14922_),
    .C(_14933_),
    .Y(_14934_));
 sky130_fd_sc_hd__and4_2 _36983_ (.A(_19348_),
    .B(_19351_),
    .C(_10055_),
    .D(_08921_),
    .X(_14935_));
 sky130_fd_sc_hd__a22o_2 _36984_ (.A1(_10210_),
    .A2(_09219_),
    .B1(_08816_),
    .B2(_09216_),
    .X(_14936_));
 sky130_fd_sc_hd__inv_2 _36985_ (.A(_14936_),
    .Y(_14937_));
 sky130_fd_sc_hd__a211o_2 _36986_ (.A1(_19353_),
    .A2(_19560_),
    .B1(_14935_),
    .C1(_14937_),
    .X(_14938_));
 sky130_fd_sc_hd__buf_1 _36987_ (.A(_11374_),
    .X(_14939_));
 sky130_fd_sc_hd__nor2_2 _36988_ (.A(_07053_),
    .B(_14939_),
    .Y(_14940_));
 sky130_fd_sc_hd__o21ai_2 _36989_ (.A1(_14935_),
    .A2(_14937_),
    .B1(_14940_),
    .Y(_14941_));
 sky130_fd_sc_hd__nand2_2 _36990_ (.A(_14938_),
    .B(_14941_),
    .Y(_14942_));
 sky130_fd_sc_hd__a21oi_2 _36991_ (.A1(_14931_),
    .A2(_14934_),
    .B1(_14942_),
    .Y(_14943_));
 sky130_fd_sc_hd__and3_2 _36992_ (.A(_14931_),
    .B(_14934_),
    .C(_14942_),
    .X(_14944_));
 sky130_fd_sc_hd__nand2_2 _36993_ (.A(_14581_),
    .B(_14584_),
    .Y(_14945_));
 sky130_fd_sc_hd__nand2_2 _36994_ (.A(_14945_),
    .B(_14578_),
    .Y(_14946_));
 sky130_fd_sc_hd__o21bai_2 _36995_ (.A1(_14943_),
    .A2(_14944_),
    .B1_N(_14946_),
    .Y(_14947_));
 sky130_fd_sc_hd__a21o_2 _36996_ (.A1(_14931_),
    .A2(_14934_),
    .B1(_14942_),
    .X(_14948_));
 sky130_fd_sc_hd__nand3_2 _36997_ (.A(_14931_),
    .B(_14934_),
    .C(_14942_),
    .Y(_14949_));
 sky130_fd_sc_hd__nand3_2 _36998_ (.A(_14948_),
    .B(_14946_),
    .C(_14949_),
    .Y(_14950_));
 sky130_fd_sc_hd__nand2_2 _36999_ (.A(_14664_),
    .B(_14656_),
    .Y(_14951_));
 sky130_fd_sc_hd__nand2_2 _37000_ (.A(_14951_),
    .B(_14653_),
    .Y(_14952_));
 sky130_fd_sc_hd__inv_2 _37001_ (.A(_14952_),
    .Y(_14953_));
 sky130_fd_sc_hd__a21oi_2 _37002_ (.A1(_14947_),
    .A2(_14950_),
    .B1(_14953_),
    .Y(_14954_));
 sky130_fd_sc_hd__nand3_2 _37003_ (.A(_14947_),
    .B(_14950_),
    .C(_14953_),
    .Y(_14955_));
 sky130_fd_sc_hd__inv_2 _37004_ (.A(_14955_),
    .Y(_14956_));
 sky130_fd_sc_hd__o2bb2ai_2 _37005_ (.A1_N(_14913_),
    .A2_N(_14921_),
    .B1(_14954_),
    .B2(_14956_),
    .Y(_14957_));
 sky130_fd_sc_hd__a21oi_2 _37006_ (.A1(_14948_),
    .A2(_14949_),
    .B1(_14946_),
    .Y(_14958_));
 sky130_fd_sc_hd__nand2_2 _37007_ (.A(_14953_),
    .B(_14950_),
    .Y(_14959_));
 sky130_fd_sc_hd__a21o_2 _37008_ (.A1(_14947_),
    .A2(_14950_),
    .B1(_14953_),
    .X(_14960_));
 sky130_fd_sc_hd__o2111ai_2 _37009_ (.A1(_14958_),
    .A2(_14959_),
    .B1(_14960_),
    .C1(_14913_),
    .D1(_14921_),
    .Y(_14961_));
 sky130_fd_sc_hd__nand2_2 _37010_ (.A(_14686_),
    .B(_14636_),
    .Y(_14962_));
 sky130_fd_sc_hd__a21oi_2 _37011_ (.A1(_14957_),
    .A2(_14961_),
    .B1(_14962_),
    .Y(_14963_));
 sky130_fd_sc_hd__inv_2 _37012_ (.A(_14315_),
    .Y(_14964_));
 sky130_fd_sc_hd__and3_2 _37013_ (.A(_14312_),
    .B(_14319_),
    .C(_14322_),
    .X(_14965_));
 sky130_fd_sc_hd__and3_2 _37014_ (.A(_14665_),
    .B(_14669_),
    .C(_14668_),
    .X(_14966_));
 sky130_fd_sc_hd__o22ai_2 _37015_ (.A1(_14964_),
    .A2(_14965_),
    .B1(_14679_),
    .B2(_14966_),
    .Y(_14967_));
 sky130_fd_sc_hd__nand2_2 _37016_ (.A(_14967_),
    .B(_14675_),
    .Y(_14968_));
 sky130_fd_sc_hd__a31oi_2 _37017_ (.A1(_14638_),
    .A2(_14637_),
    .A3(_14641_),
    .B1(_14968_),
    .Y(_14969_));
 sky130_fd_sc_hd__o211a_2 _37018_ (.A1(_14685_),
    .A2(_14969_),
    .B1(_14961_),
    .C1(_14957_),
    .X(_14970_));
 sky130_fd_sc_hd__nand2_2 _37019_ (.A(_09018_),
    .B(_09722_),
    .Y(_14971_));
 sky130_fd_sc_hd__nand2_2 _37020_ (.A(_09019_),
    .B(_11765_),
    .Y(_14972_));
 sky130_fd_sc_hd__nor2_2 _37021_ (.A(_14971_),
    .B(_14972_),
    .Y(_14973_));
 sky130_fd_sc_hd__and2_2 _37022_ (.A(_14971_),
    .B(_14972_),
    .X(_14974_));
 sky130_fd_sc_hd__nor2_2 _37023_ (.A(_11300_),
    .B(_11764_),
    .Y(_14975_));
 sky130_fd_sc_hd__o21bai_2 _37024_ (.A1(_14973_),
    .A2(_14974_),
    .B1_N(_14975_),
    .Y(_14976_));
 sky130_fd_sc_hd__or2_2 _37025_ (.A(_14971_),
    .B(_14972_),
    .X(_14977_));
 sky130_fd_sc_hd__nand2_2 _37026_ (.A(_14971_),
    .B(_14972_),
    .Y(_14978_));
 sky130_fd_sc_hd__nand3_2 _37027_ (.A(_14977_),
    .B(_14975_),
    .C(_14978_),
    .Y(_14979_));
 sky130_fd_sc_hd__nor2_2 _37028_ (.A(_14658_),
    .B(_14659_),
    .Y(_14980_));
 sky130_fd_sc_hd__o2bb2ai_2 _37029_ (.A1_N(_14976_),
    .A2_N(_14979_),
    .B1(_14661_),
    .B2(_14980_),
    .Y(_14981_));
 sky130_fd_sc_hd__a21o_2 _37030_ (.A1(_14658_),
    .A2(_14660_),
    .B1(_14659_),
    .X(_14982_));
 sky130_fd_sc_hd__nand3_2 _37031_ (.A(_14982_),
    .B(_14976_),
    .C(_14979_),
    .Y(_14983_));
 sky130_fd_sc_hd__nand2_2 _37032_ (.A(_14694_),
    .B(_14693_),
    .Y(_14984_));
 sky130_fd_sc_hd__a21oi_2 _37033_ (.A1(_14981_),
    .A2(_14983_),
    .B1(_14984_),
    .Y(_14985_));
 sky130_fd_sc_hd__and3_2 _37034_ (.A(_14981_),
    .B(_14984_),
    .C(_14983_),
    .X(_14986_));
 sky130_fd_sc_hd__a21oi_2 _37035_ (.A1(_14700_),
    .A2(_14702_),
    .B1(_14698_),
    .Y(_14987_));
 sky130_fd_sc_hd__o21bai_2 _37036_ (.A1(_14985_),
    .A2(_14986_),
    .B1_N(_14987_),
    .Y(_14988_));
 sky130_fd_sc_hd__a21o_2 _37037_ (.A1(_14981_),
    .A2(_14983_),
    .B1(_14984_),
    .X(_14989_));
 sky130_fd_sc_hd__nand3_2 _37038_ (.A(_14981_),
    .B(_14984_),
    .C(_14983_),
    .Y(_14990_));
 sky130_fd_sc_hd__nand3_2 _37039_ (.A(_14989_),
    .B(_14990_),
    .C(_14987_),
    .Y(_14991_));
 sky130_fd_sc_hd__nand2_2 _37040_ (.A(_06790_),
    .B(_11427_),
    .Y(_14992_));
 sky130_fd_sc_hd__nand2_2 _37041_ (.A(_14153_),
    .B(_08320_),
    .Y(_14993_));
 sky130_fd_sc_hd__o21ai_2 _37042_ (.A1(_14992_),
    .A2(_14993_),
    .B1(_14712_),
    .Y(_14994_));
 sky130_fd_sc_hd__a21o_2 _37043_ (.A1(_14992_),
    .A2(_14993_),
    .B1(_14994_),
    .X(_14995_));
 sky130_fd_sc_hd__nor2_2 _37044_ (.A(_14992_),
    .B(_14993_),
    .Y(_14996_));
 sky130_fd_sc_hd__and2_2 _37045_ (.A(_14992_),
    .B(_14993_),
    .X(_14997_));
 sky130_fd_sc_hd__o21ai_2 _37046_ (.A1(_14996_),
    .A2(_14997_),
    .B1(_14715_),
    .Y(_14998_));
 sky130_fd_sc_hd__nand2_2 _37047_ (.A(_14995_),
    .B(_14998_),
    .Y(_14999_));
 sky130_fd_sc_hd__a21oi_2 _37048_ (.A1(_14715_),
    .A2(_14710_),
    .B1(_14709_),
    .Y(_15000_));
 sky130_fd_sc_hd__inv_2 _37049_ (.A(_15000_),
    .Y(_15001_));
 sky130_fd_sc_hd__nand2_2 _37050_ (.A(_14999_),
    .B(_15001_),
    .Y(_15002_));
 sky130_fd_sc_hd__nand3_2 _37051_ (.A(_14995_),
    .B(_14998_),
    .C(_15000_),
    .Y(_15003_));
 sky130_fd_sc_hd__a21o_2 _37052_ (.A1(_15002_),
    .A2(_15003_),
    .B1(_14430_),
    .X(_15004_));
 sky130_fd_sc_hd__nand2_2 _37053_ (.A(_15003_),
    .B(_14429_),
    .Y(_15005_));
 sky130_fd_sc_hd__a21o_2 _37054_ (.A1(_15001_),
    .A2(_14999_),
    .B1(_15005_),
    .X(_15006_));
 sky130_fd_sc_hd__nand2_2 _37055_ (.A(_15004_),
    .B(_15006_),
    .Y(_15007_));
 sky130_fd_sc_hd__a21boi_2 _37056_ (.A1(_14988_),
    .A2(_14991_),
    .B1_N(_15007_),
    .Y(_15008_));
 sky130_fd_sc_hd__a21oi_2 _37057_ (.A1(_14989_),
    .A2(_14990_),
    .B1(_14987_),
    .Y(_15009_));
 sky130_fd_sc_hd__and3_2 _37058_ (.A(_14989_),
    .B(_14990_),
    .C(_14987_),
    .X(_15010_));
 sky130_fd_sc_hd__nor3_2 _37059_ (.A(_15007_),
    .B(_15009_),
    .C(_15010_),
    .Y(_15011_));
 sky130_fd_sc_hd__o21ai_2 _37060_ (.A1(_14678_),
    .A2(_14679_),
    .B1(_14671_),
    .Y(_15012_));
 sky130_fd_sc_hd__o21bai_2 _37061_ (.A1(_15008_),
    .A2(_15011_),
    .B1_N(_15012_),
    .Y(_15013_));
 sky130_fd_sc_hd__o21ai_2 _37062_ (.A1(_15009_),
    .A2(_15010_),
    .B1(_15007_),
    .Y(_15014_));
 sky130_fd_sc_hd__nand3b_2 _37063_ (.A_N(_15007_),
    .B(_14988_),
    .C(_14991_),
    .Y(_15015_));
 sky130_fd_sc_hd__nand3_2 _37064_ (.A(_15014_),
    .B(_15012_),
    .C(_15015_),
    .Y(_15016_));
 sky130_fd_sc_hd__nand2_2 _37065_ (.A(_14723_),
    .B(_14730_),
    .Y(_15017_));
 sky130_fd_sc_hd__a21oi_2 _37066_ (.A1(_15013_),
    .A2(_15016_),
    .B1(_15017_),
    .Y(_15018_));
 sky130_fd_sc_hd__nand2_2 _37067_ (.A(_15014_),
    .B(_15012_),
    .Y(_15019_));
 sky130_fd_sc_hd__o211a_2 _37068_ (.A1(_15011_),
    .A2(_15019_),
    .B1(_15017_),
    .C1(_15013_),
    .X(_15020_));
 sky130_fd_sc_hd__nor2_2 _37069_ (.A(_15018_),
    .B(_15020_),
    .Y(_15021_));
 sky130_fd_sc_hd__o21ai_2 _37070_ (.A1(_14963_),
    .A2(_14970_),
    .B1(_15021_),
    .Y(_15022_));
 sky130_fd_sc_hd__nand2_2 _37071_ (.A(_14747_),
    .B(_14744_),
    .Y(_15023_));
 sky130_fd_sc_hd__nand2_2 _37072_ (.A(_15023_),
    .B(_14743_),
    .Y(_15024_));
 sky130_fd_sc_hd__a22oi_2 _37073_ (.A1(_14960_),
    .A2(_14955_),
    .B1(_14921_),
    .B2(_14913_),
    .Y(_15025_));
 sky130_fd_sc_hd__o2111a_2 _37074_ (.A1(_14958_),
    .A2(_14959_),
    .B1(_14960_),
    .C1(_14913_),
    .D1(_14921_),
    .X(_15026_));
 sky130_fd_sc_hd__nor2_2 _37075_ (.A(_14685_),
    .B(_14969_),
    .Y(_15027_));
 sky130_fd_sc_hd__o21ai_2 _37076_ (.A1(_15025_),
    .A2(_15026_),
    .B1(_15027_),
    .Y(_15028_));
 sky130_fd_sc_hd__a21o_2 _37077_ (.A1(_15013_),
    .A2(_15016_),
    .B1(_15017_),
    .X(_15029_));
 sky130_fd_sc_hd__nand3_2 _37078_ (.A(_15013_),
    .B(_15016_),
    .C(_15017_),
    .Y(_15030_));
 sky130_fd_sc_hd__nand2_2 _37079_ (.A(_15029_),
    .B(_15030_),
    .Y(_15031_));
 sky130_fd_sc_hd__nand3_2 _37080_ (.A(_14962_),
    .B(_14961_),
    .C(_14957_),
    .Y(_15032_));
 sky130_fd_sc_hd__nand3_2 _37081_ (.A(_15028_),
    .B(_15031_),
    .C(_15032_),
    .Y(_15033_));
 sky130_fd_sc_hd__nand3_2 _37082_ (.A(_15022_),
    .B(_15024_),
    .C(_15033_),
    .Y(_15034_));
 sky130_fd_sc_hd__o21ai_2 _37083_ (.A1(_14963_),
    .A2(_14970_),
    .B1(_15031_),
    .Y(_15035_));
 sky130_fd_sc_hd__o21ai_2 _37084_ (.A1(_14747_),
    .A2(_14684_),
    .B1(_14744_),
    .Y(_15036_));
 sky130_fd_sc_hd__nand3_2 _37085_ (.A(_15028_),
    .B(_15021_),
    .C(_15032_),
    .Y(_15037_));
 sky130_fd_sc_hd__nand3_2 _37086_ (.A(_15035_),
    .B(_15036_),
    .C(_15037_),
    .Y(_15038_));
 sky130_fd_sc_hd__nand2_2 _37087_ (.A(_14784_),
    .B(_14482_),
    .Y(_15039_));
 sky130_fd_sc_hd__a31oi_2 _37088_ (.A1(_14728_),
    .A2(_14725_),
    .A3(_14731_),
    .B1(_14734_),
    .Y(_15040_));
 sky130_fd_sc_hd__a21oi_2 _37089_ (.A1(_14713_),
    .A2(_14716_),
    .B1(_14717_),
    .Y(_15041_));
 sky130_fd_sc_hd__o21a_2 _37090_ (.A1(_14759_),
    .A2(_15041_),
    .B1(_14719_),
    .X(_15042_));
 sky130_fd_sc_hd__o21ai_2 _37091_ (.A1(_14757_),
    .A2(_14758_),
    .B1(_15042_),
    .Y(_15043_));
 sky130_fd_sc_hd__o21ai_2 _37092_ (.A1(_14759_),
    .A2(_15041_),
    .B1(_14719_),
    .Y(_15044_));
 sky130_fd_sc_hd__nand3_2 _37093_ (.A(_15044_),
    .B(_14766_),
    .C(_14768_),
    .Y(_15045_));
 sky130_fd_sc_hd__a21oi_2 _37094_ (.A1(_14755_),
    .A2(_14217_),
    .B1(_14764_),
    .Y(_15046_));
 sky130_fd_sc_hd__inv_2 _37095_ (.A(_15046_),
    .Y(_15047_));
 sky130_fd_sc_hd__a21oi_2 _37096_ (.A1(_15043_),
    .A2(_15045_),
    .B1(_15047_),
    .Y(_15048_));
 sky130_fd_sc_hd__and3_2 _37097_ (.A(_15043_),
    .B(_15045_),
    .C(_15047_),
    .X(_15049_));
 sky130_fd_sc_hd__nand2_2 _37098_ (.A(_14762_),
    .B(_14771_),
    .Y(_15050_));
 sky130_fd_sc_hd__o21a_2 _37099_ (.A1(_14758_),
    .A2(_14773_),
    .B1(_15050_),
    .X(_15051_));
 sky130_fd_sc_hd__o21ai_2 _37100_ (.A1(_15048_),
    .A2(_15049_),
    .B1(_15051_),
    .Y(_15052_));
 sky130_fd_sc_hd__a21o_2 _37101_ (.A1(_15043_),
    .A2(_15045_),
    .B1(_15047_),
    .X(_15053_));
 sky130_fd_sc_hd__nand2_2 _37102_ (.A(_15050_),
    .B(_14769_),
    .Y(_15054_));
 sky130_fd_sc_hd__nand3_2 _37103_ (.A(_15043_),
    .B(_15045_),
    .C(_15047_),
    .Y(_15055_));
 sky130_fd_sc_hd__nand3_2 _37104_ (.A(_15053_),
    .B(_15054_),
    .C(_15055_),
    .Y(_15056_));
 sky130_fd_sc_hd__a21oi_2 _37105_ (.A1(_15052_),
    .A2(_15056_),
    .B1(_13702_),
    .Y(_15057_));
 sky130_fd_sc_hd__nand2_2 _37106_ (.A(_15053_),
    .B(_15054_),
    .Y(_15058_));
 sky130_fd_sc_hd__o211a_2 _37107_ (.A1(_15049_),
    .A2(_15058_),
    .B1(_13702_),
    .C1(_15052_),
    .X(_15059_));
 sky130_fd_sc_hd__o22ai_2 _37108_ (.A1(_14737_),
    .A2(_15040_),
    .B1(_15057_),
    .B2(_15059_),
    .Y(_15060_));
 sky130_fd_sc_hd__and2_2 _37109_ (.A(_14728_),
    .B(_14731_),
    .X(_15061_));
 sky130_fd_sc_hd__o21ai_2 _37110_ (.A1(_14452_),
    .A2(_14736_),
    .B1(_14745_),
    .Y(_15062_));
 sky130_fd_sc_hd__nand3_2 _37111_ (.A(_15052_),
    .B(_13397_),
    .C(_15056_),
    .Y(_15063_));
 sky130_fd_sc_hd__o2bb2ai_2 _37112_ (.A1_N(_15056_),
    .A2_N(_15052_),
    .B1(_13352_),
    .B2(_13354_),
    .Y(_15064_));
 sky130_fd_sc_hd__o2111ai_2 _37113_ (.A1(_14725_),
    .A2(_15061_),
    .B1(_15062_),
    .C1(_15063_),
    .D1(_15064_),
    .Y(_15065_));
 sky130_fd_sc_hd__a22oi_2 _37114_ (.A1(_15039_),
    .A2(_14778_),
    .B1(_15060_),
    .B2(_15065_),
    .Y(_15066_));
 sky130_fd_sc_hd__inv_2 _37115_ (.A(_14784_),
    .Y(_15067_));
 sky130_fd_sc_hd__and2_2 _37116_ (.A(_14778_),
    .B(_13702_),
    .X(_15068_));
 sky130_fd_sc_hd__o211a_2 _37117_ (.A1(_15067_),
    .A2(_15068_),
    .B1(_15065_),
    .C1(_15060_),
    .X(_15069_));
 sky130_fd_sc_hd__o2bb2ai_2 _37118_ (.A1_N(_15034_),
    .A2_N(_15038_),
    .B1(_15066_),
    .B2(_15069_),
    .Y(_15070_));
 sky130_fd_sc_hd__nor2_2 _37119_ (.A(_15066_),
    .B(_15069_),
    .Y(_15071_));
 sky130_fd_sc_hd__nand3_2 _37120_ (.A(_15034_),
    .B(_15038_),
    .C(_15071_),
    .Y(_15072_));
 sky130_fd_sc_hd__nand3_2 _37121_ (.A(_14852_),
    .B(_15070_),
    .C(_15072_),
    .Y(_15073_));
 sky130_fd_sc_hd__nand2_2 _37122_ (.A(_15034_),
    .B(_15038_),
    .Y(_15074_));
 sky130_fd_sc_hd__nand2_2 _37123_ (.A(_15074_),
    .B(_15071_),
    .Y(_15075_));
 sky130_fd_sc_hd__a21oi_2 _37124_ (.A1(_14740_),
    .A2(_14748_),
    .B1(_14742_),
    .Y(_15076_));
 sky130_fd_sc_hd__a21oi_2 _37125_ (.A1(_14749_),
    .A2(_14801_),
    .B1(_15076_),
    .Y(_15077_));
 sky130_fd_sc_hd__nand3b_2 _37126_ (.A_N(_15071_),
    .B(_15034_),
    .C(_15038_),
    .Y(_15078_));
 sky130_fd_sc_hd__nand3_2 _37127_ (.A(_15075_),
    .B(_15077_),
    .C(_15078_),
    .Y(_15079_));
 sky130_fd_sc_hd__a31o_2 _37128_ (.A1(_14792_),
    .A2(_14790_),
    .A3(_14791_),
    .B1(_14799_),
    .X(_15080_));
 sky130_fd_sc_hd__buf_1 _37129_ (.A(_13735_),
    .X(_15081_));
 sky130_fd_sc_hd__nand2_2 _37130_ (.A(_15080_),
    .B(_15081_),
    .Y(_15082_));
 sky130_fd_sc_hd__inv_2 _37131_ (.A(_15082_),
    .Y(_15083_));
 sky130_fd_sc_hd__nand2_2 _37132_ (.A(_14793_),
    .B(_14017_),
    .Y(_15084_));
 sky130_fd_sc_hd__nor2_2 _37133_ (.A(_15084_),
    .B(_14799_),
    .Y(_15085_));
 sky130_fd_sc_hd__o2bb2ai_2 _37134_ (.A1_N(_15073_),
    .A2_N(_15079_),
    .B1(_15083_),
    .B2(_15085_),
    .Y(_15086_));
 sky130_fd_sc_hd__o21a_2 _37135_ (.A1(_14799_),
    .A2(_15084_),
    .B1(_15082_),
    .X(_15087_));
 sky130_fd_sc_hd__nand3_2 _37136_ (.A(_15079_),
    .B(_15087_),
    .C(_15073_),
    .Y(_15088_));
 sky130_fd_sc_hd__o21ai_2 _37137_ (.A1(_14815_),
    .A2(_14804_),
    .B1(_14820_),
    .Y(_15089_));
 sky130_fd_sc_hd__a21oi_2 _37138_ (.A1(_15086_),
    .A2(_15088_),
    .B1(_15089_),
    .Y(_15090_));
 sky130_fd_sc_hd__a21oi_2 _37139_ (.A1(_15075_),
    .A2(_15078_),
    .B1(_15077_),
    .Y(_15091_));
 sky130_fd_sc_hd__nand2_2 _37140_ (.A(_15079_),
    .B(_15087_),
    .Y(_15092_));
 sky130_fd_sc_hd__o211a_2 _37141_ (.A1(_15091_),
    .A2(_15092_),
    .B1(_15086_),
    .C1(_15089_),
    .X(_15093_));
 sky130_fd_sc_hd__o22ai_2 _37142_ (.A1(_14019_),
    .A2(_14824_),
    .B1(_15090_),
    .B2(_15093_),
    .Y(_15094_));
 sky130_fd_sc_hd__a21o_2 _37143_ (.A1(_15086_),
    .A2(_15088_),
    .B1(_15089_),
    .X(_15095_));
 sky130_fd_sc_hd__nand3_2 _37144_ (.A(_15089_),
    .B(_15086_),
    .C(_15088_),
    .Y(_15096_));
 sky130_fd_sc_hd__nand3_2 _37145_ (.A(_15095_),
    .B(_14825_),
    .C(_15096_),
    .Y(_15097_));
 sky130_fd_sc_hd__inv_2 _37146_ (.A(_14828_),
    .Y(_15098_));
 sky130_fd_sc_hd__nand2_2 _37147_ (.A(_14827_),
    .B(_14829_),
    .Y(_15099_));
 sky130_fd_sc_hd__o2bb2ai_2 _37148_ (.A1_N(_14549_),
    .A2_N(_14822_),
    .B1(_15098_),
    .B2(_15099_),
    .Y(_15100_));
 sky130_fd_sc_hd__a21o_2 _37149_ (.A1(_15094_),
    .A2(_15097_),
    .B1(_15100_),
    .X(_15101_));
 sky130_fd_sc_hd__nand3_2 _37150_ (.A(_15094_),
    .B(_15100_),
    .C(_15097_),
    .Y(_15102_));
 sky130_fd_sc_hd__nand2_2 _37151_ (.A(_15101_),
    .B(_15102_),
    .Y(_15103_));
 sky130_fd_sc_hd__a21oi_2 _37152_ (.A1(_14850_),
    .A2(_14839_),
    .B1(_14836_),
    .Y(_15104_));
 sky130_fd_sc_hd__xor2_2 _37153_ (.A(_15103_),
    .B(_15104_),
    .X(_02664_));
 sky130_fd_sc_hd__o211ai_2 _37154_ (.A1(_15067_),
    .A2(_15068_),
    .B1(_15065_),
    .C1(_15060_),
    .Y(_15105_));
 sky130_fd_sc_hd__nand2_2 _37155_ (.A(_15105_),
    .B(_15065_),
    .Y(_15106_));
 sky130_fd_sc_hd__inv_2 _37156_ (.A(_15106_),
    .Y(_15107_));
 sky130_fd_sc_hd__nor2_2 _37157_ (.A(_14018_),
    .B(_15107_),
    .Y(_15108_));
 sky130_fd_sc_hd__buf_1 _37158_ (.A(_15081_),
    .X(_15109_));
 sky130_fd_sc_hd__nor2_2 _37159_ (.A(_15109_),
    .B(_15106_),
    .Y(_15110_));
 sky130_fd_sc_hd__o21a_2 _37160_ (.A1(_14952_),
    .A2(_14958_),
    .B1(_14950_),
    .X(_15111_));
 sky130_fd_sc_hd__nand2_2 _37161_ (.A(_19355_),
    .B(_10371_),
    .Y(_15112_));
 sky130_fd_sc_hd__nand2_2 _37162_ (.A(_19358_),
    .B(_11038_),
    .Y(_15113_));
 sky130_fd_sc_hd__nand2_2 _37163_ (.A(_15112_),
    .B(_15113_),
    .Y(_15114_));
 sky130_fd_sc_hd__or2_2 _37164_ (.A(_15112_),
    .B(_15113_),
    .X(_15115_));
 sky130_fd_sc_hd__buf_1 _37165_ (.A(_10520_),
    .X(_15116_));
 sky130_fd_sc_hd__o2bb2ai_2 _37166_ (.A1_N(_15114_),
    .A2_N(_15115_),
    .B1(_11300_),
    .B2(_15116_),
    .Y(_15117_));
 sky130_fd_sc_hd__nor2_2 _37167_ (.A(_11300_),
    .B(_10520_),
    .Y(_15118_));
 sky130_fd_sc_hd__nand3_2 _37168_ (.A(_15115_),
    .B(_15118_),
    .C(_15114_),
    .Y(_15119_));
 sky130_fd_sc_hd__a21o_2 _37169_ (.A1(_14940_),
    .A2(_14936_),
    .B1(_14935_),
    .X(_15120_));
 sky130_fd_sc_hd__a21o_2 _37170_ (.A1(_15117_),
    .A2(_15119_),
    .B1(_15120_),
    .X(_15121_));
 sky130_fd_sc_hd__nand3_2 _37171_ (.A(_15117_),
    .B(_15119_),
    .C(_15120_),
    .Y(_15122_));
 sky130_fd_sc_hd__nand2_2 _37172_ (.A(_14979_),
    .B(_14977_),
    .Y(_15123_));
 sky130_fd_sc_hd__a21o_2 _37173_ (.A1(_15121_),
    .A2(_15122_),
    .B1(_15123_),
    .X(_15124_));
 sky130_fd_sc_hd__nand3_2 _37174_ (.A(_15121_),
    .B(_15123_),
    .C(_15122_),
    .Y(_15125_));
 sky130_fd_sc_hd__nand2_2 _37175_ (.A(_14990_),
    .B(_14983_),
    .Y(_15126_));
 sky130_fd_sc_hd__a21oi_2 _37176_ (.A1(_15124_),
    .A2(_15125_),
    .B1(_15126_),
    .Y(_15127_));
 sky130_fd_sc_hd__and3_2 _37177_ (.A(_15124_),
    .B(_15126_),
    .C(_15125_),
    .X(_15128_));
 sky130_fd_sc_hd__o21ai_2 _37178_ (.A1(_06790_),
    .A2(_06115_),
    .B1(_11429_),
    .Y(_15129_));
 sky130_fd_sc_hd__and3_2 _37179_ (.A(_11759_),
    .B(_19362_),
    .C(_07015_),
    .X(_15130_));
 sky130_fd_sc_hd__nor2_2 _37180_ (.A(_15129_),
    .B(_15130_),
    .Y(_15131_));
 sky130_fd_sc_hd__o21ai_2 _37181_ (.A1(_06121_),
    .A2(_14997_),
    .B1(_14994_),
    .Y(_15132_));
 sky130_fd_sc_hd__or2_2 _37182_ (.A(_15131_),
    .B(_15132_),
    .X(_15133_));
 sky130_fd_sc_hd__nand2_2 _37183_ (.A(_15132_),
    .B(_15131_),
    .Y(_15134_));
 sky130_fd_sc_hd__a21oi_2 _37184_ (.A1(_15133_),
    .A2(_15134_),
    .B1(_14759_),
    .Y(_15135_));
 sky130_fd_sc_hd__nand2_2 _37185_ (.A(_15133_),
    .B(_15134_),
    .Y(_15136_));
 sky130_fd_sc_hd__nor2_2 _37186_ (.A(_14430_),
    .B(_15136_),
    .Y(_15137_));
 sky130_fd_sc_hd__nor2_2 _37187_ (.A(_15135_),
    .B(_15137_),
    .Y(_15138_));
 sky130_fd_sc_hd__o21ai_2 _37188_ (.A1(_15127_),
    .A2(_15128_),
    .B1(_15138_),
    .Y(_15139_));
 sky130_fd_sc_hd__inv_2 _37189_ (.A(_15138_),
    .Y(_15140_));
 sky130_fd_sc_hd__a21o_2 _37190_ (.A1(_15124_),
    .A2(_15125_),
    .B1(_15126_),
    .X(_15141_));
 sky130_fd_sc_hd__nand3_2 _37191_ (.A(_15124_),
    .B(_15126_),
    .C(_15125_),
    .Y(_15142_));
 sky130_fd_sc_hd__nand3_2 _37192_ (.A(_15140_),
    .B(_15141_),
    .C(_15142_),
    .Y(_15143_));
 sky130_fd_sc_hd__nand3_2 _37193_ (.A(_15111_),
    .B(_15139_),
    .C(_15143_),
    .Y(_15144_));
 sky130_fd_sc_hd__o21ai_2 _37194_ (.A1(_15127_),
    .A2(_15128_),
    .B1(_15140_),
    .Y(_15145_));
 sky130_fd_sc_hd__o21ai_2 _37195_ (.A1(_14952_),
    .A2(_14958_),
    .B1(_14950_),
    .Y(_15146_));
 sky130_fd_sc_hd__nand3_2 _37196_ (.A(_15141_),
    .B(_15138_),
    .C(_15142_),
    .Y(_15147_));
 sky130_fd_sc_hd__nand3_2 _37197_ (.A(_15145_),
    .B(_15146_),
    .C(_15147_),
    .Y(_15148_));
 sky130_fd_sc_hd__nand2_2 _37198_ (.A(_15144_),
    .B(_15148_),
    .Y(_15149_));
 sky130_fd_sc_hd__nand2_2 _37199_ (.A(_15015_),
    .B(_14991_),
    .Y(_15150_));
 sky130_fd_sc_hd__inv_2 _37200_ (.A(_15150_),
    .Y(_15151_));
 sky130_fd_sc_hd__and2_2 _37201_ (.A(_15149_),
    .B(_15151_),
    .X(_15152_));
 sky130_fd_sc_hd__nand3_2 _37202_ (.A(_15144_),
    .B(_15148_),
    .C(_15150_),
    .Y(_15153_));
 sky130_fd_sc_hd__inv_2 _37203_ (.A(_15153_),
    .Y(_15154_));
 sky130_fd_sc_hd__nand2_2 _37204_ (.A(_10193_),
    .B(_14112_),
    .Y(_15155_));
 sky130_fd_sc_hd__nand2_2 _37205_ (.A(_08799_),
    .B(_08662_),
    .Y(_15156_));
 sky130_fd_sc_hd__nor2_2 _37206_ (.A(_15155_),
    .B(_15156_),
    .Y(_15157_));
 sky130_fd_sc_hd__and2_2 _37207_ (.A(_15155_),
    .B(_15156_),
    .X(_15158_));
 sky130_fd_sc_hd__buf_1 _37208_ (.A(_11671_),
    .X(_15159_));
 sky130_fd_sc_hd__nor2_2 _37209_ (.A(_07718_),
    .B(_15159_),
    .Y(_15160_));
 sky130_fd_sc_hd__o21bai_2 _37210_ (.A1(_15157_),
    .A2(_15158_),
    .B1_N(_15160_),
    .Y(_15161_));
 sky130_fd_sc_hd__nand2_2 _37211_ (.A(_15155_),
    .B(_15156_),
    .Y(_15162_));
 sky130_fd_sc_hd__nand3b_2 _37212_ (.A_N(_15157_),
    .B(_15160_),
    .C(_15162_),
    .Y(_15163_));
 sky130_fd_sc_hd__nand2_2 _37213_ (.A(_15161_),
    .B(_15163_),
    .Y(_15164_));
 sky130_fd_sc_hd__a21oi_2 _37214_ (.A1(_14927_),
    .A2(_14924_),
    .B1(_14923_),
    .Y(_15165_));
 sky130_fd_sc_hd__nand2_2 _37215_ (.A(_15164_),
    .B(_15165_),
    .Y(_15166_));
 sky130_fd_sc_hd__a21o_2 _37216_ (.A1(_14927_),
    .A2(_14924_),
    .B1(_14923_),
    .X(_15167_));
 sky130_fd_sc_hd__nand3_2 _37217_ (.A(_15167_),
    .B(_15161_),
    .C(_15163_),
    .Y(_15168_));
 sky130_fd_sc_hd__and4_2 _37218_ (.A(_19348_),
    .B(_19351_),
    .C(_09733_),
    .D(_09216_),
    .X(_15169_));
 sky130_fd_sc_hd__o22a_2 _37219_ (.A1(_12596_),
    .A2(_10523_),
    .B1(_12597_),
    .B2(_13274_),
    .X(_15170_));
 sky130_fd_sc_hd__nor2_2 _37220_ (.A(_07053_),
    .B(_10543_),
    .Y(_15171_));
 sky130_fd_sc_hd__o21ai_2 _37221_ (.A1(_15169_),
    .A2(_15170_),
    .B1(_15171_),
    .Y(_15172_));
 sky130_fd_sc_hd__inv_2 _37222_ (.A(_15171_),
    .Y(_15173_));
 sky130_fd_sc_hd__a22o_2 _37223_ (.A1(_19348_),
    .A2(_10055_),
    .B1(_19351_),
    .B2(_19559_),
    .X(_15174_));
 sky130_fd_sc_hd__nand3b_2 _37224_ (.A_N(_15169_),
    .B(_15173_),
    .C(_15174_),
    .Y(_15175_));
 sky130_fd_sc_hd__nand2_2 _37225_ (.A(_15172_),
    .B(_15175_),
    .Y(_15176_));
 sky130_fd_sc_hd__a21oi_2 _37226_ (.A1(_15166_),
    .A2(_15168_),
    .B1(_15176_),
    .Y(_15177_));
 sky130_fd_sc_hd__and3_2 _37227_ (.A(_15166_),
    .B(_15168_),
    .C(_15176_),
    .X(_15178_));
 sky130_fd_sc_hd__a21oi_2 _37228_ (.A1(_14900_),
    .A2(_14903_),
    .B1(_14917_),
    .Y(_15179_));
 sky130_fd_sc_hd__o21ai_2 _37229_ (.A1(_15177_),
    .A2(_15178_),
    .B1(_15179_),
    .Y(_15180_));
 sky130_fd_sc_hd__a21o_2 _37230_ (.A1(_15166_),
    .A2(_15168_),
    .B1(_15176_),
    .X(_15181_));
 sky130_fd_sc_hd__o21ai_2 _37231_ (.A1(_14908_),
    .A2(_14909_),
    .B1(_14901_),
    .Y(_15182_));
 sky130_fd_sc_hd__nand3_2 _37232_ (.A(_15166_),
    .B(_15168_),
    .C(_15176_),
    .Y(_15183_));
 sky130_fd_sc_hd__nand3_2 _37233_ (.A(_15181_),
    .B(_15182_),
    .C(_15183_),
    .Y(_15184_));
 sky130_fd_sc_hd__a21boi_2 _37234_ (.A1(_14931_),
    .A2(_14942_),
    .B1_N(_14934_),
    .Y(_15185_));
 sky130_fd_sc_hd__a21boi_2 _37235_ (.A1(_15180_),
    .A2(_15184_),
    .B1_N(_15185_),
    .Y(_15186_));
 sky130_fd_sc_hd__nand2_2 _37236_ (.A(_15181_),
    .B(_15183_),
    .Y(_15187_));
 sky130_fd_sc_hd__a21oi_2 _37237_ (.A1(_15187_),
    .A2(_15179_),
    .B1(_15185_),
    .Y(_15188_));
 sky130_fd_sc_hd__and2_2 _37238_ (.A(_15188_),
    .B(_15184_),
    .X(_15189_));
 sky130_fd_sc_hd__nor2_2 _37239_ (.A(_14339_),
    .B(_14646_),
    .Y(_15190_));
 sky130_fd_sc_hd__nand2_2 _37240_ (.A(_09819_),
    .B(_07358_),
    .Y(_15191_));
 sky130_fd_sc_hd__a21o_2 _37241_ (.A1(_10156_),
    .A2(_08651_),
    .B1(_15191_),
    .X(_15192_));
 sky130_fd_sc_hd__nand2_2 _37242_ (.A(_10158_),
    .B(_19577_),
    .Y(_15193_));
 sky130_fd_sc_hd__a21o_2 _37243_ (.A1(_19328_),
    .A2(_19580_),
    .B1(_15193_),
    .X(_15194_));
 sky130_fd_sc_hd__nand3b_2 _37244_ (.A_N(_15190_),
    .B(_15192_),
    .C(_15194_),
    .Y(_15195_));
 sky130_fd_sc_hd__nand2_2 _37245_ (.A(_15192_),
    .B(_15194_),
    .Y(_15196_));
 sky130_fd_sc_hd__nand2_2 _37246_ (.A(_15196_),
    .B(_15190_),
    .Y(_15197_));
 sky130_fd_sc_hd__nor2_2 _37247_ (.A(_14872_),
    .B(_14867_),
    .Y(_15198_));
 sky130_fd_sc_hd__nor2_2 _37248_ (.A(_14870_),
    .B(_15198_),
    .Y(_15199_));
 sky130_fd_sc_hd__a21o_2 _37249_ (.A1(_15195_),
    .A2(_15197_),
    .B1(_15199_),
    .X(_15200_));
 sky130_fd_sc_hd__nand3_2 _37250_ (.A(_15199_),
    .B(_15195_),
    .C(_15197_),
    .Y(_15201_));
 sky130_fd_sc_hd__nand2_2 _37251_ (.A(_14897_),
    .B(_14894_),
    .Y(_15202_));
 sky130_fd_sc_hd__a21oi_2 _37252_ (.A1(_15200_),
    .A2(_15201_),
    .B1(_15202_),
    .Y(_15203_));
 sky130_fd_sc_hd__nand3_2 _37253_ (.A(_15200_),
    .B(_15202_),
    .C(_15201_),
    .Y(_15204_));
 sky130_fd_sc_hd__inv_2 _37254_ (.A(_15204_),
    .Y(_15205_));
 sky130_fd_sc_hd__nand3_2 _37255_ (.A(_11169_),
    .B(_13146_),
    .C(_19594_),
    .Y(_15206_));
 sky130_fd_sc_hd__nor2_2 _37256_ (.A(_06388_),
    .B(_15206_),
    .Y(_15207_));
 sky130_fd_sc_hd__o22a_2 _37257_ (.A1(_06388_),
    .A2(_18182_),
    .B1(_14855_),
    .B2(_06958_),
    .X(_15208_));
 sky130_fd_sc_hd__nor2_2 _37258_ (.A(_10150_),
    .B(_08053_),
    .Y(_15209_));
 sky130_fd_sc_hd__o21bai_2 _37259_ (.A1(_15207_),
    .A2(_15208_),
    .B1_N(_15209_),
    .Y(_15210_));
 sky130_fd_sc_hd__a22o_2 _37260_ (.A1(_19308_),
    .A2(_06557_),
    .B1(_06396_),
    .B2(_14356_),
    .X(_15211_));
 sky130_fd_sc_hd__nand3b_2 _37261_ (.A_N(_15207_),
    .B(_15211_),
    .C(_15209_),
    .Y(_15212_));
 sky130_fd_sc_hd__o21ai_2 _37262_ (.A1(_14857_),
    .A2(_14856_),
    .B1(_14861_),
    .Y(_15213_));
 sky130_fd_sc_hd__a21oi_2 _37263_ (.A1(_15210_),
    .A2(_15212_),
    .B1(_15213_),
    .Y(_15214_));
 sky130_fd_sc_hd__and3_2 _37264_ (.A(_15213_),
    .B(_15210_),
    .C(_15212_),
    .X(_15215_));
 sky130_fd_sc_hd__nor2_2 _37265_ (.A(_09357_),
    .B(_08947_),
    .Y(_15216_));
 sky130_fd_sc_hd__and4_2 _37266_ (.A(_19316_),
    .B(_10136_),
    .C(_07153_),
    .D(_06945_),
    .X(_15217_));
 sky130_fd_sc_hd__nand2_2 _37267_ (.A(_19316_),
    .B(_06945_),
    .Y(_15218_));
 sky130_fd_sc_hd__o21a_2 _37268_ (.A1(_14868_),
    .A2(_08604_),
    .B1(_15218_),
    .X(_15219_));
 sky130_fd_sc_hd__nor3_2 _37269_ (.A(_15216_),
    .B(_15217_),
    .C(_15219_),
    .Y(_15220_));
 sky130_fd_sc_hd__o21a_2 _37270_ (.A1(_15217_),
    .A2(_15219_),
    .B1(_15216_),
    .X(_15221_));
 sky130_fd_sc_hd__nor2_2 _37271_ (.A(_15220_),
    .B(_15221_),
    .Y(_15222_));
 sky130_fd_sc_hd__o21ai_2 _37272_ (.A1(_15214_),
    .A2(_15215_),
    .B1(_15222_),
    .Y(_15223_));
 sky130_fd_sc_hd__a21o_2 _37273_ (.A1(_15210_),
    .A2(_15212_),
    .B1(_15213_),
    .X(_15224_));
 sky130_fd_sc_hd__o21ai_2 _37274_ (.A1(_15217_),
    .A2(_15219_),
    .B1(_15216_),
    .Y(_15225_));
 sky130_fd_sc_hd__or2b_2 _37275_ (.A(_15220_),
    .B_N(_15225_),
    .X(_15226_));
 sky130_fd_sc_hd__nand3_2 _37276_ (.A(_15213_),
    .B(_15210_),
    .C(_15212_),
    .Y(_15227_));
 sky130_fd_sc_hd__nand3_2 _37277_ (.A(_15224_),
    .B(_15226_),
    .C(_15227_),
    .Y(_15228_));
 sky130_fd_sc_hd__o21ai_2 _37278_ (.A1(_14876_),
    .A2(_14865_),
    .B1(_14881_),
    .Y(_15229_));
 sky130_fd_sc_hd__a21oi_2 _37279_ (.A1(_15223_),
    .A2(_15228_),
    .B1(_15229_),
    .Y(_15230_));
 sky130_fd_sc_hd__nand2_2 _37280_ (.A(_15224_),
    .B(_15226_),
    .Y(_15231_));
 sky130_fd_sc_hd__o211a_2 _37281_ (.A1(_15215_),
    .A2(_15231_),
    .B1(_15229_),
    .C1(_15223_),
    .X(_15232_));
 sky130_fd_sc_hd__o22ai_2 _37282_ (.A1(_15203_),
    .A2(_15205_),
    .B1(_15230_),
    .B2(_15232_),
    .Y(_15233_));
 sky130_fd_sc_hd__a21o_2 _37283_ (.A1(_15223_),
    .A2(_15228_),
    .B1(_15229_),
    .X(_15234_));
 sky130_fd_sc_hd__nor2_2 _37284_ (.A(_15203_),
    .B(_15205_),
    .Y(_15235_));
 sky130_fd_sc_hd__nand3_2 _37285_ (.A(_15223_),
    .B(_15229_),
    .C(_15228_),
    .Y(_15236_));
 sky130_fd_sc_hd__nand3_2 _37286_ (.A(_15234_),
    .B(_15235_),
    .C(_15236_),
    .Y(_15237_));
 sky130_fd_sc_hd__nand2_2 _37287_ (.A(_14911_),
    .B(_14890_),
    .Y(_15238_));
 sky130_fd_sc_hd__nand2_2 _37288_ (.A(_15238_),
    .B(_14886_),
    .Y(_15239_));
 sky130_fd_sc_hd__a21oi_2 _37289_ (.A1(_15233_),
    .A2(_15237_),
    .B1(_15239_),
    .Y(_15240_));
 sky130_fd_sc_hd__inv_2 _37290_ (.A(_14886_),
    .Y(_15241_));
 sky130_fd_sc_hd__a31oi_2 _37291_ (.A1(_14887_),
    .A2(_14889_),
    .A3(_14888_),
    .B1(_14919_),
    .Y(_15242_));
 sky130_fd_sc_hd__o211a_2 _37292_ (.A1(_15241_),
    .A2(_15242_),
    .B1(_15237_),
    .C1(_15233_),
    .X(_15243_));
 sky130_fd_sc_hd__o22ai_2 _37293_ (.A1(_15186_),
    .A2(_15189_),
    .B1(_15240_),
    .B2(_15243_),
    .Y(_15244_));
 sky130_fd_sc_hd__a21o_2 _37294_ (.A1(_15233_),
    .A2(_15237_),
    .B1(_15239_),
    .X(_15245_));
 sky130_fd_sc_hd__a21oi_2 _37295_ (.A1(_15184_),
    .A2(_15188_),
    .B1(_15186_),
    .Y(_15246_));
 sky130_fd_sc_hd__nand3_2 _37296_ (.A(_15233_),
    .B(_15239_),
    .C(_15237_),
    .Y(_15247_));
 sky130_fd_sc_hd__nand3_2 _37297_ (.A(_15245_),
    .B(_15246_),
    .C(_15247_),
    .Y(_15248_));
 sky130_fd_sc_hd__a21oi_2 _37298_ (.A1(_14907_),
    .A2(_14912_),
    .B1(_14853_),
    .Y(_15249_));
 sky130_fd_sc_hd__nand2_2 _37299_ (.A(_14960_),
    .B(_14955_),
    .Y(_15250_));
 sky130_fd_sc_hd__o21ai_2 _37300_ (.A1(_15249_),
    .A2(_15250_),
    .B1(_14913_),
    .Y(_15251_));
 sky130_fd_sc_hd__a21oi_2 _37301_ (.A1(_15244_),
    .A2(_15248_),
    .B1(_15251_),
    .Y(_15252_));
 sky130_fd_sc_hd__nand2_2 _37302_ (.A(_15247_),
    .B(_15246_),
    .Y(_15253_));
 sky130_fd_sc_hd__o211a_2 _37303_ (.A1(_15240_),
    .A2(_15253_),
    .B1(_15251_),
    .C1(_15244_),
    .X(_15254_));
 sky130_fd_sc_hd__o22ai_2 _37304_ (.A1(_15152_),
    .A2(_15154_),
    .B1(_15252_),
    .B2(_15254_),
    .Y(_15255_));
 sky130_fd_sc_hd__nand2_2 _37305_ (.A(_15149_),
    .B(_15151_),
    .Y(_15256_));
 sky130_fd_sc_hd__nand2_2 _37306_ (.A(_15256_),
    .B(_15153_),
    .Y(_15257_));
 sky130_fd_sc_hd__nor2_2 _37307_ (.A(_15240_),
    .B(_15253_),
    .Y(_15258_));
 sky130_fd_sc_hd__a21oi_2 _37308_ (.A1(_15245_),
    .A2(_15247_),
    .B1(_15246_),
    .Y(_15259_));
 sky130_fd_sc_hd__o21bai_2 _37309_ (.A1(_15258_),
    .A2(_15259_),
    .B1_N(_15251_),
    .Y(_15260_));
 sky130_fd_sc_hd__nand3_2 _37310_ (.A(_15244_),
    .B(_15251_),
    .C(_15248_),
    .Y(_15261_));
 sky130_fd_sc_hd__nand3b_2 _37311_ (.A_N(_15257_),
    .B(_15260_),
    .C(_15261_),
    .Y(_15262_));
 sky130_fd_sc_hd__o21ai_2 _37312_ (.A1(_15031_),
    .A2(_14963_),
    .B1(_15032_),
    .Y(_15263_));
 sky130_fd_sc_hd__nand3_2 _37313_ (.A(_15255_),
    .B(_15262_),
    .C(_15263_),
    .Y(_15264_));
 sky130_fd_sc_hd__o21bai_2 _37314_ (.A1(_15252_),
    .A2(_15254_),
    .B1_N(_15257_),
    .Y(_15265_));
 sky130_fd_sc_hd__a21oi_2 _37315_ (.A1(_15028_),
    .A2(_15021_),
    .B1(_14970_),
    .Y(_15266_));
 sky130_fd_sc_hd__nand3_2 _37316_ (.A(_15260_),
    .B(_15261_),
    .C(_15257_),
    .Y(_15267_));
 sky130_fd_sc_hd__nand3_2 _37317_ (.A(_15265_),
    .B(_15266_),
    .C(_15267_),
    .Y(_15268_));
 sky130_fd_sc_hd__inv_2 _37318_ (.A(_15017_),
    .Y(_15269_));
 sky130_fd_sc_hd__a21oi_2 _37319_ (.A1(_15014_),
    .A2(_15015_),
    .B1(_15012_),
    .Y(_15270_));
 sky130_fd_sc_hd__o21a_2 _37320_ (.A1(_15269_),
    .A2(_15270_),
    .B1(_15016_),
    .X(_15271_));
 sky130_fd_sc_hd__nand2_2 _37321_ (.A(_15005_),
    .B(_15002_),
    .Y(_15272_));
 sky130_fd_sc_hd__a21o_2 _37322_ (.A1(_14766_),
    .A2(_14768_),
    .B1(_15272_),
    .X(_15273_));
 sky130_fd_sc_hd__nand3_2 _37323_ (.A(_14766_),
    .B(_15272_),
    .C(_14768_),
    .Y(_15274_));
 sky130_fd_sc_hd__a21oi_2 _37324_ (.A1(_15273_),
    .A2(_15274_),
    .B1(_15047_),
    .Y(_15275_));
 sky130_fd_sc_hd__nand2_2 _37325_ (.A(_15273_),
    .B(_15274_),
    .Y(_15276_));
 sky130_fd_sc_hd__nor2_2 _37326_ (.A(_15046_),
    .B(_15276_),
    .Y(_15277_));
 sky130_fd_sc_hd__nand2_2 _37327_ (.A(_15055_),
    .B(_15045_),
    .Y(_15278_));
 sky130_fd_sc_hd__o21bai_2 _37328_ (.A1(_15275_),
    .A2(_15277_),
    .B1_N(_15278_),
    .Y(_15279_));
 sky130_fd_sc_hd__nand2_2 _37329_ (.A(_15276_),
    .B(_15046_),
    .Y(_15280_));
 sky130_fd_sc_hd__nand3_2 _37330_ (.A(_15273_),
    .B(_15047_),
    .C(_15274_),
    .Y(_15281_));
 sky130_fd_sc_hd__nand3_2 _37331_ (.A(_15280_),
    .B(_15278_),
    .C(_15281_),
    .Y(_15282_));
 sky130_fd_sc_hd__nand2_2 _37332_ (.A(_15279_),
    .B(_15282_),
    .Y(_15283_));
 sky130_fd_sc_hd__nand2_2 _37333_ (.A(_15283_),
    .B(_14794_),
    .Y(_15284_));
 sky130_fd_sc_hd__nand3_2 _37334_ (.A(_15279_),
    .B(_14482_),
    .C(_15282_),
    .Y(_15285_));
 sky130_fd_sc_hd__nand3_2 _37335_ (.A(_15271_),
    .B(_15284_),
    .C(_15285_),
    .Y(_15286_));
 sky130_fd_sc_hd__nand2_2 _37336_ (.A(_15283_),
    .B(_14482_),
    .Y(_15287_));
 sky130_fd_sc_hd__o21ai_2 _37337_ (.A1(_15269_),
    .A2(_15270_),
    .B1(_15016_),
    .Y(_15288_));
 sky130_fd_sc_hd__nand3_2 _37338_ (.A(_15279_),
    .B(_14794_),
    .C(_15282_),
    .Y(_15289_));
 sky130_fd_sc_hd__nand3_2 _37339_ (.A(_15287_),
    .B(_15288_),
    .C(_15289_),
    .Y(_15290_));
 sky130_fd_sc_hd__nand2_2 _37340_ (.A(_15063_),
    .B(_15056_),
    .Y(_15291_));
 sky130_fd_sc_hd__a21oi_2 _37341_ (.A1(_15286_),
    .A2(_15290_),
    .B1(_15291_),
    .Y(_15292_));
 sky130_fd_sc_hd__and3_2 _37342_ (.A(_15286_),
    .B(_15290_),
    .C(_15291_),
    .X(_15293_));
 sky130_fd_sc_hd__o2bb2ai_2 _37343_ (.A1_N(_15264_),
    .A2_N(_15268_),
    .B1(_15292_),
    .B2(_15293_),
    .Y(_15294_));
 sky130_fd_sc_hd__inv_2 _37344_ (.A(_15291_),
    .Y(_15295_));
 sky130_fd_sc_hd__a31oi_2 _37345_ (.A1(_15284_),
    .A2(_15271_),
    .A3(_15285_),
    .B1(_15295_),
    .Y(_15296_));
 sky130_fd_sc_hd__a21oi_2 _37346_ (.A1(_15290_),
    .A2(_15296_),
    .B1(_15292_),
    .Y(_15297_));
 sky130_fd_sc_hd__nand3_2 _37347_ (.A(_15268_),
    .B(_15264_),
    .C(_15297_),
    .Y(_15298_));
 sky130_fd_sc_hd__inv_2 _37348_ (.A(_15037_),
    .Y(_15299_));
 sky130_fd_sc_hd__nand2_2 _37349_ (.A(_15035_),
    .B(_15036_),
    .Y(_15300_));
 sky130_fd_sc_hd__o2bb2ai_2 _37350_ (.A1_N(_15071_),
    .A2_N(_15034_),
    .B1(_15299_),
    .B2(_15300_),
    .Y(_15301_));
 sky130_fd_sc_hd__a21oi_2 _37351_ (.A1(_15294_),
    .A2(_15298_),
    .B1(_15301_),
    .Y(_15302_));
 sky130_fd_sc_hd__a21oi_2 _37352_ (.A1(_15268_),
    .A2(_15264_),
    .B1(_15297_),
    .Y(_15303_));
 sky130_fd_sc_hd__nand2_2 _37353_ (.A(_15301_),
    .B(_15298_),
    .Y(_15304_));
 sky130_fd_sc_hd__nor2_2 _37354_ (.A(_15303_),
    .B(_15304_),
    .Y(_15305_));
 sky130_fd_sc_hd__o22ai_2 _37355_ (.A1(_15108_),
    .A2(_15110_),
    .B1(_15302_),
    .B2(_15305_),
    .Y(_15306_));
 sky130_fd_sc_hd__a21o_2 _37356_ (.A1(_15294_),
    .A2(_15298_),
    .B1(_15301_),
    .X(_15307_));
 sky130_fd_sc_hd__nor2_2 _37357_ (.A(_13725_),
    .B(_15106_),
    .Y(_15308_));
 sky130_fd_sc_hd__nor2_2 _37358_ (.A(_13735_),
    .B(_15107_),
    .Y(_15309_));
 sky130_fd_sc_hd__nor2_2 _37359_ (.A(_15308_),
    .B(_15309_),
    .Y(_15310_));
 sky130_fd_sc_hd__inv_2 _37360_ (.A(_15310_),
    .Y(_15311_));
 sky130_fd_sc_hd__nand3_2 _37361_ (.A(_15294_),
    .B(_15298_),
    .C(_15301_),
    .Y(_15312_));
 sky130_fd_sc_hd__nand3_2 _37362_ (.A(_15307_),
    .B(_15311_),
    .C(_15312_),
    .Y(_15313_));
 sky130_fd_sc_hd__nand2_2 _37363_ (.A(_15092_),
    .B(_15073_),
    .Y(_15314_));
 sky130_fd_sc_hd__nand3_2 _37364_ (.A(_15306_),
    .B(_15313_),
    .C(_15314_),
    .Y(_15315_));
 sky130_fd_sc_hd__o22ai_2 _37365_ (.A1(_15309_),
    .A2(_15308_),
    .B1(_15302_),
    .B2(_15305_),
    .Y(_15316_));
 sky130_fd_sc_hd__nand3_2 _37366_ (.A(_15307_),
    .B(_15312_),
    .C(_15310_),
    .Y(_15317_));
 sky130_fd_sc_hd__a21oi_2 _37367_ (.A1(_15087_),
    .A2(_15079_),
    .B1(_15091_),
    .Y(_15318_));
 sky130_fd_sc_hd__nand3_2 _37368_ (.A(_15316_),
    .B(_15317_),
    .C(_15318_),
    .Y(_15319_));
 sky130_fd_sc_hd__buf_1 _37369_ (.A(_14019_),
    .X(_15320_));
 sky130_fd_sc_hd__inv_2 _37370_ (.A(_15080_),
    .Y(_15321_));
 sky130_fd_sc_hd__o2bb2ai_2 _37371_ (.A1_N(_15315_),
    .A2_N(_15319_),
    .B1(_15320_),
    .B2(_15321_),
    .Y(_15322_));
 sky130_fd_sc_hd__nand3_2 _37372_ (.A(_15319_),
    .B(_15315_),
    .C(_15083_),
    .Y(_15323_));
 sky130_fd_sc_hd__inv_2 _37373_ (.A(_14825_),
    .Y(_15324_));
 sky130_fd_sc_hd__o21ai_2 _37374_ (.A1(_15324_),
    .A2(_15090_),
    .B1(_15096_),
    .Y(_15325_));
 sky130_fd_sc_hd__a21o_2 _37375_ (.A1(_15322_),
    .A2(_15323_),
    .B1(_15325_),
    .X(_15326_));
 sky130_fd_sc_hd__nand3_2 _37376_ (.A(_15322_),
    .B(_15325_),
    .C(_15323_),
    .Y(_15327_));
 sky130_fd_sc_hd__and2_2 _37377_ (.A(_15326_),
    .B(_15327_),
    .X(_15328_));
 sky130_fd_sc_hd__inv_2 _37378_ (.A(_15328_),
    .Y(_15329_));
 sky130_fd_sc_hd__and3_2 _37379_ (.A(_15095_),
    .B(_14825_),
    .C(_15096_),
    .X(_15330_));
 sky130_fd_sc_hd__nand2_2 _37380_ (.A(_15094_),
    .B(_15100_),
    .Y(_15331_));
 sky130_fd_sc_hd__o2111ai_2 _37381_ (.A1(_15330_),
    .A2(_15331_),
    .B1(_14835_),
    .C1(_14839_),
    .D1(_15101_),
    .Y(_15332_));
 sky130_fd_sc_hd__inv_2 _37382_ (.A(_15332_),
    .Y(_15333_));
 sky130_fd_sc_hd__nand2_2 _37383_ (.A(_14835_),
    .B(_15102_),
    .Y(_15334_));
 sky130_fd_sc_hd__nand2_2 _37384_ (.A(_15334_),
    .B(_15101_),
    .Y(_15335_));
 sky130_fd_sc_hd__a21boi_2 _37385_ (.A1(_14850_),
    .A2(_15333_),
    .B1_N(_15335_),
    .Y(_15336_));
 sky130_fd_sc_hd__xor2_2 _37386_ (.A(_15329_),
    .B(_15336_),
    .X(_02665_));
 sky130_fd_sc_hd__nand3_2 _37387_ (.A(_10818_),
    .B(_10699_),
    .C(_06946_),
    .Y(_15337_));
 sky130_fd_sc_hd__nor2_2 _37388_ (.A(_06557_),
    .B(_15337_),
    .Y(_15338_));
 sky130_fd_sc_hd__o22a_2 _37389_ (.A1(_06954_),
    .A2(_10830_),
    .B1(_10832_),
    .B2(_08053_),
    .X(_15339_));
 sky130_fd_sc_hd__nand2_2 _37390_ (.A(_19311_),
    .B(_08447_),
    .Y(_15340_));
 sky130_fd_sc_hd__o21ai_2 _37391_ (.A1(_15338_),
    .A2(_15339_),
    .B1(_15340_),
    .Y(_15341_));
 sky130_fd_sc_hd__o2bb2ai_2 _37392_ (.A1_N(_15209_),
    .A2_N(_15211_),
    .B1(_19598_),
    .B2(_15206_),
    .Y(_15342_));
 sky130_fd_sc_hd__a22o_2 _37393_ (.A1(_19308_),
    .A2(_06750_),
    .B1(_06958_),
    .B2(_14356_),
    .X(_15343_));
 sky130_fd_sc_hd__inv_2 _37394_ (.A(_15340_),
    .Y(_15344_));
 sky130_fd_sc_hd__nand3b_2 _37395_ (.A_N(_15338_),
    .B(_15343_),
    .C(_15344_),
    .Y(_15345_));
 sky130_fd_sc_hd__nand3_2 _37396_ (.A(_15341_),
    .B(_15342_),
    .C(_15345_),
    .Y(_15346_));
 sky130_fd_sc_hd__o21ai_2 _37397_ (.A1(_15338_),
    .A2(_15339_),
    .B1(_15344_),
    .Y(_15347_));
 sky130_fd_sc_hd__a21oi_2 _37398_ (.A1(_15211_),
    .A2(_15209_),
    .B1(_15207_),
    .Y(_15348_));
 sky130_fd_sc_hd__nand3b_2 _37399_ (.A_N(_15338_),
    .B(_15343_),
    .C(_15340_),
    .Y(_15349_));
 sky130_fd_sc_hd__nand3_2 _37400_ (.A(_15347_),
    .B(_15348_),
    .C(_15349_),
    .Y(_15350_));
 sky130_fd_sc_hd__a22oi_2 _37401_ (.A1(_10146_),
    .A2(_07153_),
    .B1(_09838_),
    .B2(_08490_),
    .Y(_15351_));
 sky130_fd_sc_hd__nor2_2 _37402_ (.A(_09357_),
    .B(_09246_),
    .Y(_15352_));
 sky130_fd_sc_hd__and4_2 _37403_ (.A(_09842_),
    .B(_10136_),
    .C(_09248_),
    .D(_19585_),
    .X(_15353_));
 sky130_fd_sc_hd__nor3_2 _37404_ (.A(_15351_),
    .B(_15352_),
    .C(_15353_),
    .Y(_15354_));
 sky130_fd_sc_hd__o21ai_2 _37405_ (.A1(_15351_),
    .A2(_15353_),
    .B1(_15352_),
    .Y(_15355_));
 sky130_fd_sc_hd__or2b_2 _37406_ (.A(_15354_),
    .B_N(_15355_),
    .X(_15356_));
 sky130_fd_sc_hd__a21oi_2 _37407_ (.A1(_15346_),
    .A2(_15350_),
    .B1(_15356_),
    .Y(_15357_));
 sky130_fd_sc_hd__inv_2 _37408_ (.A(_15355_),
    .Y(_15358_));
 sky130_fd_sc_hd__o211a_2 _37409_ (.A1(_15354_),
    .A2(_15358_),
    .B1(_15350_),
    .C1(_15346_),
    .X(_15359_));
 sky130_fd_sc_hd__o21a_2 _37410_ (.A1(_15222_),
    .A2(_15214_),
    .B1(_15227_),
    .X(_15360_));
 sky130_fd_sc_hd__o21ai_2 _37411_ (.A1(_15357_),
    .A2(_15359_),
    .B1(_15360_),
    .Y(_15361_));
 sky130_fd_sc_hd__o21ai_2 _37412_ (.A1(_15222_),
    .A2(_15214_),
    .B1(_15227_),
    .Y(_15362_));
 sky130_fd_sc_hd__nand2_2 _37413_ (.A(_15346_),
    .B(_15350_),
    .Y(_15363_));
 sky130_fd_sc_hd__nor2_2 _37414_ (.A(_15354_),
    .B(_15358_),
    .Y(_15364_));
 sky130_fd_sc_hd__nand2_2 _37415_ (.A(_15363_),
    .B(_15364_),
    .Y(_15365_));
 sky130_fd_sc_hd__nand3_2 _37416_ (.A(_15356_),
    .B(_15350_),
    .C(_15346_),
    .Y(_15366_));
 sky130_fd_sc_hd__nand3_2 _37417_ (.A(_15362_),
    .B(_15365_),
    .C(_15366_),
    .Y(_15367_));
 sky130_fd_sc_hd__o21ai_2 _37418_ (.A1(_14868_),
    .A2(_08604_),
    .B1(_15218_),
    .Y(_15368_));
 sky130_fd_sc_hd__a21oi_2 _37419_ (.A1(_15368_),
    .A2(_15216_),
    .B1(_15217_),
    .Y(_15369_));
 sky130_fd_sc_hd__nand3_2 _37420_ (.A(_09826_),
    .B(_10158_),
    .C(_19573_),
    .Y(_15370_));
 sky130_fd_sc_hd__nor2_2 _37421_ (.A(_09678_),
    .B(_15370_),
    .Y(_15371_));
 sky130_fd_sc_hd__a22o_2 _37422_ (.A1(_09826_),
    .A2(_19577_),
    .B1(_10158_),
    .B2(_19573_),
    .X(_15372_));
 sky130_fd_sc_hd__inv_2 _37423_ (.A(_15372_),
    .Y(_15373_));
 sky130_fd_sc_hd__nor2_2 _37424_ (.A(_08423_),
    .B(_12088_),
    .Y(_15374_));
 sky130_fd_sc_hd__inv_2 _37425_ (.A(_15374_),
    .Y(_15375_));
 sky130_fd_sc_hd__o21ai_2 _37426_ (.A1(_15371_),
    .A2(_15373_),
    .B1(_15375_),
    .Y(_15376_));
 sky130_fd_sc_hd__nand3b_2 _37427_ (.A_N(_15371_),
    .B(_15372_),
    .C(_15374_),
    .Y(_15377_));
 sky130_fd_sc_hd__nand3b_2 _37428_ (.A_N(_15369_),
    .B(_15376_),
    .C(_15377_),
    .Y(_15378_));
 sky130_fd_sc_hd__o21ai_2 _37429_ (.A1(_15371_),
    .A2(_15373_),
    .B1(_15374_),
    .Y(_15379_));
 sky130_fd_sc_hd__nand3b_2 _37430_ (.A_N(_15371_),
    .B(_15375_),
    .C(_15372_),
    .Y(_15380_));
 sky130_fd_sc_hd__nand3_2 _37431_ (.A(_15379_),
    .B(_15380_),
    .C(_15369_),
    .Y(_15381_));
 sky130_fd_sc_hd__o21ai_2 _37432_ (.A1(_15191_),
    .A2(_15193_),
    .B1(_15197_),
    .Y(_15382_));
 sky130_fd_sc_hd__a21oi_2 _37433_ (.A1(_15378_),
    .A2(_15381_),
    .B1(_15382_),
    .Y(_15383_));
 sky130_fd_sc_hd__and3_2 _37434_ (.A(_15378_),
    .B(_15381_),
    .C(_15382_),
    .X(_15384_));
 sky130_fd_sc_hd__nor2_2 _37435_ (.A(_15383_),
    .B(_15384_),
    .Y(_15385_));
 sky130_fd_sc_hd__a21oi_2 _37436_ (.A1(_15361_),
    .A2(_15367_),
    .B1(_15385_),
    .Y(_15386_));
 sky130_fd_sc_hd__nand2_2 _37437_ (.A(_15362_),
    .B(_15365_),
    .Y(_15387_));
 sky130_fd_sc_hd__o211a_2 _37438_ (.A1(_15359_),
    .A2(_15387_),
    .B1(_15361_),
    .C1(_15385_),
    .X(_15388_));
 sky130_fd_sc_hd__a21o_2 _37439_ (.A1(_15200_),
    .A2(_15201_),
    .B1(_15202_),
    .X(_15389_));
 sky130_fd_sc_hd__nand2_2 _37440_ (.A(_15389_),
    .B(_15204_),
    .Y(_15390_));
 sky130_fd_sc_hd__o21a_2 _37441_ (.A1(_15390_),
    .A2(_15230_),
    .B1(_15236_),
    .X(_15391_));
 sky130_fd_sc_hd__o21ai_2 _37442_ (.A1(_15386_),
    .A2(_15388_),
    .B1(_15391_),
    .Y(_15392_));
 sky130_fd_sc_hd__inv_2 _37443_ (.A(_15228_),
    .Y(_15393_));
 sky130_fd_sc_hd__nand2_2 _37444_ (.A(_15223_),
    .B(_15229_),
    .Y(_15394_));
 sky130_fd_sc_hd__o22ai_2 _37445_ (.A1(_15393_),
    .A2(_15394_),
    .B1(_15390_),
    .B2(_15230_),
    .Y(_15395_));
 sky130_fd_sc_hd__o2bb2ai_2 _37446_ (.A1_N(_15367_),
    .A2_N(_15361_),
    .B1(_15383_),
    .B2(_15384_),
    .Y(_15396_));
 sky130_fd_sc_hd__nand3_2 _37447_ (.A(_15361_),
    .B(_15385_),
    .C(_15367_),
    .Y(_15397_));
 sky130_fd_sc_hd__nand3_2 _37448_ (.A(_15395_),
    .B(_15396_),
    .C(_15397_),
    .Y(_15398_));
 sky130_fd_sc_hd__and2_2 _37449_ (.A(_14897_),
    .B(_14894_),
    .X(_15399_));
 sky130_fd_sc_hd__a21oi_2 _37450_ (.A1(_15197_),
    .A2(_15195_),
    .B1(_15199_),
    .Y(_15400_));
 sky130_fd_sc_hd__o21ai_2 _37451_ (.A1(_15399_),
    .A2(_15400_),
    .B1(_15201_),
    .Y(_15401_));
 sky130_fd_sc_hd__and4_2 _37452_ (.A(_10655_),
    .B(_13454_),
    .C(_19565_),
    .D(_08922_),
    .X(_15402_));
 sky130_fd_sc_hd__o22a_2 _37453_ (.A1(_14645_),
    .A2(_08487_),
    .B1(_14097_),
    .B2(_15159_),
    .X(_15403_));
 sky130_fd_sc_hd__nor2_2 _37454_ (.A(_07718_),
    .B(_10523_),
    .Y(_15404_));
 sky130_fd_sc_hd__o21bai_2 _37455_ (.A1(_15402_),
    .A2(_15403_),
    .B1_N(_15404_),
    .Y(_15405_));
 sky130_fd_sc_hd__a22o_2 _37456_ (.A1(_14095_),
    .A2(_09223_),
    .B1(_19341_),
    .B2(_08921_),
    .X(_15406_));
 sky130_fd_sc_hd__nand3b_2 _37457_ (.A_N(_15402_),
    .B(_15406_),
    .C(_15404_),
    .Y(_15407_));
 sky130_fd_sc_hd__a21oi_2 _37458_ (.A1(_15160_),
    .A2(_15162_),
    .B1(_15157_),
    .Y(_15408_));
 sky130_fd_sc_hd__inv_2 _37459_ (.A(_15408_),
    .Y(_15409_));
 sky130_fd_sc_hd__a21oi_2 _37460_ (.A1(_15405_),
    .A2(_15407_),
    .B1(_15409_),
    .Y(_15410_));
 sky130_fd_sc_hd__nand2_2 _37461_ (.A(_15405_),
    .B(_15407_),
    .Y(_15411_));
 sky130_fd_sc_hd__nor2_2 _37462_ (.A(_15408_),
    .B(_15411_),
    .Y(_15412_));
 sky130_fd_sc_hd__nor2_2 _37463_ (.A(_11251_),
    .B(_10533_),
    .Y(_15413_));
 sky130_fd_sc_hd__nand2_2 _37464_ (.A(_09101_),
    .B(_19350_),
    .Y(_15414_));
 sky130_fd_sc_hd__nand2_2 _37465_ (.A(_10050_),
    .B(_19558_),
    .Y(_15415_));
 sky130_fd_sc_hd__a22o_2 _37466_ (.A1(_07481_),
    .A2(_09736_),
    .B1(_08809_),
    .B2(_19553_),
    .X(_15416_));
 sky130_fd_sc_hd__o21ai_2 _37467_ (.A1(_15414_),
    .A2(_15415_),
    .B1(_15416_),
    .Y(_15417_));
 sky130_fd_sc_hd__xor2_2 _37468_ (.A(_15413_),
    .B(_15417_),
    .X(_15418_));
 sky130_fd_sc_hd__inv_2 _37469_ (.A(_15418_),
    .Y(_15419_));
 sky130_fd_sc_hd__o21ai_2 _37470_ (.A1(_15410_),
    .A2(_15412_),
    .B1(_15419_),
    .Y(_15420_));
 sky130_fd_sc_hd__nand2_2 _37471_ (.A(_15411_),
    .B(_15408_),
    .Y(_15421_));
 sky130_fd_sc_hd__nand3_2 _37472_ (.A(_15409_),
    .B(_15405_),
    .C(_15407_),
    .Y(_15422_));
 sky130_fd_sc_hd__nand3_2 _37473_ (.A(_15421_),
    .B(_15418_),
    .C(_15422_),
    .Y(_15423_));
 sky130_fd_sc_hd__nand3b_2 _37474_ (.A_N(_15401_),
    .B(_15420_),
    .C(_15423_),
    .Y(_15424_));
 sky130_fd_sc_hd__o21ai_2 _37475_ (.A1(_15410_),
    .A2(_15412_),
    .B1(_15418_),
    .Y(_15425_));
 sky130_fd_sc_hd__nand3_2 _37476_ (.A(_15419_),
    .B(_15421_),
    .C(_15422_),
    .Y(_15426_));
 sky130_fd_sc_hd__nand3_2 _37477_ (.A(_15425_),
    .B(_15401_),
    .C(_15426_),
    .Y(_15427_));
 sky130_fd_sc_hd__inv_2 _37478_ (.A(_15166_),
    .Y(_15428_));
 sky130_fd_sc_hd__and3_2 _37479_ (.A(_15168_),
    .B(_15175_),
    .C(_15172_),
    .X(_15429_));
 sky130_fd_sc_hd__nor2_2 _37480_ (.A(_15428_),
    .B(_15429_),
    .Y(_15430_));
 sky130_fd_sc_hd__a21oi_2 _37481_ (.A1(_15424_),
    .A2(_15427_),
    .B1(_15430_),
    .Y(_15431_));
 sky130_fd_sc_hd__and3_2 _37482_ (.A(_15424_),
    .B(_15427_),
    .C(_15430_),
    .X(_15432_));
 sky130_fd_sc_hd__nor2_2 _37483_ (.A(_15431_),
    .B(_15432_),
    .Y(_15433_));
 sky130_fd_sc_hd__a21o_2 _37484_ (.A1(_15392_),
    .A2(_15398_),
    .B1(_15433_),
    .X(_15434_));
 sky130_fd_sc_hd__a21o_2 _37485_ (.A1(_15184_),
    .A2(_15188_),
    .B1(_15186_),
    .X(_15435_));
 sky130_fd_sc_hd__o21ai_2 _37486_ (.A1(_15435_),
    .A2(_15240_),
    .B1(_15247_),
    .Y(_15436_));
 sky130_fd_sc_hd__nand3_2 _37487_ (.A(_15433_),
    .B(_15392_),
    .C(_15398_),
    .Y(_15437_));
 sky130_fd_sc_hd__nand3_2 _37488_ (.A(_15434_),
    .B(_15436_),
    .C(_15437_),
    .Y(_15438_));
 sky130_fd_sc_hd__o21a_2 _37489_ (.A1(_15186_),
    .A2(_15189_),
    .B1(_15247_),
    .X(_15439_));
 sky130_fd_sc_hd__o2bb2ai_2 _37490_ (.A1_N(_15424_),
    .A2_N(_15427_),
    .B1(_15428_),
    .B2(_15429_),
    .Y(_15440_));
 sky130_fd_sc_hd__nand3_2 _37491_ (.A(_15424_),
    .B(_15427_),
    .C(_15430_),
    .Y(_15441_));
 sky130_fd_sc_hd__a22oi_2 _37492_ (.A1(_15440_),
    .A2(_15441_),
    .B1(_15392_),
    .B2(_15398_),
    .Y(_15442_));
 sky130_fd_sc_hd__nand2_2 _37493_ (.A(_15440_),
    .B(_15441_),
    .Y(_15443_));
 sky130_fd_sc_hd__a21oi_2 _37494_ (.A1(_15396_),
    .A2(_15397_),
    .B1(_15395_),
    .Y(_15444_));
 sky130_fd_sc_hd__nor3b_2 _37495_ (.A(_15443_),
    .B(_15444_),
    .C_N(_15398_),
    .Y(_15445_));
 sky130_fd_sc_hd__o22ai_2 _37496_ (.A1(_15240_),
    .A2(_15439_),
    .B1(_15442_),
    .B2(_15445_),
    .Y(_15446_));
 sky130_fd_sc_hd__nand2_2 _37497_ (.A(_19355_),
    .B(_19545_),
    .Y(_15447_));
 sky130_fd_sc_hd__nand2_2 _37498_ (.A(_19358_),
    .B(_19541_),
    .Y(_15448_));
 sky130_fd_sc_hd__nor2_2 _37499_ (.A(_15447_),
    .B(_15448_),
    .Y(_15449_));
 sky130_fd_sc_hd__and2_2 _37500_ (.A(_15447_),
    .B(_15448_),
    .X(_15450_));
 sky130_fd_sc_hd__nand2_2 _37501_ (.A(_14153_),
    .B(_09386_),
    .Y(_15451_));
 sky130_fd_sc_hd__o21ai_2 _37502_ (.A1(_15449_),
    .A2(_15450_),
    .B1(_15451_),
    .Y(_15452_));
 sky130_fd_sc_hd__or2_2 _37503_ (.A(_15447_),
    .B(_15448_),
    .X(_15453_));
 sky130_fd_sc_hd__inv_2 _37504_ (.A(_15451_),
    .Y(_15454_));
 sky130_fd_sc_hd__nand2_2 _37505_ (.A(_15447_),
    .B(_15448_),
    .Y(_15455_));
 sky130_fd_sc_hd__nand3_2 _37506_ (.A(_15453_),
    .B(_15454_),
    .C(_15455_),
    .Y(_15456_));
 sky130_fd_sc_hd__a21o_2 _37507_ (.A1(_15171_),
    .A2(_15174_),
    .B1(_15169_),
    .X(_15457_));
 sky130_fd_sc_hd__a21o_2 _37508_ (.A1(_15452_),
    .A2(_15456_),
    .B1(_15457_),
    .X(_15458_));
 sky130_fd_sc_hd__nand3_2 _37509_ (.A(_15457_),
    .B(_15452_),
    .C(_15456_),
    .Y(_15459_));
 sky130_fd_sc_hd__nand2_2 _37510_ (.A(_15119_),
    .B(_15115_),
    .Y(_15460_));
 sky130_fd_sc_hd__a21oi_2 _37511_ (.A1(_15458_),
    .A2(_15459_),
    .B1(_15460_),
    .Y(_15461_));
 sky130_fd_sc_hd__and3_2 _37512_ (.A(_15458_),
    .B(_15459_),
    .C(_15460_),
    .X(_15462_));
 sky130_fd_sc_hd__inv_2 _37513_ (.A(_15123_),
    .Y(_15463_));
 sky130_fd_sc_hd__a21oi_2 _37514_ (.A1(_15117_),
    .A2(_15119_),
    .B1(_15120_),
    .Y(_15464_));
 sky130_fd_sc_hd__o21ai_2 _37515_ (.A1(_15463_),
    .A2(_15464_),
    .B1(_15122_),
    .Y(_15465_));
 sky130_fd_sc_hd__o21bai_2 _37516_ (.A1(_15461_),
    .A2(_15462_),
    .B1_N(_15465_),
    .Y(_15466_));
 sky130_fd_sc_hd__a21o_2 _37517_ (.A1(_15458_),
    .A2(_15459_),
    .B1(_15460_),
    .X(_15467_));
 sky130_fd_sc_hd__nand3_2 _37518_ (.A(_15458_),
    .B(_15459_),
    .C(_15460_),
    .Y(_15468_));
 sky130_fd_sc_hd__nand3_2 _37519_ (.A(_15467_),
    .B(_15465_),
    .C(_15468_),
    .Y(_15469_));
 sky130_fd_sc_hd__and2_2 _37520_ (.A(_15130_),
    .B(_06628_),
    .X(_15470_));
 sky130_fd_sc_hd__a21oi_2 _37521_ (.A1(_14712_),
    .A2(_15129_),
    .B1(_15470_),
    .Y(_15471_));
 sky130_fd_sc_hd__nor2_2 _37522_ (.A(_15471_),
    .B(_14429_),
    .Y(_15472_));
 sky130_fd_sc_hd__and2b_2 _37523_ (.A_N(_14759_),
    .B(_15471_),
    .X(_15473_));
 sky130_fd_sc_hd__nor2_2 _37524_ (.A(_15472_),
    .B(_15473_),
    .Y(_15474_));
 sky130_fd_sc_hd__buf_1 _37525_ (.A(_15474_),
    .X(_15475_));
 sky130_fd_sc_hd__buf_1 _37526_ (.A(_15475_),
    .X(_15476_));
 sky130_fd_sc_hd__a21oi_2 _37527_ (.A1(_15466_),
    .A2(_15469_),
    .B1(_15476_),
    .Y(_15477_));
 sky130_fd_sc_hd__buf_1 _37528_ (.A(_15474_),
    .X(_15478_));
 sky130_fd_sc_hd__and3_2 _37529_ (.A(_15466_),
    .B(_15469_),
    .C(_15478_),
    .X(_15479_));
 sky130_fd_sc_hd__a21oi_2 _37530_ (.A1(_15181_),
    .A2(_15183_),
    .B1(_15182_),
    .Y(_15480_));
 sky130_fd_sc_hd__o21ai_2 _37531_ (.A1(_15185_),
    .A2(_15480_),
    .B1(_15184_),
    .Y(_15481_));
 sky130_fd_sc_hd__inv_2 _37532_ (.A(_15481_),
    .Y(_15482_));
 sky130_fd_sc_hd__o21ai_2 _37533_ (.A1(_15477_),
    .A2(_15479_),
    .B1(_15482_),
    .Y(_15483_));
 sky130_fd_sc_hd__a21o_2 _37534_ (.A1(_15466_),
    .A2(_15469_),
    .B1(_15475_),
    .X(_15484_));
 sky130_fd_sc_hd__nand3_2 _37535_ (.A(_15466_),
    .B(_15469_),
    .C(_15475_),
    .Y(_15485_));
 sky130_fd_sc_hd__nand3_2 _37536_ (.A(_15484_),
    .B(_15485_),
    .C(_15481_),
    .Y(_15486_));
 sky130_fd_sc_hd__o21ai_2 _37537_ (.A1(_15127_),
    .A2(_15140_),
    .B1(_15142_),
    .Y(_15487_));
 sky130_fd_sc_hd__a21oi_2 _37538_ (.A1(_15483_),
    .A2(_15486_),
    .B1(_15487_),
    .Y(_15488_));
 sky130_fd_sc_hd__and3_2 _37539_ (.A(_15483_),
    .B(_15486_),
    .C(_15487_),
    .X(_15489_));
 sky130_fd_sc_hd__o2bb2ai_2 _37540_ (.A1_N(_15438_),
    .A2_N(_15446_),
    .B1(_15488_),
    .B2(_15489_),
    .Y(_15490_));
 sky130_fd_sc_hd__nand2_2 _37541_ (.A(_15484_),
    .B(_15485_),
    .Y(_15491_));
 sky130_fd_sc_hd__a21boi_2 _37542_ (.A1(_15491_),
    .A2(_15482_),
    .B1_N(_15487_),
    .Y(_15492_));
 sky130_fd_sc_hd__a21oi_2 _37543_ (.A1(_15486_),
    .A2(_15492_),
    .B1(_15488_),
    .Y(_15493_));
 sky130_fd_sc_hd__nand3_2 _37544_ (.A(_15493_),
    .B(_15446_),
    .C(_15438_),
    .Y(_15494_));
 sky130_fd_sc_hd__nand2_2 _37545_ (.A(_15244_),
    .B(_15251_),
    .Y(_15495_));
 sky130_fd_sc_hd__o22ai_2 _37546_ (.A1(_15258_),
    .A2(_15495_),
    .B1(_15257_),
    .B2(_15252_),
    .Y(_15496_));
 sky130_fd_sc_hd__a21oi_2 _37547_ (.A1(_15490_),
    .A2(_15494_),
    .B1(_15496_),
    .Y(_15497_));
 sky130_fd_sc_hd__a21oi_2 _37548_ (.A1(_15434_),
    .A2(_15437_),
    .B1(_15436_),
    .Y(_15498_));
 sky130_fd_sc_hd__nand2_2 _37549_ (.A(_15493_),
    .B(_15438_),
    .Y(_15499_));
 sky130_fd_sc_hd__o211a_2 _37550_ (.A1(_15498_),
    .A2(_15499_),
    .B1(_15490_),
    .C1(_15496_),
    .X(_15500_));
 sky130_fd_sc_hd__nand2_2 _37551_ (.A(_15145_),
    .B(_15147_),
    .Y(_15501_));
 sky130_fd_sc_hd__nand2_2 _37552_ (.A(_14764_),
    .B(_13965_),
    .Y(_15502_));
 sky130_fd_sc_hd__nand2_2 _37553_ (.A(_14763_),
    .B(_14765_),
    .Y(_15503_));
 sky130_fd_sc_hd__nand2_2 _37554_ (.A(_15502_),
    .B(_15503_),
    .Y(_15504_));
 sky130_fd_sc_hd__a211o_2 _37555_ (.A1(_15136_),
    .A2(_14430_),
    .B1(_15470_),
    .C1(_15504_),
    .X(_15505_));
 sky130_fd_sc_hd__o21ai_2 _37556_ (.A1(_15470_),
    .A2(_15135_),
    .B1(_15504_),
    .Y(_15506_));
 sky130_fd_sc_hd__and3_2 _37557_ (.A(_15505_),
    .B(_15274_),
    .C(_15506_),
    .X(_15507_));
 sky130_fd_sc_hd__nand2_2 _37558_ (.A(_15507_),
    .B(_15281_),
    .Y(_15508_));
 sky130_fd_sc_hd__a22o_2 _37559_ (.A1(_15505_),
    .A2(_15506_),
    .B1(_15281_),
    .B2(_15274_),
    .X(_15509_));
 sky130_fd_sc_hd__nand3_2 _37560_ (.A(_15508_),
    .B(_14482_),
    .C(_15509_),
    .Y(_15510_));
 sky130_fd_sc_hd__a21o_2 _37561_ (.A1(_15508_),
    .A2(_15509_),
    .B1(_14482_),
    .X(_15511_));
 sky130_fd_sc_hd__o2111ai_2 _37562_ (.A1(_15111_),
    .A2(_15501_),
    .B1(_15510_),
    .C1(_15153_),
    .D1(_15511_),
    .Y(_15512_));
 sky130_fd_sc_hd__nand2_2 _37563_ (.A(_15511_),
    .B(_15510_),
    .Y(_15513_));
 sky130_fd_sc_hd__nand2_2 _37564_ (.A(_15153_),
    .B(_15148_),
    .Y(_15514_));
 sky130_fd_sc_hd__nand2_2 _37565_ (.A(_15279_),
    .B(_14794_),
    .Y(_15515_));
 sky130_fd_sc_hd__and2_2 _37566_ (.A(_15515_),
    .B(_15282_),
    .X(_15516_));
 sky130_fd_sc_hd__a21oi_2 _37567_ (.A1(_15513_),
    .A2(_15514_),
    .B1(_15516_),
    .Y(_15517_));
 sky130_fd_sc_hd__nand2_2 _37568_ (.A(_15513_),
    .B(_15514_),
    .Y(_15518_));
 sky130_fd_sc_hd__a21boi_2 _37569_ (.A1(_15518_),
    .A2(_15512_),
    .B1_N(_15516_),
    .Y(_15519_));
 sky130_fd_sc_hd__a21oi_2 _37570_ (.A1(_15512_),
    .A2(_15517_),
    .B1(_15519_),
    .Y(_15520_));
 sky130_fd_sc_hd__o21ai_2 _37571_ (.A1(_15497_),
    .A2(_15500_),
    .B1(_15520_),
    .Y(_15521_));
 sky130_fd_sc_hd__a21boi_2 _37572_ (.A1(_15268_),
    .A2(_15297_),
    .B1_N(_15264_),
    .Y(_15522_));
 sky130_fd_sc_hd__nand2_2 _37573_ (.A(_15518_),
    .B(_15512_),
    .Y(_15523_));
 sky130_fd_sc_hd__nor2_2 _37574_ (.A(_15516_),
    .B(_15523_),
    .Y(_15524_));
 sky130_fd_sc_hd__nand3_2 _37575_ (.A(_15496_),
    .B(_15490_),
    .C(_15494_),
    .Y(_15525_));
 sky130_fd_sc_hd__a21o_2 _37576_ (.A1(_15490_),
    .A2(_15494_),
    .B1(_15496_),
    .X(_15526_));
 sky130_fd_sc_hd__o211ai_2 _37577_ (.A1(_15519_),
    .A2(_15524_),
    .B1(_15525_),
    .C1(_15526_),
    .Y(_15527_));
 sky130_fd_sc_hd__nand3_2 _37578_ (.A(_15521_),
    .B(_15522_),
    .C(_15527_),
    .Y(_15528_));
 sky130_fd_sc_hd__o22ai_2 _37579_ (.A1(_15524_),
    .A2(_15519_),
    .B1(_15497_),
    .B2(_15500_),
    .Y(_15529_));
 sky130_fd_sc_hd__inv_2 _37580_ (.A(_15262_),
    .Y(_15530_));
 sky130_fd_sc_hd__nand2_2 _37581_ (.A(_15255_),
    .B(_15263_),
    .Y(_15531_));
 sky130_fd_sc_hd__o2bb2ai_2 _37582_ (.A1_N(_15297_),
    .A2_N(_15268_),
    .B1(_15530_),
    .B2(_15531_),
    .Y(_15532_));
 sky130_fd_sc_hd__nand3_2 _37583_ (.A(_15526_),
    .B(_15520_),
    .C(_15525_),
    .Y(_15533_));
 sky130_fd_sc_hd__nand3_2 _37584_ (.A(_15529_),
    .B(_15532_),
    .C(_15533_),
    .Y(_15534_));
 sky130_fd_sc_hd__nor2b_2 _37585_ (.A(_15296_),
    .B_N(_15290_),
    .Y(_15535_));
 sky130_fd_sc_hd__nor2_2 _37586_ (.A(_15081_),
    .B(_15535_),
    .Y(_15536_));
 sky130_fd_sc_hd__and2_2 _37587_ (.A(_15535_),
    .B(_13736_),
    .X(_15537_));
 sky130_fd_sc_hd__nor2_2 _37588_ (.A(_15536_),
    .B(_15537_),
    .Y(_15538_));
 sky130_fd_sc_hd__nand3_2 _37589_ (.A(_15528_),
    .B(_15534_),
    .C(_15538_),
    .Y(_15539_));
 sky130_fd_sc_hd__o2bb2ai_2 _37590_ (.A1_N(_15534_),
    .A2_N(_15528_),
    .B1(_15536_),
    .B2(_15537_),
    .Y(_15540_));
 sky130_fd_sc_hd__o2111ai_2 _37591_ (.A1(_15302_),
    .A2(_15310_),
    .B1(_15312_),
    .C1(_15539_),
    .D1(_15540_),
    .Y(_15541_));
 sky130_fd_sc_hd__o21ai_2 _37592_ (.A1(_15310_),
    .A2(_15302_),
    .B1(_15312_),
    .Y(_15542_));
 sky130_fd_sc_hd__nor2_2 _37593_ (.A(_14018_),
    .B(_15535_),
    .Y(_15543_));
 sky130_fd_sc_hd__and2_2 _37594_ (.A(_15535_),
    .B(_14823_),
    .X(_15544_));
 sky130_fd_sc_hd__o2bb2ai_2 _37595_ (.A1_N(_15534_),
    .A2_N(_15528_),
    .B1(_15543_),
    .B2(_15544_),
    .Y(_15545_));
 sky130_fd_sc_hd__nand3b_2 _37596_ (.A_N(_15538_),
    .B(_15528_),
    .C(_15534_),
    .Y(_15546_));
 sky130_fd_sc_hd__nand3_2 _37597_ (.A(_15542_),
    .B(_15545_),
    .C(_15546_),
    .Y(_15547_));
 sky130_fd_sc_hd__a21oi_2 _37598_ (.A1(_15541_),
    .A2(_15547_),
    .B1(_15108_),
    .Y(_15548_));
 sky130_fd_sc_hd__and3_2 _37599_ (.A(_15541_),
    .B(_15547_),
    .C(_15108_),
    .X(_15549_));
 sky130_fd_sc_hd__inv_2 _37600_ (.A(_15313_),
    .Y(_15550_));
 sky130_fd_sc_hd__nand2_2 _37601_ (.A(_15306_),
    .B(_15314_),
    .Y(_15551_));
 sky130_fd_sc_hd__o2bb2ai_2 _37602_ (.A1_N(_15083_),
    .A2_N(_15319_),
    .B1(_15550_),
    .B2(_15551_),
    .Y(_15552_));
 sky130_fd_sc_hd__o21bai_2 _37603_ (.A1(_15548_),
    .A2(_15549_),
    .B1_N(_15552_),
    .Y(_15553_));
 sky130_fd_sc_hd__a21o_2 _37604_ (.A1(_15541_),
    .A2(_15547_),
    .B1(_15108_),
    .X(_15554_));
 sky130_fd_sc_hd__nand3_2 _37605_ (.A(_15541_),
    .B(_15547_),
    .C(_15108_),
    .Y(_15555_));
 sky130_fd_sc_hd__nand3_2 _37606_ (.A(_15554_),
    .B(_15552_),
    .C(_15555_),
    .Y(_15556_));
 sky130_fd_sc_hd__and2_2 _37607_ (.A(_15553_),
    .B(_15556_),
    .X(_15557_));
 sky130_fd_sc_hd__o21ai_2 _37608_ (.A1(_15329_),
    .A2(_15336_),
    .B1(_15327_),
    .Y(_15558_));
 sky130_fd_sc_hd__xor2_2 _37609_ (.A(_15557_),
    .B(_15558_),
    .X(_02666_));
 sky130_fd_sc_hd__inv_2 _37610_ (.A(_15534_),
    .Y(_15559_));
 sky130_fd_sc_hd__o21a_2 _37611_ (.A1(_15536_),
    .A2(_15537_),
    .B1(_15528_),
    .X(_15560_));
 sky130_fd_sc_hd__o31a_2 _37612_ (.A1(_15488_),
    .A2(_15489_),
    .A3(_15498_),
    .B1(_15438_),
    .X(_15561_));
 sky130_fd_sc_hd__nand2_2 _37613_ (.A(_15441_),
    .B(_15427_),
    .Y(_15562_));
 sky130_fd_sc_hd__nand2_2 _37614_ (.A(_06822_),
    .B(_19540_),
    .Y(_15563_));
 sky130_fd_sc_hd__nand2_2 _37615_ (.A(_11023_),
    .B(_07652_),
    .Y(_15564_));
 sky130_fd_sc_hd__nor2_2 _37616_ (.A(_15563_),
    .B(_15564_),
    .Y(_15565_));
 sky130_fd_sc_hd__nand2_2 _37617_ (.A(_15563_),
    .B(_15564_),
    .Y(_15566_));
 sky130_fd_sc_hd__and2b_2 _37618_ (.A_N(_15565_),
    .B(_15566_),
    .X(_15567_));
 sky130_fd_sc_hd__nand2_2 _37619_ (.A(_15567_),
    .B(_15454_),
    .Y(_15568_));
 sky130_fd_sc_hd__or2_2 _37620_ (.A(_15563_),
    .B(_15564_),
    .X(_15569_));
 sky130_fd_sc_hd__a21o_2 _37621_ (.A1(_15569_),
    .A2(_15566_),
    .B1(_15454_),
    .X(_15570_));
 sky130_fd_sc_hd__nand2_2 _37622_ (.A(_15568_),
    .B(_15570_),
    .Y(_15571_));
 sky130_fd_sc_hd__o2bb2a_2 _37623_ (.A1_N(_15416_),
    .A2_N(_15413_),
    .B1(_15414_),
    .B2(_15415_),
    .X(_15572_));
 sky130_fd_sc_hd__nand2_2 _37624_ (.A(_15571_),
    .B(_15572_),
    .Y(_15573_));
 sky130_fd_sc_hd__nand3b_2 _37625_ (.A_N(_15572_),
    .B(_15568_),
    .C(_15570_),
    .Y(_15574_));
 sky130_fd_sc_hd__nand2_2 _37626_ (.A(_15456_),
    .B(_15453_),
    .Y(_15575_));
 sky130_fd_sc_hd__nand3_2 _37627_ (.A(_15573_),
    .B(_15574_),
    .C(_15575_),
    .Y(_15576_));
 sky130_fd_sc_hd__a21o_2 _37628_ (.A1(_15573_),
    .A2(_15574_),
    .B1(_15575_),
    .X(_15577_));
 sky130_fd_sc_hd__and2_2 _37629_ (.A(_15468_),
    .B(_15459_),
    .X(_15578_));
 sky130_fd_sc_hd__a21boi_2 _37630_ (.A1(_15576_),
    .A2(_15577_),
    .B1_N(_15578_),
    .Y(_15579_));
 sky130_fd_sc_hd__nand2_2 _37631_ (.A(_15577_),
    .B(_15576_),
    .Y(_15580_));
 sky130_fd_sc_hd__nor2_2 _37632_ (.A(_15578_),
    .B(_15580_),
    .Y(_15581_));
 sky130_fd_sc_hd__o21ai_2 _37633_ (.A1(_15579_),
    .A2(_15581_),
    .B1(_15476_),
    .Y(_15582_));
 sky130_fd_sc_hd__a21o_2 _37634_ (.A1(_15459_),
    .A2(_15468_),
    .B1(_15580_),
    .X(_15583_));
 sky130_fd_sc_hd__or2_2 _37635_ (.A(_15472_),
    .B(_15473_),
    .X(_15584_));
 sky130_fd_sc_hd__buf_1 _37636_ (.A(_15584_),
    .X(_15585_));
 sky130_fd_sc_hd__buf_1 _37637_ (.A(_15585_),
    .X(_15586_));
 sky130_fd_sc_hd__nand2_2 _37638_ (.A(_15580_),
    .B(_15578_),
    .Y(_15587_));
 sky130_fd_sc_hd__nand3_2 _37639_ (.A(_15583_),
    .B(_15586_),
    .C(_15587_),
    .Y(_15588_));
 sky130_fd_sc_hd__nand3b_2 _37640_ (.A_N(_15562_),
    .B(_15582_),
    .C(_15588_),
    .Y(_15589_));
 sky130_fd_sc_hd__nand2_2 _37641_ (.A(_15587_),
    .B(_15478_),
    .Y(_15590_));
 sky130_fd_sc_hd__o21ai_2 _37642_ (.A1(_15579_),
    .A2(_15581_),
    .B1(_15586_),
    .Y(_15591_));
 sky130_fd_sc_hd__o211ai_2 _37643_ (.A1(_15581_),
    .A2(_15590_),
    .B1(_15562_),
    .C1(_15591_),
    .Y(_15592_));
 sky130_fd_sc_hd__nand2_2 _37644_ (.A(_15589_),
    .B(_15592_),
    .Y(_15593_));
 sky130_fd_sc_hd__inv_2 _37645_ (.A(_15466_),
    .Y(_15594_));
 sky130_fd_sc_hd__and2_2 _37646_ (.A(_15469_),
    .B(_15585_),
    .X(_15595_));
 sky130_fd_sc_hd__nor2_2 _37647_ (.A(_15594_),
    .B(_15595_),
    .Y(_15596_));
 sky130_fd_sc_hd__inv_2 _37648_ (.A(_15596_),
    .Y(_15597_));
 sky130_fd_sc_hd__nand2_2 _37649_ (.A(_15593_),
    .B(_15597_),
    .Y(_15598_));
 sky130_fd_sc_hd__inv_2 _37650_ (.A(_15598_),
    .Y(_15599_));
 sky130_fd_sc_hd__nand3_2 _37651_ (.A(_15589_),
    .B(_15592_),
    .C(_15596_),
    .Y(_15600_));
 sky130_fd_sc_hd__inv_2 _37652_ (.A(_15600_),
    .Y(_15601_));
 sky130_fd_sc_hd__and4_2 _37653_ (.A(_08045_),
    .B(_11514_),
    .C(_19307_),
    .D(_06944_),
    .X(_15602_));
 sky130_fd_sc_hd__o22a_2 _37654_ (.A1(_06750_),
    .A2(_10830_),
    .B1(_10832_),
    .B2(_07833_),
    .X(_15603_));
 sky130_fd_sc_hd__nor2_2 _37655_ (.A(_15602_),
    .B(_15603_),
    .Y(_15604_));
 sky130_fd_sc_hd__nand3_2 _37656_ (.A(_15604_),
    .B(_19314_),
    .C(_19586_),
    .Y(_15605_));
 sky130_fd_sc_hd__nand2_2 _37657_ (.A(_10827_),
    .B(_19586_),
    .Y(_15606_));
 sky130_fd_sc_hd__o21ai_2 _37658_ (.A1(_15602_),
    .A2(_15603_),
    .B1(_15606_),
    .Y(_15607_));
 sky130_fd_sc_hd__a21o_2 _37659_ (.A1(_15343_),
    .A2(_15344_),
    .B1(_15338_),
    .X(_15608_));
 sky130_fd_sc_hd__a21o_2 _37660_ (.A1(_15605_),
    .A2(_15607_),
    .B1(_15608_),
    .X(_15609_));
 sky130_fd_sc_hd__nand3_2 _37661_ (.A(_15605_),
    .B(_15607_),
    .C(_15608_),
    .Y(_15610_));
 sky130_fd_sc_hd__nor2_2 _37662_ (.A(_09357_),
    .B(_11660_),
    .Y(_15611_));
 sky130_fd_sc_hd__a22o_2 _37663_ (.A1(_10146_),
    .A2(_08490_),
    .B1(_19320_),
    .B2(_07848_),
    .X(_15612_));
 sky130_fd_sc_hd__o311a_2 _37664_ (.A1(_11178_),
    .A2(_09246_),
    .A3(_08947_),
    .B1(_15611_),
    .C1(_15612_),
    .X(_15613_));
 sky130_fd_sc_hd__or3_2 _37665_ (.A(_10705_),
    .B(_09246_),
    .C(_08957_),
    .X(_15614_));
 sky130_fd_sc_hd__a21oi_2 _37666_ (.A1(_15614_),
    .A2(_15612_),
    .B1(_15611_),
    .Y(_15615_));
 sky130_fd_sc_hd__nor2_2 _37667_ (.A(_15613_),
    .B(_15615_),
    .Y(_15616_));
 sky130_fd_sc_hd__a21oi_2 _37668_ (.A1(_15609_),
    .A2(_15610_),
    .B1(_15616_),
    .Y(_15617_));
 sky130_fd_sc_hd__and3_2 _37669_ (.A(_15609_),
    .B(_15616_),
    .C(_15610_),
    .X(_15618_));
 sky130_fd_sc_hd__nand2_2 _37670_ (.A(_15366_),
    .B(_15346_),
    .Y(_15619_));
 sky130_fd_sc_hd__o21bai_2 _37671_ (.A1(_15617_),
    .A2(_15618_),
    .B1_N(_15619_),
    .Y(_15620_));
 sky130_fd_sc_hd__a21o_2 _37672_ (.A1(_15609_),
    .A2(_15610_),
    .B1(_15616_),
    .X(_15621_));
 sky130_fd_sc_hd__nand3_2 _37673_ (.A(_15609_),
    .B(_15616_),
    .C(_15610_),
    .Y(_15622_));
 sky130_fd_sc_hd__nand3_2 _37674_ (.A(_15621_),
    .B(_15619_),
    .C(_15622_),
    .Y(_15623_));
 sky130_fd_sc_hd__nand2_2 _37675_ (.A(_11205_),
    .B(_12349_),
    .Y(_15624_));
 sky130_fd_sc_hd__nand2_2 _37676_ (.A(_10867_),
    .B(_14112_),
    .Y(_15625_));
 sky130_fd_sc_hd__nand2_2 _37677_ (.A(_15624_),
    .B(_15625_),
    .Y(_15626_));
 sky130_fd_sc_hd__o21ai_2 _37678_ (.A1(_12090_),
    .A2(_15370_),
    .B1(_15626_),
    .Y(_15627_));
 sky130_fd_sc_hd__or3_2 _37679_ (.A(_08424_),
    .B(_09226_),
    .C(_15627_),
    .X(_15628_));
 sky130_fd_sc_hd__o21ai_2 _37680_ (.A1(_08424_),
    .A2(_09226_),
    .B1(_15627_),
    .Y(_15629_));
 sky130_fd_sc_hd__nor2_2 _37681_ (.A(_15352_),
    .B(_15353_),
    .Y(_15630_));
 sky130_fd_sc_hd__nor2_2 _37682_ (.A(_15351_),
    .B(_15630_),
    .Y(_15631_));
 sky130_fd_sc_hd__a21o_2 _37683_ (.A1(_15628_),
    .A2(_15629_),
    .B1(_15631_),
    .X(_15632_));
 sky130_fd_sc_hd__nand3_2 _37684_ (.A(_15628_),
    .B(_15629_),
    .C(_15631_),
    .Y(_15633_));
 sky130_fd_sc_hd__a21o_2 _37685_ (.A1(_15374_),
    .A2(_15372_),
    .B1(_15371_),
    .X(_15634_));
 sky130_fd_sc_hd__a21o_2 _37686_ (.A1(_15632_),
    .A2(_15633_),
    .B1(_15634_),
    .X(_15635_));
 sky130_fd_sc_hd__nand3_2 _37687_ (.A(_15632_),
    .B(_15633_),
    .C(_15634_),
    .Y(_15636_));
 sky130_fd_sc_hd__nand2_2 _37688_ (.A(_15635_),
    .B(_15636_),
    .Y(_15637_));
 sky130_fd_sc_hd__a21o_2 _37689_ (.A1(_15620_),
    .A2(_15623_),
    .B1(_15637_),
    .X(_15638_));
 sky130_fd_sc_hd__and2_2 _37690_ (.A(_15397_),
    .B(_15367_),
    .X(_15639_));
 sky130_fd_sc_hd__nand3_2 _37691_ (.A(_15620_),
    .B(_15623_),
    .C(_15637_),
    .Y(_15640_));
 sky130_fd_sc_hd__nand3_2 _37692_ (.A(_15638_),
    .B(_15639_),
    .C(_15640_),
    .Y(_15641_));
 sky130_fd_sc_hd__nand2_2 _37693_ (.A(_15620_),
    .B(_15623_),
    .Y(_15642_));
 sky130_fd_sc_hd__nand2_2 _37694_ (.A(_15642_),
    .B(_15637_),
    .Y(_15643_));
 sky130_fd_sc_hd__nand3b_2 _37695_ (.A_N(_15637_),
    .B(_15620_),
    .C(_15623_),
    .Y(_15644_));
 sky130_fd_sc_hd__nand3b_2 _37696_ (.A_N(_15639_),
    .B(_15643_),
    .C(_15644_),
    .Y(_15645_));
 sky130_fd_sc_hd__nand2_2 _37697_ (.A(_10655_),
    .B(_19565_),
    .Y(_15646_));
 sky130_fd_sc_hd__a21o_2 _37698_ (.A1(_10656_),
    .A2(_10055_),
    .B1(_15646_),
    .X(_15647_));
 sky130_fd_sc_hd__nand2_2 _37699_ (.A(_13454_),
    .B(_19562_),
    .Y(_15648_));
 sky130_fd_sc_hd__a21o_2 _37700_ (.A1(_14095_),
    .A2(_08921_),
    .B1(_15648_),
    .X(_15649_));
 sky130_fd_sc_hd__a211o_2 _37701_ (.A1(_15647_),
    .A2(_15649_),
    .B1(_12602_),
    .C1(_14939_),
    .X(_15650_));
 sky130_fd_sc_hd__o211ai_2 _37702_ (.A1(_12602_),
    .A2(_14939_),
    .B1(_15649_),
    .C1(_15647_),
    .Y(_15651_));
 sky130_fd_sc_hd__a21o_2 _37703_ (.A1(_15404_),
    .A2(_15406_),
    .B1(_15402_),
    .X(_15652_));
 sky130_fd_sc_hd__a21o_2 _37704_ (.A1(_15650_),
    .A2(_15651_),
    .B1(_15652_),
    .X(_15653_));
 sky130_fd_sc_hd__nand3_2 _37705_ (.A(_15650_),
    .B(_15652_),
    .C(_15651_),
    .Y(_15654_));
 sky130_fd_sc_hd__nand2_2 _37706_ (.A(_12069_),
    .B(_19546_),
    .Y(_15655_));
 sky130_fd_sc_hd__nand2_2 _37707_ (.A(_19549_),
    .B(_19553_),
    .Y(_15656_));
 sky130_fd_sc_hd__a22o_2 _37708_ (.A1(_09101_),
    .A2(_09722_),
    .B1(_08185_),
    .B2(_11765_),
    .X(_15657_));
 sky130_fd_sc_hd__o21ai_2 _37709_ (.A1(_15414_),
    .A2(_15656_),
    .B1(_15657_),
    .Y(_15658_));
 sky130_fd_sc_hd__or2_2 _37710_ (.A(_15655_),
    .B(_15658_),
    .X(_15659_));
 sky130_fd_sc_hd__nand2_2 _37711_ (.A(_15658_),
    .B(_15655_),
    .Y(_15660_));
 sky130_fd_sc_hd__and2_2 _37712_ (.A(_15659_),
    .B(_15660_),
    .X(_15661_));
 sky130_fd_sc_hd__a21o_2 _37713_ (.A1(_15653_),
    .A2(_15654_),
    .B1(_15661_),
    .X(_15662_));
 sky130_fd_sc_hd__nand3_2 _37714_ (.A(_15653_),
    .B(_15654_),
    .C(_15661_),
    .Y(_15663_));
 sky130_fd_sc_hd__a21bo_2 _37715_ (.A1(_15382_),
    .A2(_15381_),
    .B1_N(_15378_),
    .X(_15664_));
 sky130_fd_sc_hd__a21oi_2 _37716_ (.A1(_15662_),
    .A2(_15663_),
    .B1(_15664_),
    .Y(_15665_));
 sky130_fd_sc_hd__and3_2 _37717_ (.A(_15662_),
    .B(_15664_),
    .C(_15663_),
    .X(_15666_));
 sky130_fd_sc_hd__o21a_2 _37718_ (.A1(_15418_),
    .A2(_15410_),
    .B1(_15422_),
    .X(_15667_));
 sky130_fd_sc_hd__o21a_2 _37719_ (.A1(_15665_),
    .A2(_15666_),
    .B1(_15667_),
    .X(_15668_));
 sky130_fd_sc_hd__nor3_2 _37720_ (.A(_15667_),
    .B(_15665_),
    .C(_15666_),
    .Y(_15669_));
 sky130_fd_sc_hd__o2bb2ai_2 _37721_ (.A1_N(_15641_),
    .A2_N(_15645_),
    .B1(_15668_),
    .B2(_15669_),
    .Y(_15670_));
 sky130_fd_sc_hd__nor2_2 _37722_ (.A(_15669_),
    .B(_15668_),
    .Y(_15671_));
 sky130_fd_sc_hd__nand3_2 _37723_ (.A(_15671_),
    .B(_15645_),
    .C(_15641_),
    .Y(_15672_));
 sky130_fd_sc_hd__nand2_2 _37724_ (.A(_15433_),
    .B(_15392_),
    .Y(_15673_));
 sky130_fd_sc_hd__nand2_2 _37725_ (.A(_15673_),
    .B(_15398_),
    .Y(_15674_));
 sky130_fd_sc_hd__a21oi_2 _37726_ (.A1(_15670_),
    .A2(_15672_),
    .B1(_15674_),
    .Y(_15675_));
 sky130_fd_sc_hd__nand3_2 _37727_ (.A(_15670_),
    .B(_15672_),
    .C(_15674_),
    .Y(_15676_));
 sky130_fd_sc_hd__inv_2 _37728_ (.A(_15676_),
    .Y(_15677_));
 sky130_fd_sc_hd__o22ai_2 _37729_ (.A1(_15599_),
    .A2(_15601_),
    .B1(_15675_),
    .B2(_15677_),
    .Y(_15678_));
 sky130_fd_sc_hd__nand2_2 _37730_ (.A(_15670_),
    .B(_15672_),
    .Y(_15679_));
 sky130_fd_sc_hd__inv_2 _37731_ (.A(_15674_),
    .Y(_15680_));
 sky130_fd_sc_hd__nand2_2 _37732_ (.A(_15598_),
    .B(_15600_),
    .Y(_15681_));
 sky130_fd_sc_hd__a21oi_2 _37733_ (.A1(_15679_),
    .A2(_15680_),
    .B1(_15681_),
    .Y(_15682_));
 sky130_fd_sc_hd__nand2_2 _37734_ (.A(_15682_),
    .B(_15676_),
    .Y(_15683_));
 sky130_fd_sc_hd__nand3b_2 _37735_ (.A_N(_15561_),
    .B(_15678_),
    .C(_15683_),
    .Y(_15684_));
 sky130_fd_sc_hd__o21bai_2 _37736_ (.A1(_15675_),
    .A2(_15677_),
    .B1_N(_15681_),
    .Y(_15685_));
 sky130_fd_sc_hd__nand3b_2 _37737_ (.A_N(_15675_),
    .B(_15676_),
    .C(_15681_),
    .Y(_15686_));
 sky130_fd_sc_hd__nand3_2 _37738_ (.A(_15685_),
    .B(_15561_),
    .C(_15686_),
    .Y(_15687_));
 sky130_fd_sc_hd__nand2_2 _37739_ (.A(_15684_),
    .B(_15687_),
    .Y(_15688_));
 sky130_fd_sc_hd__nand2_2 _37740_ (.A(_15492_),
    .B(_15486_),
    .Y(_15689_));
 sky130_fd_sc_hd__or2_2 _37741_ (.A(_15470_),
    .B(_15473_),
    .X(_15690_));
 sky130_fd_sc_hd__inv_2 _37742_ (.A(_15690_),
    .Y(_15691_));
 sky130_fd_sc_hd__nor2_2 _37743_ (.A(_14488_),
    .B(_14755_),
    .Y(_15692_));
 sky130_fd_sc_hd__o31ai_2 _37744_ (.A1(_15470_),
    .A2(_15692_),
    .A3(_15135_),
    .B1(_15502_),
    .Y(_15693_));
 sky130_fd_sc_hd__or2_2 _37745_ (.A(_15691_),
    .B(_15693_),
    .X(_15694_));
 sky130_fd_sc_hd__nand2_2 _37746_ (.A(_15693_),
    .B(_15691_),
    .Y(_15695_));
 sky130_fd_sc_hd__a21o_2 _37747_ (.A1(_15694_),
    .A2(_15695_),
    .B1(_13405_),
    .X(_15696_));
 sky130_fd_sc_hd__nand3_2 _37748_ (.A(_15694_),
    .B(_13406_),
    .C(_15695_),
    .Y(_15697_));
 sky130_fd_sc_hd__nand2_2 _37749_ (.A(_15696_),
    .B(_15697_),
    .Y(_15698_));
 sky130_fd_sc_hd__a21o_2 _37750_ (.A1(_15689_),
    .A2(_15486_),
    .B1(_15698_),
    .X(_15699_));
 sky130_fd_sc_hd__nand3_2 _37751_ (.A(_15689_),
    .B(_15698_),
    .C(_15486_),
    .Y(_15700_));
 sky130_fd_sc_hd__a21bo_2 _37752_ (.A1(_15508_),
    .A2(_14248_),
    .B1_N(_15509_),
    .X(_15701_));
 sky130_fd_sc_hd__and2_2 _37753_ (.A(_15700_),
    .B(_15701_),
    .X(_15702_));
 sky130_fd_sc_hd__a21oi_2 _37754_ (.A1(_15699_),
    .A2(_15700_),
    .B1(_15701_),
    .Y(_15703_));
 sky130_fd_sc_hd__a21oi_2 _37755_ (.A1(_15699_),
    .A2(_15702_),
    .B1(_15703_),
    .Y(_15704_));
 sky130_fd_sc_hd__nand2_2 _37756_ (.A(_15688_),
    .B(_15704_),
    .Y(_15705_));
 sky130_fd_sc_hd__nand2_2 _37757_ (.A(_15702_),
    .B(_15699_),
    .Y(_15706_));
 sky130_fd_sc_hd__a21o_2 _37758_ (.A1(_15699_),
    .A2(_15700_),
    .B1(_15701_),
    .X(_15707_));
 sky130_fd_sc_hd__nand2_2 _37759_ (.A(_15706_),
    .B(_15707_),
    .Y(_15708_));
 sky130_fd_sc_hd__nand3_2 _37760_ (.A(_15684_),
    .B(_15687_),
    .C(_15708_),
    .Y(_15709_));
 sky130_fd_sc_hd__a21oi_2 _37761_ (.A1(_15526_),
    .A2(_15520_),
    .B1(_15500_),
    .Y(_15710_));
 sky130_fd_sc_hd__a21oi_2 _37762_ (.A1(_15705_),
    .A2(_15709_),
    .B1(_15710_),
    .Y(_15711_));
 sky130_fd_sc_hd__nand3_2 _37763_ (.A(_15705_),
    .B(_15709_),
    .C(_15710_),
    .Y(_15712_));
 sky130_fd_sc_hd__nand2_2 _37764_ (.A(_15518_),
    .B(_14018_),
    .Y(_15713_));
 sky130_fd_sc_hd__o21a_2 _37765_ (.A1(_15516_),
    .A2(_15523_),
    .B1(_15518_),
    .X(_15714_));
 sky130_fd_sc_hd__or2_2 _37766_ (.A(_14017_),
    .B(_15714_),
    .X(_15715_));
 sky130_fd_sc_hd__o21a_2 _37767_ (.A1(_15524_),
    .A2(_15713_),
    .B1(_15715_),
    .X(_15716_));
 sky130_fd_sc_hd__nand2_2 _37768_ (.A(_15712_),
    .B(_15716_),
    .Y(_15717_));
 sky130_fd_sc_hd__a31oi_2 _37769_ (.A1(_15561_),
    .A2(_15685_),
    .A3(_15686_),
    .B1(_15708_),
    .Y(_15718_));
 sky130_fd_sc_hd__nand2_2 _37770_ (.A(_15718_),
    .B(_15684_),
    .Y(_15719_));
 sky130_fd_sc_hd__nand2_2 _37771_ (.A(_15688_),
    .B(_15708_),
    .Y(_15720_));
 sky130_fd_sc_hd__nand3b_2 _37772_ (.A_N(_15710_),
    .B(_15719_),
    .C(_15720_),
    .Y(_15721_));
 sky130_fd_sc_hd__a21o_2 _37773_ (.A1(_15721_),
    .A2(_15712_),
    .B1(_15716_),
    .X(_15722_));
 sky130_fd_sc_hd__o221ai_2 _37774_ (.A1(_15559_),
    .A2(_15560_),
    .B1(_15711_),
    .B2(_15717_),
    .C1(_15722_),
    .Y(_15723_));
 sky130_fd_sc_hd__o21ai_2 _37775_ (.A1(_15524_),
    .A2(_15713_),
    .B1(_15715_),
    .Y(_15724_));
 sky130_fd_sc_hd__a21o_2 _37776_ (.A1(_15721_),
    .A2(_15712_),
    .B1(_15724_),
    .X(_15725_));
 sky130_fd_sc_hd__nor2_2 _37777_ (.A(_15559_),
    .B(_15560_),
    .Y(_15726_));
 sky130_fd_sc_hd__nand3_2 _37778_ (.A(_15721_),
    .B(_15712_),
    .C(_15724_),
    .Y(_15727_));
 sky130_fd_sc_hd__nand3_2 _37779_ (.A(_15725_),
    .B(_15726_),
    .C(_15727_),
    .Y(_15728_));
 sky130_fd_sc_hd__buf_1 _37780_ (.A(_15320_),
    .X(_15729_));
 sky130_fd_sc_hd__o2bb2ai_2 _37781_ (.A1_N(_15723_),
    .A2_N(_15728_),
    .B1(_15729_),
    .B2(_15535_),
    .Y(_15730_));
 sky130_fd_sc_hd__nand3_2 _37782_ (.A(_15723_),
    .B(_15728_),
    .C(_15543_),
    .Y(_15731_));
 sky130_fd_sc_hd__a21bo_2 _37783_ (.A1(_15108_),
    .A2(_15541_),
    .B1_N(_15547_),
    .X(_15732_));
 sky130_fd_sc_hd__a21oi_2 _37784_ (.A1(_15730_),
    .A2(_15731_),
    .B1(_15732_),
    .Y(_15733_));
 sky130_fd_sc_hd__and3_2 _37785_ (.A(_15730_),
    .B(_15732_),
    .C(_15731_),
    .X(_15734_));
 sky130_fd_sc_hd__nor2_2 _37786_ (.A(_15733_),
    .B(_15734_),
    .Y(_15735_));
 sky130_fd_sc_hd__a21oi_2 _37787_ (.A1(_15315_),
    .A2(_15319_),
    .B1(_15083_),
    .Y(_15736_));
 sky130_fd_sc_hd__nand2_2 _37788_ (.A(_15325_),
    .B(_15323_),
    .Y(_15737_));
 sky130_fd_sc_hd__o2111ai_2 _37789_ (.A1(_15736_),
    .A2(_15737_),
    .B1(_15556_),
    .C1(_15553_),
    .D1(_15326_),
    .Y(_15738_));
 sky130_fd_sc_hd__nor3_2 _37790_ (.A(_15332_),
    .B(_15738_),
    .C(_14842_),
    .Y(_15739_));
 sky130_fd_sc_hd__nand3_2 _37791_ (.A(_11157_),
    .B(_13760_),
    .C(_15739_),
    .Y(_15740_));
 sky130_fd_sc_hd__nor2_2 _37792_ (.A(_15332_),
    .B(_15738_),
    .Y(_15741_));
 sky130_fd_sc_hd__a21oi_2 _37793_ (.A1(_15554_),
    .A2(_15555_),
    .B1(_15552_),
    .Y(_15742_));
 sky130_fd_sc_hd__o21a_2 _37794_ (.A1(_15327_),
    .A2(_15742_),
    .B1(_15556_),
    .X(_15743_));
 sky130_fd_sc_hd__o21ai_2 _37795_ (.A1(_15335_),
    .A2(_15738_),
    .B1(_15743_),
    .Y(_15744_));
 sky130_fd_sc_hd__a21oi_2 _37796_ (.A1(_15741_),
    .A2(_14849_),
    .B1(_15744_),
    .Y(_15745_));
 sky130_fd_sc_hd__nand2_2 _37797_ (.A(_13765_),
    .B(_15739_),
    .Y(_15746_));
 sky130_fd_sc_hd__nand3_2 _37798_ (.A(_15740_),
    .B(_15745_),
    .C(_15746_),
    .Y(_15747_));
 sky130_fd_sc_hd__xor2_2 _37799_ (.A(_15735_),
    .B(_15747_),
    .X(_02667_));
 sky130_fd_sc_hd__nand2_2 _37800_ (.A(_15589_),
    .B(_15596_),
    .Y(_15748_));
 sky130_fd_sc_hd__nand2_2 _37801_ (.A(_15691_),
    .B(_15692_),
    .Y(_15749_));
 sky130_fd_sc_hd__inv_2 _37802_ (.A(_15502_),
    .Y(_15750_));
 sky130_fd_sc_hd__nand2_2 _37803_ (.A(_15690_),
    .B(_15750_),
    .Y(_15751_));
 sky130_fd_sc_hd__nand2_2 _37804_ (.A(_15749_),
    .B(_15751_),
    .Y(_15752_));
 sky130_fd_sc_hd__nor2_2 _37805_ (.A(_13405_),
    .B(_15752_),
    .Y(_15753_));
 sky130_fd_sc_hd__nand2_2 _37806_ (.A(_15752_),
    .B(_13405_),
    .Y(_15754_));
 sky130_fd_sc_hd__or2b_2 _37807_ (.A(_15753_),
    .B_N(_15754_),
    .X(_15755_));
 sky130_fd_sc_hd__buf_1 _37808_ (.A(_15755_),
    .X(_15756_));
 sky130_fd_sc_hd__a21o_2 _37809_ (.A1(_15748_),
    .A2(_15592_),
    .B1(_15756_),
    .X(_15757_));
 sky130_fd_sc_hd__nand3_2 _37810_ (.A(_15748_),
    .B(_15756_),
    .C(_15592_),
    .Y(_15758_));
 sky130_fd_sc_hd__nand2_2 _37811_ (.A(_15757_),
    .B(_15758_),
    .Y(_15759_));
 sky130_fd_sc_hd__nand2_2 _37812_ (.A(_15696_),
    .B(_15751_),
    .Y(_15760_));
 sky130_fd_sc_hd__inv_2 _37813_ (.A(_15760_),
    .Y(_15761_));
 sky130_fd_sc_hd__nand2_2 _37814_ (.A(_15759_),
    .B(_15761_),
    .Y(_15762_));
 sky130_fd_sc_hd__inv_2 _37815_ (.A(_15762_),
    .Y(_15763_));
 sky130_fd_sc_hd__nand3_2 _37816_ (.A(_15757_),
    .B(_15760_),
    .C(_15758_),
    .Y(_15764_));
 sky130_fd_sc_hd__inv_2 _37817_ (.A(_15764_),
    .Y(_15765_));
 sky130_fd_sc_hd__and4_2 _37818_ (.A(_07832_),
    .B(_14356_),
    .C(_19308_),
    .D(_08950_),
    .X(_15766_));
 sky130_fd_sc_hd__o22a_2 _37819_ (.A1(_07380_),
    .A2(_18182_),
    .B1(_14855_),
    .B2(_08604_),
    .X(_15767_));
 sky130_fd_sc_hd__nor2_2 _37820_ (.A(_15766_),
    .B(_15767_),
    .Y(_15768_));
 sky130_fd_sc_hd__nand3_2 _37821_ (.A(_15768_),
    .B(_19313_),
    .C(_19583_),
    .Y(_15769_));
 sky130_fd_sc_hd__nand2_2 _37822_ (.A(_19313_),
    .B(_19583_),
    .Y(_15770_));
 sky130_fd_sc_hd__o21ai_2 _37823_ (.A1(_15766_),
    .A2(_15767_),
    .B1(_15770_),
    .Y(_15771_));
 sky130_fd_sc_hd__nand2_2 _37824_ (.A(_15769_),
    .B(_15771_),
    .Y(_15772_));
 sky130_fd_sc_hd__inv_2 _37825_ (.A(_15602_),
    .Y(_15773_));
 sky130_fd_sc_hd__o21ai_2 _37826_ (.A1(_15606_),
    .A2(_15603_),
    .B1(_15773_),
    .Y(_15774_));
 sky130_fd_sc_hd__inv_2 _37827_ (.A(_15774_),
    .Y(_15775_));
 sky130_fd_sc_hd__nand2_2 _37828_ (.A(_15772_),
    .B(_15775_),
    .Y(_15776_));
 sky130_fd_sc_hd__nand3_2 _37829_ (.A(_15769_),
    .B(_15771_),
    .C(_15774_),
    .Y(_15777_));
 sky130_fd_sc_hd__buf_1 _37830_ (.A(_19324_),
    .X(_15778_));
 sky130_fd_sc_hd__nand2_2 _37831_ (.A(_15778_),
    .B(_19575_),
    .Y(_15779_));
 sky130_fd_sc_hd__inv_2 _37832_ (.A(_10703_),
    .Y(_15780_));
 sky130_fd_sc_hd__buf_1 _37833_ (.A(_15780_),
    .X(_15781_));
 sky130_fd_sc_hd__o22a_2 _37834_ (.A1(_14370_),
    .A2(_09256_),
    .B1(_14868_),
    .B2(_09678_),
    .X(_15782_));
 sky130_fd_sc_hd__a31o_2 _37835_ (.A1(_19579_),
    .A2(_19581_),
    .A3(_15781_),
    .B1(_15782_),
    .X(_15783_));
 sky130_fd_sc_hd__xor2_2 _37836_ (.A(_15779_),
    .B(_15783_),
    .X(_15784_));
 sky130_fd_sc_hd__a21o_2 _37837_ (.A1(_15776_),
    .A2(_15777_),
    .B1(_15784_),
    .X(_15785_));
 sky130_fd_sc_hd__nand3_2 _37838_ (.A(_15784_),
    .B(_15776_),
    .C(_15777_),
    .Y(_15786_));
 sky130_fd_sc_hd__nand2_2 _37839_ (.A(_15622_),
    .B(_15610_),
    .Y(_15787_));
 sky130_fd_sc_hd__a21oi_2 _37840_ (.A1(_15785_),
    .A2(_15786_),
    .B1(_15787_),
    .Y(_15788_));
 sky130_fd_sc_hd__a21boi_2 _37841_ (.A1(_15609_),
    .A2(_15616_),
    .B1_N(_15610_),
    .Y(_15789_));
 sky130_fd_sc_hd__a21oi_2 _37842_ (.A1(_15776_),
    .A2(_15777_),
    .B1(_15784_),
    .Y(_15790_));
 sky130_fd_sc_hd__nor3b_2 _37843_ (.A(_15789_),
    .B(_15790_),
    .C_N(_15786_),
    .Y(_15791_));
 sky130_fd_sc_hd__o21a_2 _37844_ (.A1(_15624_),
    .A2(_15625_),
    .B1(_15628_),
    .X(_15792_));
 sky130_fd_sc_hd__nor2_2 _37845_ (.A(_14339_),
    .B(_15159_),
    .Y(_15793_));
 sky130_fd_sc_hd__nand2_2 _37846_ (.A(_10166_),
    .B(_09199_),
    .Y(_15794_));
 sky130_fd_sc_hd__nand2_2 _37847_ (.A(_19331_),
    .B(_19567_),
    .Y(_15795_));
 sky130_fd_sc_hd__nor2_2 _37848_ (.A(_15794_),
    .B(_15795_),
    .Y(_15796_));
 sky130_fd_sc_hd__and2_2 _37849_ (.A(_15794_),
    .B(_15795_),
    .X(_15797_));
 sky130_fd_sc_hd__nor2_2 _37850_ (.A(_15796_),
    .B(_15797_),
    .Y(_15798_));
 sky130_fd_sc_hd__or2_2 _37851_ (.A(_15793_),
    .B(_15798_),
    .X(_15799_));
 sky130_fd_sc_hd__nand2_2 _37852_ (.A(_15798_),
    .B(_15793_),
    .Y(_15800_));
 sky130_fd_sc_hd__a31o_2 _37853_ (.A1(_19581_),
    .A2(_19583_),
    .A3(_15781_),
    .B1(_15613_),
    .X(_15801_));
 sky130_fd_sc_hd__a21oi_2 _37854_ (.A1(_15799_),
    .A2(_15800_),
    .B1(_15801_),
    .Y(_15802_));
 sky130_fd_sc_hd__nand3_2 _37855_ (.A(_15801_),
    .B(_15799_),
    .C(_15800_),
    .Y(_15803_));
 sky130_fd_sc_hd__inv_2 _37856_ (.A(_15803_),
    .Y(_15804_));
 sky130_fd_sc_hd__nor3_2 _37857_ (.A(_15792_),
    .B(_15802_),
    .C(_15804_),
    .Y(_15805_));
 sky130_fd_sc_hd__o21a_2 _37858_ (.A1(_15802_),
    .A2(_15804_),
    .B1(_15792_),
    .X(_15806_));
 sky130_fd_sc_hd__nor2_2 _37859_ (.A(_15805_),
    .B(_15806_),
    .Y(_15807_));
 sky130_fd_sc_hd__o21ai_2 _37860_ (.A1(_15788_),
    .A2(_15791_),
    .B1(_15807_),
    .Y(_15808_));
 sky130_fd_sc_hd__a21oi_2 _37861_ (.A1(_15621_),
    .A2(_15622_),
    .B1(_15619_),
    .Y(_15809_));
 sky130_fd_sc_hd__o21a_2 _37862_ (.A1(_15637_),
    .A2(_15809_),
    .B1(_15623_),
    .X(_15810_));
 sky130_fd_sc_hd__nand2_2 _37863_ (.A(_15785_),
    .B(_15786_),
    .Y(_15811_));
 sky130_fd_sc_hd__nand2_2 _37864_ (.A(_15811_),
    .B(_15789_),
    .Y(_15812_));
 sky130_fd_sc_hd__nand3_2 _37865_ (.A(_15785_),
    .B(_15787_),
    .C(_15786_),
    .Y(_15813_));
 sky130_fd_sc_hd__o21ai_2 _37866_ (.A1(_15802_),
    .A2(_15804_),
    .B1(_15792_),
    .Y(_15814_));
 sky130_fd_sc_hd__a21o_2 _37867_ (.A1(_15799_),
    .A2(_15800_),
    .B1(_15801_),
    .X(_15815_));
 sky130_fd_sc_hd__nand3b_2 _37868_ (.A_N(_15792_),
    .B(_15815_),
    .C(_15803_),
    .Y(_15816_));
 sky130_fd_sc_hd__nand2_2 _37869_ (.A(_15814_),
    .B(_15816_),
    .Y(_15817_));
 sky130_fd_sc_hd__nand3_2 _37870_ (.A(_15812_),
    .B(_15813_),
    .C(_15817_),
    .Y(_15818_));
 sky130_fd_sc_hd__nand3_2 _37871_ (.A(_15808_),
    .B(_15810_),
    .C(_15818_),
    .Y(_15819_));
 sky130_fd_sc_hd__o22ai_2 _37872_ (.A1(_15806_),
    .A2(_15805_),
    .B1(_15788_),
    .B2(_15791_),
    .Y(_15820_));
 sky130_fd_sc_hd__o21ai_2 _37873_ (.A1(_15637_),
    .A2(_15809_),
    .B1(_15623_),
    .Y(_15821_));
 sky130_fd_sc_hd__nand3_2 _37874_ (.A(_15812_),
    .B(_15807_),
    .C(_15813_),
    .Y(_15822_));
 sky130_fd_sc_hd__nand3_2 _37875_ (.A(_15820_),
    .B(_15821_),
    .C(_15822_),
    .Y(_15823_));
 sky130_fd_sc_hd__nand2_2 _37876_ (.A(_15819_),
    .B(_15823_),
    .Y(_15824_));
 sky130_fd_sc_hd__a21boi_2 _37877_ (.A1(_15632_),
    .A2(_15634_),
    .B1_N(_15633_),
    .Y(_15825_));
 sky130_fd_sc_hd__nand2_2 _37878_ (.A(_10193_),
    .B(_09220_),
    .Y(_15826_));
 sky130_fd_sc_hd__nand2_2 _37879_ (.A(_08799_),
    .B(_19558_),
    .Y(_15827_));
 sky130_fd_sc_hd__xor2_2 _37880_ (.A(_15826_),
    .B(_15827_),
    .X(_15828_));
 sky130_fd_sc_hd__a21o_2 _37881_ (.A1(_19344_),
    .A2(_19555_),
    .B1(_15828_),
    .X(_15829_));
 sky130_fd_sc_hd__nand3_2 _37882_ (.A(_15828_),
    .B(_19344_),
    .C(_19555_),
    .Y(_15830_));
 sky130_fd_sc_hd__o21ai_2 _37883_ (.A1(_15646_),
    .A2(_15648_),
    .B1(_15650_),
    .Y(_15831_));
 sky130_fd_sc_hd__a21o_2 _37884_ (.A1(_15829_),
    .A2(_15830_),
    .B1(_15831_),
    .X(_15832_));
 sky130_fd_sc_hd__nand3_2 _37885_ (.A(_15831_),
    .B(_15829_),
    .C(_15830_),
    .Y(_15833_));
 sky130_fd_sc_hd__nor2_2 _37886_ (.A(_07053_),
    .B(_10519_),
    .Y(_15834_));
 sky130_fd_sc_hd__a22o_2 _37887_ (.A1(_19348_),
    .A2(_10371_),
    .B1(_19351_),
    .B2(_11038_),
    .X(_15835_));
 sky130_fd_sc_hd__o21ai_2 _37888_ (.A1(_10539_),
    .A2(_15414_),
    .B1(_15835_),
    .Y(_15836_));
 sky130_fd_sc_hd__or2_2 _37889_ (.A(_15834_),
    .B(_15836_),
    .X(_15837_));
 sky130_fd_sc_hd__nand2_2 _37890_ (.A(_15836_),
    .B(_15834_),
    .Y(_15838_));
 sky130_fd_sc_hd__nand2_2 _37891_ (.A(_15837_),
    .B(_15838_),
    .Y(_15839_));
 sky130_fd_sc_hd__a21o_2 _37892_ (.A1(_15832_),
    .A2(_15833_),
    .B1(_15839_),
    .X(_15840_));
 sky130_fd_sc_hd__nand3_2 _37893_ (.A(_15832_),
    .B(_15833_),
    .C(_15839_),
    .Y(_15841_));
 sky130_fd_sc_hd__nand3b_2 _37894_ (.A_N(_15825_),
    .B(_15840_),
    .C(_15841_),
    .Y(_15842_));
 sky130_fd_sc_hd__a21bo_2 _37895_ (.A1(_15832_),
    .A2(_15833_),
    .B1_N(_15839_),
    .X(_15843_));
 sky130_fd_sc_hd__nand3b_2 _37896_ (.A_N(_15839_),
    .B(_15832_),
    .C(_15833_),
    .Y(_15844_));
 sky130_fd_sc_hd__nand3_2 _37897_ (.A(_15843_),
    .B(_15825_),
    .C(_15844_),
    .Y(_15845_));
 sky130_fd_sc_hd__nand2_2 _37898_ (.A(_15663_),
    .B(_15654_),
    .Y(_15846_));
 sky130_fd_sc_hd__a21o_2 _37899_ (.A1(_15842_),
    .A2(_15845_),
    .B1(_15846_),
    .X(_15847_));
 sky130_fd_sc_hd__nand3_2 _37900_ (.A(_15842_),
    .B(_15845_),
    .C(_15846_),
    .Y(_15848_));
 sky130_fd_sc_hd__and2_2 _37901_ (.A(_15847_),
    .B(_15848_),
    .X(_15849_));
 sky130_fd_sc_hd__nand2_2 _37902_ (.A(_15824_),
    .B(_15849_),
    .Y(_15850_));
 sky130_fd_sc_hd__a21oi_2 _37903_ (.A1(_15638_),
    .A2(_15640_),
    .B1(_15639_),
    .Y(_15851_));
 sky130_fd_sc_hd__a21oi_2 _37904_ (.A1(_15671_),
    .A2(_15641_),
    .B1(_15851_),
    .Y(_15852_));
 sky130_fd_sc_hd__nand2_2 _37905_ (.A(_15847_),
    .B(_15848_),
    .Y(_15853_));
 sky130_fd_sc_hd__nand3_2 _37906_ (.A(_15819_),
    .B(_15823_),
    .C(_15853_),
    .Y(_15854_));
 sky130_fd_sc_hd__nand3_2 _37907_ (.A(_15850_),
    .B(_15852_),
    .C(_15854_),
    .Y(_15855_));
 sky130_fd_sc_hd__a21o_2 _37908_ (.A1(_15671_),
    .A2(_15641_),
    .B1(_15851_),
    .X(_15856_));
 sky130_fd_sc_hd__nand2_2 _37909_ (.A(_15824_),
    .B(_15853_),
    .Y(_15857_));
 sky130_fd_sc_hd__nand3_2 _37910_ (.A(_15849_),
    .B(_15819_),
    .C(_15823_),
    .Y(_15858_));
 sky130_fd_sc_hd__nand3_2 _37911_ (.A(_15856_),
    .B(_15857_),
    .C(_15858_),
    .Y(_15859_));
 sky130_fd_sc_hd__nand3_2 _37912_ (.A(_15662_),
    .B(_15664_),
    .C(_15663_),
    .Y(_15860_));
 sky130_fd_sc_hd__o21ai_2 _37913_ (.A1(_15667_),
    .A2(_15665_),
    .B1(_15860_),
    .Y(_15861_));
 sky130_fd_sc_hd__o21ai_2 _37914_ (.A1(_08182_),
    .A2(_19357_),
    .B1(_18156_),
    .Y(_15862_));
 sky130_fd_sc_hd__nor2_2 _37915_ (.A(_15564_),
    .B(_06826_),
    .Y(_15863_));
 sky130_fd_sc_hd__o21ai_2 _37916_ (.A1(_15862_),
    .A2(_15863_),
    .B1(_15451_),
    .Y(_15864_));
 sky130_fd_sc_hd__nor2_2 _37917_ (.A(_08352_),
    .B(_15862_),
    .Y(_15865_));
 sky130_fd_sc_hd__o21ai_2 _37918_ (.A1(_06826_),
    .A2(_15564_),
    .B1(_15865_),
    .Y(_15866_));
 sky130_fd_sc_hd__o21ai_2 _37919_ (.A1(_15414_),
    .A2(_15656_),
    .B1(_15659_),
    .Y(_15867_));
 sky130_fd_sc_hd__a21o_2 _37920_ (.A1(_15864_),
    .A2(_15866_),
    .B1(_15867_),
    .X(_15868_));
 sky130_fd_sc_hd__and2_2 _37921_ (.A(_15864_),
    .B(_15866_),
    .X(_15869_));
 sky130_fd_sc_hd__nand2_2 _37922_ (.A(_15867_),
    .B(_15869_),
    .Y(_15870_));
 sky130_fd_sc_hd__nand2_2 _37923_ (.A(_15868_),
    .B(_15870_),
    .Y(_15871_));
 sky130_fd_sc_hd__nand2_2 _37924_ (.A(_15568_),
    .B(_15569_),
    .Y(_15872_));
 sky130_fd_sc_hd__nand2_2 _37925_ (.A(_15871_),
    .B(_15872_),
    .Y(_15873_));
 sky130_fd_sc_hd__and2_2 _37926_ (.A(_15576_),
    .B(_15574_),
    .X(_15874_));
 sky130_fd_sc_hd__inv_2 _37927_ (.A(_15872_),
    .Y(_15875_));
 sky130_fd_sc_hd__nand3_2 _37928_ (.A(_15868_),
    .B(_15875_),
    .C(_15870_),
    .Y(_15876_));
 sky130_fd_sc_hd__nand3_2 _37929_ (.A(_15873_),
    .B(_15874_),
    .C(_15876_),
    .Y(_15877_));
 sky130_fd_sc_hd__nand2_2 _37930_ (.A(_15871_),
    .B(_15875_),
    .Y(_15878_));
 sky130_fd_sc_hd__nand3_2 _37931_ (.A(_15868_),
    .B(_15872_),
    .C(_15870_),
    .Y(_15879_));
 sky130_fd_sc_hd__nand2_2 _37932_ (.A(_15576_),
    .B(_15574_),
    .Y(_15880_));
 sky130_fd_sc_hd__nand3_2 _37933_ (.A(_15878_),
    .B(_15879_),
    .C(_15880_),
    .Y(_15881_));
 sky130_fd_sc_hd__nand2_2 _37934_ (.A(_15877_),
    .B(_15881_),
    .Y(_15882_));
 sky130_fd_sc_hd__nand2_2 _37935_ (.A(_15882_),
    .B(_15476_),
    .Y(_15883_));
 sky130_fd_sc_hd__nand3_2 _37936_ (.A(_15877_),
    .B(_15881_),
    .C(_15586_),
    .Y(_15884_));
 sky130_fd_sc_hd__nand3b_2 _37937_ (.A_N(_15861_),
    .B(_15883_),
    .C(_15884_),
    .Y(_15885_));
 sky130_fd_sc_hd__buf_1 _37938_ (.A(_15585_),
    .X(_15886_));
 sky130_fd_sc_hd__nand2_2 _37939_ (.A(_15882_),
    .B(_15886_),
    .Y(_15887_));
 sky130_fd_sc_hd__nand3_2 _37940_ (.A(_15877_),
    .B(_15881_),
    .C(_15475_),
    .Y(_15888_));
 sky130_fd_sc_hd__nand3_2 _37941_ (.A(_15887_),
    .B(_15861_),
    .C(_15888_),
    .Y(_15889_));
 sky130_fd_sc_hd__buf_1 _37942_ (.A(_15889_),
    .X(_15890_));
 sky130_fd_sc_hd__nand2_2 _37943_ (.A(_15590_),
    .B(_15583_),
    .Y(_15891_));
 sky130_fd_sc_hd__a21oi_2 _37944_ (.A1(_15885_),
    .A2(_15890_),
    .B1(_15891_),
    .Y(_15892_));
 sky130_fd_sc_hd__and3_2 _37945_ (.A(_15885_),
    .B(_15889_),
    .C(_15891_),
    .X(_15893_));
 sky130_fd_sc_hd__o2bb2ai_2 _37946_ (.A1_N(_15855_),
    .A2_N(_15859_),
    .B1(_15892_),
    .B2(_15893_),
    .Y(_15894_));
 sky130_fd_sc_hd__nor2_2 _37947_ (.A(_15892_),
    .B(_15893_),
    .Y(_15895_));
 sky130_fd_sc_hd__nand3_2 _37948_ (.A(_15895_),
    .B(_15859_),
    .C(_15855_),
    .Y(_15896_));
 sky130_fd_sc_hd__o21ai_2 _37949_ (.A1(_15681_),
    .A2(_15675_),
    .B1(_15676_),
    .Y(_15897_));
 sky130_fd_sc_hd__a21oi_2 _37950_ (.A1(_15894_),
    .A2(_15896_),
    .B1(_15897_),
    .Y(_15898_));
 sky130_fd_sc_hd__o211a_2 _37951_ (.A1(_15677_),
    .A2(_15682_),
    .B1(_15896_),
    .C1(_15894_),
    .X(_15899_));
 sky130_fd_sc_hd__o22ai_2 _37952_ (.A1(_15763_),
    .A2(_15765_),
    .B1(_15898_),
    .B2(_15899_),
    .Y(_15900_));
 sky130_fd_sc_hd__nand2_2 _37953_ (.A(_15762_),
    .B(_15764_),
    .Y(_15901_));
 sky130_fd_sc_hd__a21o_2 _37954_ (.A1(_15894_),
    .A2(_15896_),
    .B1(_15897_),
    .X(_15902_));
 sky130_fd_sc_hd__nand3_2 _37955_ (.A(_15894_),
    .B(_15897_),
    .C(_15896_),
    .Y(_15903_));
 sky130_fd_sc_hd__nand3b_2 _37956_ (.A_N(_15901_),
    .B(_15902_),
    .C(_15903_),
    .Y(_15904_));
 sky130_fd_sc_hd__nand2_2 _37957_ (.A(_15687_),
    .B(_15704_),
    .Y(_15905_));
 sky130_fd_sc_hd__nand2_2 _37958_ (.A(_15905_),
    .B(_15684_),
    .Y(_15906_));
 sky130_fd_sc_hd__a21oi_2 _37959_ (.A1(_15900_),
    .A2(_15904_),
    .B1(_15906_),
    .Y(_15907_));
 sky130_fd_sc_hd__a21oi_2 _37960_ (.A1(_15685_),
    .A2(_15686_),
    .B1(_15561_),
    .Y(_15908_));
 sky130_fd_sc_hd__o211a_2 _37961_ (.A1(_15908_),
    .A2(_15718_),
    .B1(_15904_),
    .C1(_15900_),
    .X(_15909_));
 sky130_fd_sc_hd__or2b_2 _37962_ (.A(_15702_),
    .B_N(_15699_),
    .X(_15910_));
 sky130_fd_sc_hd__nor2_2 _37963_ (.A(_13737_),
    .B(_15910_),
    .Y(_15911_));
 sky130_fd_sc_hd__and2_2 _37964_ (.A(_15910_),
    .B(_13735_),
    .X(_15912_));
 sky130_fd_sc_hd__buf_1 _37965_ (.A(_15912_),
    .X(_15913_));
 sky130_fd_sc_hd__or2_2 _37966_ (.A(_15911_),
    .B(_15913_),
    .X(_15914_));
 sky130_fd_sc_hd__o21ai_2 _37967_ (.A1(_15907_),
    .A2(_15909_),
    .B1(_15914_),
    .Y(_15915_));
 sky130_fd_sc_hd__nand2_2 _37968_ (.A(_15717_),
    .B(_15721_),
    .Y(_15916_));
 sky130_fd_sc_hd__a21o_2 _37969_ (.A1(_15900_),
    .A2(_15904_),
    .B1(_15906_),
    .X(_15917_));
 sky130_fd_sc_hd__nor2_2 _37970_ (.A(_15911_),
    .B(_15913_),
    .Y(_15918_));
 sky130_fd_sc_hd__nand3_2 _37971_ (.A(_15906_),
    .B(_15900_),
    .C(_15904_),
    .Y(_15919_));
 sky130_fd_sc_hd__nand3_2 _37972_ (.A(_15917_),
    .B(_15918_),
    .C(_15919_),
    .Y(_15920_));
 sky130_fd_sc_hd__nand3_2 _37973_ (.A(_15915_),
    .B(_15916_),
    .C(_15920_),
    .Y(_15921_));
 sky130_fd_sc_hd__o21ai_2 _37974_ (.A1(_15907_),
    .A2(_15909_),
    .B1(_15918_),
    .Y(_15922_));
 sky130_fd_sc_hd__a21oi_2 _37975_ (.A1(_15712_),
    .A2(_15716_),
    .B1(_15711_),
    .Y(_15923_));
 sky130_fd_sc_hd__nand3_2 _37976_ (.A(_15917_),
    .B(_15914_),
    .C(_15919_),
    .Y(_15924_));
 sky130_fd_sc_hd__nand3_2 _37977_ (.A(_15922_),
    .B(_15923_),
    .C(_15924_),
    .Y(_15925_));
 sky130_fd_sc_hd__o2bb2ai_2 _37978_ (.A1_N(_15921_),
    .A2_N(_15925_),
    .B1(_15320_),
    .B2(_15714_),
    .Y(_15926_));
 sky130_fd_sc_hd__inv_2 _37979_ (.A(_15715_),
    .Y(_15927_));
 sky130_fd_sc_hd__nand3_2 _37980_ (.A(_15925_),
    .B(_15921_),
    .C(_15927_),
    .Y(_15928_));
 sky130_fd_sc_hd__nand2_2 _37981_ (.A(_15728_),
    .B(_15543_),
    .Y(_15929_));
 sky130_fd_sc_hd__nand2_2 _37982_ (.A(_15929_),
    .B(_15723_),
    .Y(_15930_));
 sky130_fd_sc_hd__a21oi_2 _37983_ (.A1(_15926_),
    .A2(_15928_),
    .B1(_15930_),
    .Y(_15931_));
 sky130_fd_sc_hd__and3_2 _37984_ (.A(_15930_),
    .B(_15926_),
    .C(_15928_),
    .X(_15932_));
 sky130_fd_sc_hd__nor2_2 _37985_ (.A(_15931_),
    .B(_15932_),
    .Y(_15933_));
 sky130_fd_sc_hd__inv_2 _37986_ (.A(_15747_),
    .Y(_15934_));
 sky130_fd_sc_hd__nand3_2 _37987_ (.A(_15730_),
    .B(_15732_),
    .C(_15731_),
    .Y(_15935_));
 sky130_fd_sc_hd__o21ai_2 _37988_ (.A1(_15733_),
    .A2(_15934_),
    .B1(_15935_),
    .Y(_15936_));
 sky130_fd_sc_hd__xor2_2 _37989_ (.A(_15933_),
    .B(_15936_),
    .X(_02668_));
 sky130_fd_sc_hd__nand2_2 _37990_ (.A(_15902_),
    .B(_15903_),
    .Y(_15937_));
 sky130_fd_sc_hd__a22oi_2 _37991_ (.A1(_15905_),
    .A2(_15684_),
    .B1(_15937_),
    .B2(_15901_),
    .Y(_15938_));
 sky130_fd_sc_hd__a22oi_2 _37992_ (.A1(_15904_),
    .A2(_15938_),
    .B1(_15917_),
    .B2(_15918_),
    .Y(_15939_));
 sky130_fd_sc_hd__nand2_2 _37993_ (.A(_10193_),
    .B(_09736_),
    .Y(_15940_));
 sky130_fd_sc_hd__nand2_2 _37994_ (.A(_08799_),
    .B(_19553_),
    .Y(_15941_));
 sky130_fd_sc_hd__nor2_2 _37995_ (.A(_15940_),
    .B(_15941_),
    .Y(_15942_));
 sky130_fd_sc_hd__inv_2 _37996_ (.A(_15942_),
    .Y(_15943_));
 sky130_fd_sc_hd__nand2_2 _37997_ (.A(_15940_),
    .B(_15941_),
    .Y(_15944_));
 sky130_fd_sc_hd__nor2_2 _37998_ (.A(_12602_),
    .B(_11036_),
    .Y(_15945_));
 sky130_fd_sc_hd__a21o_2 _37999_ (.A1(_15943_),
    .A2(_15944_),
    .B1(_15945_),
    .X(_15946_));
 sky130_fd_sc_hd__nand3_2 _38000_ (.A(_15943_),
    .B(_15945_),
    .C(_15944_),
    .Y(_15947_));
 sky130_fd_sc_hd__o21ai_2 _38001_ (.A1(_15826_),
    .A2(_15827_),
    .B1(_15830_),
    .Y(_15948_));
 sky130_fd_sc_hd__a21o_2 _38002_ (.A1(_15946_),
    .A2(_15947_),
    .B1(_15948_),
    .X(_15949_));
 sky130_fd_sc_hd__nand3_2 _38003_ (.A(_15948_),
    .B(_15946_),
    .C(_15947_),
    .Y(_15950_));
 sky130_fd_sc_hd__nand2_2 _38004_ (.A(_14153_),
    .B(_19352_),
    .Y(_15951_));
 sky130_fd_sc_hd__inv_2 _38005_ (.A(_15951_),
    .Y(_15952_));
 sky130_fd_sc_hd__and4_2 _38006_ (.A(_19347_),
    .B(_08159_),
    .C(_11901_),
    .D(_11037_),
    .X(_15953_));
 sky130_fd_sc_hd__o22a_2 _38007_ (.A1(_12596_),
    .A2(_10535_),
    .B1(_12597_),
    .B2(_10518_),
    .X(_15954_));
 sky130_fd_sc_hd__nor2_2 _38008_ (.A(_15953_),
    .B(_15954_),
    .Y(_15955_));
 sky130_fd_sc_hd__xor2_2 _38009_ (.A(_15952_),
    .B(_15955_),
    .X(_15956_));
 sky130_fd_sc_hd__a21oi_2 _38010_ (.A1(_15949_),
    .A2(_15950_),
    .B1(_15956_),
    .Y(_15957_));
 sky130_fd_sc_hd__and3_2 _38011_ (.A(_15949_),
    .B(_15956_),
    .C(_15950_),
    .X(_15958_));
 sky130_fd_sc_hd__o21ai_2 _38012_ (.A1(_15792_),
    .A2(_15802_),
    .B1(_15803_),
    .Y(_15959_));
 sky130_fd_sc_hd__o21bai_2 _38013_ (.A1(_15957_),
    .A2(_15958_),
    .B1_N(_15959_),
    .Y(_15960_));
 sky130_fd_sc_hd__a21o_2 _38014_ (.A1(_15949_),
    .A2(_15950_),
    .B1(_15956_),
    .X(_15961_));
 sky130_fd_sc_hd__nand3_2 _38015_ (.A(_15949_),
    .B(_15956_),
    .C(_15950_),
    .Y(_15962_));
 sky130_fd_sc_hd__nand3_2 _38016_ (.A(_15961_),
    .B(_15962_),
    .C(_15959_),
    .Y(_15963_));
 sky130_fd_sc_hd__nand2_2 _38017_ (.A(_15832_),
    .B(_15839_),
    .Y(_15964_));
 sky130_fd_sc_hd__nand2_2 _38018_ (.A(_15964_),
    .B(_15833_),
    .Y(_15965_));
 sky130_fd_sc_hd__a21oi_2 _38019_ (.A1(_15960_),
    .A2(_15963_),
    .B1(_15965_),
    .Y(_15966_));
 sky130_fd_sc_hd__and3_2 _38020_ (.A(_15960_),
    .B(_15963_),
    .C(_15965_),
    .X(_15967_));
 sky130_fd_sc_hd__nand2_2 _38021_ (.A(_15786_),
    .B(_15777_),
    .Y(_15968_));
 sky130_fd_sc_hd__a21oi_2 _38022_ (.A1(_19313_),
    .A2(_19583_),
    .B1(_15766_),
    .Y(_15969_));
 sky130_fd_sc_hd__and4_2 _38023_ (.A(_08598_),
    .B(_11169_),
    .C(_10823_),
    .D(_19582_),
    .X(_15970_));
 sky130_fd_sc_hd__o22a_2 _38024_ (.A1(_08950_),
    .A2(_11509_),
    .B1(_10832_),
    .B2(_08947_),
    .X(_15971_));
 sky130_fd_sc_hd__nor2_2 _38025_ (.A(_15970_),
    .B(_15971_),
    .Y(_15972_));
 sky130_fd_sc_hd__nand2_2 _38026_ (.A(_10827_),
    .B(_19581_),
    .Y(_15973_));
 sky130_fd_sc_hd__nand2_2 _38027_ (.A(_15972_),
    .B(_15973_),
    .Y(_15974_));
 sky130_fd_sc_hd__or2_2 _38028_ (.A(_15973_),
    .B(_15972_),
    .X(_15975_));
 sky130_fd_sc_hd__o211ai_2 _38029_ (.A1(_15767_),
    .A2(_15969_),
    .B1(_15974_),
    .C1(_15975_),
    .Y(_15976_));
 sky130_fd_sc_hd__nor2_2 _38030_ (.A(_15770_),
    .B(_15767_),
    .Y(_15977_));
 sky130_fd_sc_hd__o21ai_2 _38031_ (.A1(_15970_),
    .A2(_15971_),
    .B1(_15973_),
    .Y(_15978_));
 sky130_fd_sc_hd__or3_2 _38032_ (.A(_15973_),
    .B(_15970_),
    .C(_15971_),
    .X(_15979_));
 sky130_fd_sc_hd__o211ai_2 _38033_ (.A1(_15766_),
    .A2(_15977_),
    .B1(_15978_),
    .C1(_15979_),
    .Y(_15980_));
 sky130_fd_sc_hd__nand2_2 _38034_ (.A(_19324_),
    .B(_19572_),
    .Y(_15981_));
 sky130_fd_sc_hd__o22a_2 _38035_ (.A1(_14370_),
    .A2(_11660_),
    .B1(_14869_),
    .B2(_14646_),
    .X(_15982_));
 sky130_fd_sc_hd__and3_2 _38036_ (.A(_15780_),
    .B(_12349_),
    .C(_07845_),
    .X(_15983_));
 sky130_fd_sc_hd__nor3_2 _38037_ (.A(_15981_),
    .B(_15982_),
    .C(_15983_),
    .Y(_15984_));
 sky130_fd_sc_hd__o21a_2 _38038_ (.A1(_15982_),
    .A2(_15983_),
    .B1(_15981_),
    .X(_15985_));
 sky130_fd_sc_hd__nor2_2 _38039_ (.A(_15984_),
    .B(_15985_),
    .Y(_15986_));
 sky130_fd_sc_hd__a21o_2 _38040_ (.A1(_15976_),
    .A2(_15980_),
    .B1(_15986_),
    .X(_15987_));
 sky130_fd_sc_hd__nand3_2 _38041_ (.A(_15976_),
    .B(_15986_),
    .C(_15980_),
    .Y(_15988_));
 sky130_fd_sc_hd__nand3_2 _38042_ (.A(_15968_),
    .B(_15987_),
    .C(_15988_),
    .Y(_15989_));
 sky130_fd_sc_hd__a21oi_2 _38043_ (.A1(_15976_),
    .A2(_15980_),
    .B1(_15986_),
    .Y(_15990_));
 sky130_fd_sc_hd__and3_2 _38044_ (.A(_15976_),
    .B(_15986_),
    .C(_15980_),
    .X(_15991_));
 sky130_fd_sc_hd__a21boi_2 _38045_ (.A1(_15784_),
    .A2(_15776_),
    .B1_N(_15777_),
    .Y(_15992_));
 sky130_fd_sc_hd__o21ai_2 _38046_ (.A1(_15990_),
    .A2(_15991_),
    .B1(_15992_),
    .Y(_15993_));
 sky130_fd_sc_hd__inv_2 _38047_ (.A(_15800_),
    .Y(_15994_));
 sky130_fd_sc_hd__nor2_2 _38048_ (.A(_15796_),
    .B(_15994_),
    .Y(_15995_));
 sky130_fd_sc_hd__nand2_2 _38049_ (.A(_19328_),
    .B(_08662_),
    .Y(_15996_));
 sky130_fd_sc_hd__nand2_2 _38050_ (.A(_10156_),
    .B(_10380_),
    .Y(_15997_));
 sky130_fd_sc_hd__or2_2 _38051_ (.A(_15996_),
    .B(_15997_),
    .X(_15998_));
 sky130_fd_sc_hd__nand2_2 _38052_ (.A(_15996_),
    .B(_15997_),
    .Y(_15999_));
 sky130_fd_sc_hd__nand2_2 _38053_ (.A(_19334_),
    .B(_10055_),
    .Y(_16000_));
 sky130_fd_sc_hd__a21bo_2 _38054_ (.A1(_15998_),
    .A2(_15999_),
    .B1_N(_16000_),
    .X(_16001_));
 sky130_fd_sc_hd__nand3b_2 _38055_ (.A_N(_16000_),
    .B(_15998_),
    .C(_15999_),
    .Y(_16002_));
 sky130_fd_sc_hd__buf_1 _38056_ (.A(_11178_),
    .X(_16003_));
 sky130_fd_sc_hd__o32ai_2 _38057_ (.A1(_09679_),
    .A2(_09263_),
    .A3(_16003_),
    .B1(_15779_),
    .B2(_15782_),
    .Y(_16004_));
 sky130_fd_sc_hd__a21o_2 _38058_ (.A1(_16001_),
    .A2(_16002_),
    .B1(_16004_),
    .X(_16005_));
 sky130_fd_sc_hd__nand3_2 _38059_ (.A(_16001_),
    .B(_16004_),
    .C(_16002_),
    .Y(_16006_));
 sky130_fd_sc_hd__nand2_2 _38060_ (.A(_16005_),
    .B(_16006_),
    .Y(_16007_));
 sky130_fd_sc_hd__nor2_2 _38061_ (.A(_15995_),
    .B(_16007_),
    .Y(_16008_));
 sky130_fd_sc_hd__inv_2 _38062_ (.A(_15995_),
    .Y(_16009_));
 sky130_fd_sc_hd__and2_2 _38063_ (.A(_16005_),
    .B(_16006_),
    .X(_16010_));
 sky130_fd_sc_hd__nor2_2 _38064_ (.A(_16009_),
    .B(_16010_),
    .Y(_16011_));
 sky130_fd_sc_hd__o2bb2ai_2 _38065_ (.A1_N(_15989_),
    .A2_N(_15993_),
    .B1(_16008_),
    .B2(_16011_),
    .Y(_16012_));
 sky130_fd_sc_hd__nor2_2 _38066_ (.A(_16008_),
    .B(_16011_),
    .Y(_16013_));
 sky130_fd_sc_hd__nand3_2 _38067_ (.A(_15993_),
    .B(_16013_),
    .C(_15989_),
    .Y(_16014_));
 sky130_fd_sc_hd__o21ai_2 _38068_ (.A1(_15817_),
    .A2(_15788_),
    .B1(_15813_),
    .Y(_16015_));
 sky130_fd_sc_hd__a21oi_2 _38069_ (.A1(_16012_),
    .A2(_16014_),
    .B1(_16015_),
    .Y(_16016_));
 sky130_fd_sc_hd__a21oi_2 _38070_ (.A1(_15811_),
    .A2(_15789_),
    .B1(_15817_),
    .Y(_16017_));
 sky130_fd_sc_hd__o211a_2 _38071_ (.A1(_15791_),
    .A2(_16017_),
    .B1(_16014_),
    .C1(_16012_),
    .X(_16018_));
 sky130_fd_sc_hd__o22ai_2 _38072_ (.A1(_15966_),
    .A2(_15967_),
    .B1(_16016_),
    .B2(_16018_),
    .Y(_16019_));
 sky130_fd_sc_hd__a21oi_2 _38073_ (.A1(_15993_),
    .A2(_15989_),
    .B1(_16013_),
    .Y(_16020_));
 sky130_fd_sc_hd__nor2_2 _38074_ (.A(_15995_),
    .B(_16010_),
    .Y(_16021_));
 sky130_fd_sc_hd__nor2_2 _38075_ (.A(_16007_),
    .B(_16009_),
    .Y(_16022_));
 sky130_fd_sc_hd__o211a_2 _38076_ (.A1(_16021_),
    .A2(_16022_),
    .B1(_15989_),
    .C1(_15993_),
    .X(_16023_));
 sky130_fd_sc_hd__o21bai_2 _38077_ (.A1(_16020_),
    .A2(_16023_),
    .B1_N(_16015_),
    .Y(_16024_));
 sky130_fd_sc_hd__nor2_2 _38078_ (.A(_15966_),
    .B(_15967_),
    .Y(_16025_));
 sky130_fd_sc_hd__nand3_2 _38079_ (.A(_16012_),
    .B(_16015_),
    .C(_16014_),
    .Y(_16026_));
 sky130_fd_sc_hd__nand3_2 _38080_ (.A(_16024_),
    .B(_16025_),
    .C(_16026_),
    .Y(_16027_));
 sky130_fd_sc_hd__a21oi_2 _38081_ (.A1(_15820_),
    .A2(_15822_),
    .B1(_15821_),
    .Y(_16028_));
 sky130_fd_sc_hd__a21oi_2 _38082_ (.A1(_15853_),
    .A2(_15823_),
    .B1(_16028_),
    .Y(_16029_));
 sky130_fd_sc_hd__a21oi_2 _38083_ (.A1(_16019_),
    .A2(_16027_),
    .B1(_16029_),
    .Y(_16030_));
 sky130_fd_sc_hd__nand2_2 _38084_ (.A(_16024_),
    .B(_16025_),
    .Y(_16031_));
 sky130_fd_sc_hd__o211a_2 _38085_ (.A1(_16018_),
    .A2(_16031_),
    .B1(_16029_),
    .C1(_16019_),
    .X(_16032_));
 sky130_fd_sc_hd__nand2_2 _38086_ (.A(_15868_),
    .B(_15872_),
    .Y(_16033_));
 sky130_fd_sc_hd__nand2_2 _38087_ (.A(_16033_),
    .B(_15870_),
    .Y(_16034_));
 sky130_fd_sc_hd__a2bb2o_2 _38088_ (.A1_N(_10539_),
    .A2_N(_15414_),
    .B1(_15835_),
    .B2(_15834_),
    .X(_16035_));
 sky130_fd_sc_hd__nor2_2 _38089_ (.A(_16035_),
    .B(_15869_),
    .Y(_16036_));
 sky130_fd_sc_hd__nor2_2 _38090_ (.A(_15863_),
    .B(_15865_),
    .Y(_16037_));
 sky130_fd_sc_hd__inv_2 _38091_ (.A(_16037_),
    .Y(_16038_));
 sky130_fd_sc_hd__nand2_2 _38092_ (.A(_15869_),
    .B(_16035_),
    .Y(_16039_));
 sky130_fd_sc_hd__or3b_2 _38093_ (.A(_16036_),
    .B(_16038_),
    .C_N(_16039_),
    .X(_16040_));
 sky130_fd_sc_hd__inv_2 _38094_ (.A(_16036_),
    .Y(_16041_));
 sky130_fd_sc_hd__nand2_2 _38095_ (.A(_16041_),
    .B(_16039_),
    .Y(_16042_));
 sky130_fd_sc_hd__nand2_2 _38096_ (.A(_16042_),
    .B(_16038_),
    .Y(_16043_));
 sky130_fd_sc_hd__nand3b_2 _38097_ (.A_N(_16034_),
    .B(_16040_),
    .C(_16043_),
    .Y(_16044_));
 sky130_fd_sc_hd__buf_1 _38098_ (.A(_16037_),
    .X(_16045_));
 sky130_fd_sc_hd__or3b_2 _38099_ (.A(_16036_),
    .B(_16045_),
    .C_N(_16039_),
    .X(_16046_));
 sky130_fd_sc_hd__nand2_2 _38100_ (.A(_16042_),
    .B(_16045_),
    .Y(_16047_));
 sky130_fd_sc_hd__nand3_2 _38101_ (.A(_16046_),
    .B(_16034_),
    .C(_16047_),
    .Y(_16048_));
 sky130_fd_sc_hd__nand2_2 _38102_ (.A(_16044_),
    .B(_16048_),
    .Y(_16049_));
 sky130_fd_sc_hd__nand2_2 _38103_ (.A(_16049_),
    .B(_15476_),
    .Y(_16050_));
 sky130_fd_sc_hd__a21boi_2 _38104_ (.A1(_15846_),
    .A2(_15845_),
    .B1_N(_15842_),
    .Y(_16051_));
 sky130_fd_sc_hd__nand3_2 _38105_ (.A(_16044_),
    .B(_16048_),
    .C(_15586_),
    .Y(_16052_));
 sky130_fd_sc_hd__nand3_2 _38106_ (.A(_16050_),
    .B(_16051_),
    .C(_16052_),
    .Y(_16053_));
 sky130_fd_sc_hd__nand2_2 _38107_ (.A(_16049_),
    .B(_15886_),
    .Y(_16054_));
 sky130_fd_sc_hd__nand2_2 _38108_ (.A(_15848_),
    .B(_15842_),
    .Y(_16055_));
 sky130_fd_sc_hd__nand3_2 _38109_ (.A(_16044_),
    .B(_16048_),
    .C(_15478_),
    .Y(_16056_));
 sky130_fd_sc_hd__nand2_2 _38110_ (.A(_15877_),
    .B(_15478_),
    .Y(_16057_));
 sky130_fd_sc_hd__nand2_2 _38111_ (.A(_16057_),
    .B(_15881_),
    .Y(_16058_));
 sky130_fd_sc_hd__inv_2 _38112_ (.A(_16058_),
    .Y(_16059_));
 sky130_fd_sc_hd__a31oi_2 _38113_ (.A1(_16054_),
    .A2(_16055_),
    .A3(_16056_),
    .B1(_16059_),
    .Y(_16060_));
 sky130_fd_sc_hd__nand3_2 _38114_ (.A(_16054_),
    .B(_16055_),
    .C(_16056_),
    .Y(_16061_));
 sky130_fd_sc_hd__a21oi_2 _38115_ (.A1(_16061_),
    .A2(_16053_),
    .B1(_16058_),
    .Y(_16062_));
 sky130_fd_sc_hd__a21oi_2 _38116_ (.A1(_16053_),
    .A2(_16060_),
    .B1(_16062_),
    .Y(_16063_));
 sky130_fd_sc_hd__o21ai_2 _38117_ (.A1(_16030_),
    .A2(_16032_),
    .B1(_16063_),
    .Y(_16064_));
 sky130_fd_sc_hd__a21boi_2 _38118_ (.A1(_15855_),
    .A2(_15895_),
    .B1_N(_15859_),
    .Y(_16065_));
 sky130_fd_sc_hd__and2_2 _38119_ (.A(_15823_),
    .B(_15853_),
    .X(_16066_));
 sky130_fd_sc_hd__o2bb2ai_2 _38120_ (.A1_N(_16027_),
    .A2_N(_16019_),
    .B1(_16028_),
    .B2(_16066_),
    .Y(_16067_));
 sky130_fd_sc_hd__nand2_2 _38121_ (.A(_16061_),
    .B(_16053_),
    .Y(_16068_));
 sky130_fd_sc_hd__nand2_2 _38122_ (.A(_16068_),
    .B(_16059_),
    .Y(_16069_));
 sky130_fd_sc_hd__nand3_2 _38123_ (.A(_16061_),
    .B(_16053_),
    .C(_16058_),
    .Y(_16070_));
 sky130_fd_sc_hd__nand2_2 _38124_ (.A(_16069_),
    .B(_16070_),
    .Y(_16071_));
 sky130_fd_sc_hd__nand3_2 _38125_ (.A(_16019_),
    .B(_16029_),
    .C(_16027_),
    .Y(_16072_));
 sky130_fd_sc_hd__nand3_2 _38126_ (.A(_16067_),
    .B(_16071_),
    .C(_16072_),
    .Y(_16073_));
 sky130_fd_sc_hd__nand3_2 _38127_ (.A(_16064_),
    .B(_16065_),
    .C(_16073_),
    .Y(_16074_));
 sky130_fd_sc_hd__inv_2 _38128_ (.A(_16070_),
    .Y(_16075_));
 sky130_fd_sc_hd__o22ai_2 _38129_ (.A1(_16062_),
    .A2(_16075_),
    .B1(_16030_),
    .B2(_16032_),
    .Y(_16076_));
 sky130_fd_sc_hd__nand2_2 _38130_ (.A(_15895_),
    .B(_15855_),
    .Y(_16077_));
 sky130_fd_sc_hd__nand2_2 _38131_ (.A(_16077_),
    .B(_15859_),
    .Y(_16078_));
 sky130_fd_sc_hd__nand3_2 _38132_ (.A(_16067_),
    .B(_16063_),
    .C(_16072_),
    .Y(_16079_));
 sky130_fd_sc_hd__nand3_2 _38133_ (.A(_16076_),
    .B(_16078_),
    .C(_16079_),
    .Y(_16080_));
 sky130_fd_sc_hd__nand2_2 _38134_ (.A(_16074_),
    .B(_16080_),
    .Y(_16081_));
 sky130_fd_sc_hd__nand3_2 _38135_ (.A(_15885_),
    .B(_15890_),
    .C(_15891_),
    .Y(_16082_));
 sky130_fd_sc_hd__buf_1 _38136_ (.A(_15756_),
    .X(_16083_));
 sky130_fd_sc_hd__a21oi_2 _38137_ (.A1(_16082_),
    .A2(_15890_),
    .B1(_16083_),
    .Y(_16084_));
 sky130_fd_sc_hd__buf_1 _38138_ (.A(_15755_),
    .X(_16085_));
 sky130_fd_sc_hd__and3_2 _38139_ (.A(_16082_),
    .B(_16085_),
    .C(_15890_),
    .X(_16086_));
 sky130_fd_sc_hd__inv_2 _38140_ (.A(_15751_),
    .Y(_16087_));
 sky130_fd_sc_hd__nor2_2 _38141_ (.A(_16087_),
    .B(_15753_),
    .Y(_16088_));
 sky130_fd_sc_hd__buf_1 _38142_ (.A(_16088_),
    .X(_16089_));
 sky130_fd_sc_hd__o21ai_2 _38143_ (.A1(_16084_),
    .A2(_16086_),
    .B1(_16089_),
    .Y(_16090_));
 sky130_fd_sc_hd__a21o_2 _38144_ (.A1(_16082_),
    .A2(_15890_),
    .B1(_16085_),
    .X(_16091_));
 sky130_fd_sc_hd__inv_2 _38145_ (.A(_16088_),
    .Y(_16092_));
 sky130_fd_sc_hd__buf_1 _38146_ (.A(_16092_),
    .X(_16093_));
 sky130_fd_sc_hd__nand3_2 _38147_ (.A(_16082_),
    .B(_16085_),
    .C(_15890_),
    .Y(_16094_));
 sky130_fd_sc_hd__nand3_2 _38148_ (.A(_16091_),
    .B(_16093_),
    .C(_16094_),
    .Y(_16095_));
 sky130_fd_sc_hd__nand2_2 _38149_ (.A(_16090_),
    .B(_16095_),
    .Y(_16096_));
 sky130_fd_sc_hd__nand2_2 _38150_ (.A(_16081_),
    .B(_16096_),
    .Y(_16097_));
 sky130_fd_sc_hd__a31oi_2 _38151_ (.A1(_16064_),
    .A2(_16065_),
    .A3(_16073_),
    .B1(_16096_),
    .Y(_16098_));
 sky130_fd_sc_hd__nand2_2 _38152_ (.A(_16098_),
    .B(_16080_),
    .Y(_16099_));
 sky130_fd_sc_hd__o21ai_2 _38153_ (.A1(_15901_),
    .A2(_15898_),
    .B1(_15903_),
    .Y(_16100_));
 sky130_fd_sc_hd__nand3_2 _38154_ (.A(_16097_),
    .B(_16099_),
    .C(_16100_),
    .Y(_16101_));
 sky130_fd_sc_hd__and2_2 _38155_ (.A(_16090_),
    .B(_16095_),
    .X(_16102_));
 sky130_fd_sc_hd__nand2_2 _38156_ (.A(_16081_),
    .B(_16102_),
    .Y(_16103_));
 sky130_fd_sc_hd__nand2_2 _38157_ (.A(_15903_),
    .B(_15901_),
    .Y(_16104_));
 sky130_fd_sc_hd__nand2_2 _38158_ (.A(_16104_),
    .B(_15902_),
    .Y(_16105_));
 sky130_fd_sc_hd__nand3_2 _38159_ (.A(_16074_),
    .B(_16080_),
    .C(_16096_),
    .Y(_16106_));
 sky130_fd_sc_hd__nand3_2 _38160_ (.A(_16103_),
    .B(_16105_),
    .C(_16106_),
    .Y(_16107_));
 sky130_fd_sc_hd__nand2_2 _38161_ (.A(_15758_),
    .B(_15760_),
    .Y(_16108_));
 sky130_fd_sc_hd__nand2_2 _38162_ (.A(_16108_),
    .B(_15757_),
    .Y(_16109_));
 sky130_fd_sc_hd__nor2_2 _38163_ (.A(_14823_),
    .B(_16109_),
    .Y(_16110_));
 sky130_fd_sc_hd__inv_2 _38164_ (.A(_16109_),
    .Y(_16111_));
 sky130_fd_sc_hd__nor2_2 _38165_ (.A(_13737_),
    .B(_16111_),
    .Y(_16112_));
 sky130_fd_sc_hd__nor2_2 _38166_ (.A(_16110_),
    .B(_16112_),
    .Y(_16113_));
 sky130_fd_sc_hd__nand3_2 _38167_ (.A(_16101_),
    .B(_16107_),
    .C(_16113_),
    .Y(_16114_));
 sky130_fd_sc_hd__o2bb2ai_2 _38168_ (.A1_N(_16107_),
    .A2_N(_16101_),
    .B1(_16110_),
    .B2(_16112_),
    .Y(_16115_));
 sky130_fd_sc_hd__nand3_2 _38169_ (.A(_15939_),
    .B(_16114_),
    .C(_16115_),
    .Y(_16116_));
 sky130_fd_sc_hd__o21ai_2 _38170_ (.A1(_15914_),
    .A2(_15907_),
    .B1(_15919_),
    .Y(_16117_));
 sky130_fd_sc_hd__buf_1 _38171_ (.A(_14018_),
    .X(_16118_));
 sky130_fd_sc_hd__nor2_2 _38172_ (.A(_16118_),
    .B(_16111_),
    .Y(_16119_));
 sky130_fd_sc_hd__buf_1 _38173_ (.A(_15109_),
    .X(_16120_));
 sky130_fd_sc_hd__nor2_2 _38174_ (.A(_16120_),
    .B(_16109_),
    .Y(_16121_));
 sky130_fd_sc_hd__o2bb2ai_2 _38175_ (.A1_N(_16107_),
    .A2_N(_16101_),
    .B1(_16119_),
    .B2(_16121_),
    .Y(_16122_));
 sky130_fd_sc_hd__a31oi_2 _38176_ (.A1(_16103_),
    .A2(_16105_),
    .A3(_16106_),
    .B1(_16113_),
    .Y(_16123_));
 sky130_fd_sc_hd__nand2_2 _38177_ (.A(_16123_),
    .B(_16101_),
    .Y(_16124_));
 sky130_fd_sc_hd__nand3_2 _38178_ (.A(_16117_),
    .B(_16122_),
    .C(_16124_),
    .Y(_16125_));
 sky130_fd_sc_hd__nand2_2 _38179_ (.A(_16116_),
    .B(_16125_),
    .Y(_16126_));
 sky130_fd_sc_hd__nand2_2 _38180_ (.A(_16126_),
    .B(_15913_),
    .Y(_16127_));
 sky130_fd_sc_hd__a21boi_2 _38181_ (.A1(_15925_),
    .A2(_15927_),
    .B1_N(_15921_),
    .Y(_16128_));
 sky130_fd_sc_hd__inv_2 _38182_ (.A(_15913_),
    .Y(_16129_));
 sky130_fd_sc_hd__nand3_2 _38183_ (.A(_16116_),
    .B(_16125_),
    .C(_16129_),
    .Y(_16130_));
 sky130_fd_sc_hd__nand3_2 _38184_ (.A(_16127_),
    .B(_16128_),
    .C(_16130_),
    .Y(_16131_));
 sky130_fd_sc_hd__nand2_2 _38185_ (.A(_16126_),
    .B(_16129_),
    .Y(_16132_));
 sky130_fd_sc_hd__and3_2 _38186_ (.A(_15917_),
    .B(_15918_),
    .C(_15919_),
    .X(_16133_));
 sky130_fd_sc_hd__nand2_2 _38187_ (.A(_15915_),
    .B(_15916_),
    .Y(_16134_));
 sky130_fd_sc_hd__o2bb2ai_2 _38188_ (.A1_N(_15927_),
    .A2_N(_15925_),
    .B1(_16133_),
    .B2(_16134_),
    .Y(_16135_));
 sky130_fd_sc_hd__nand3_2 _38189_ (.A(_16116_),
    .B(_16125_),
    .C(_15913_),
    .Y(_16136_));
 sky130_fd_sc_hd__nand3_2 _38190_ (.A(_16132_),
    .B(_16135_),
    .C(_16136_),
    .Y(_16137_));
 sky130_fd_sc_hd__nand2_2 _38191_ (.A(_16131_),
    .B(_16137_),
    .Y(_16138_));
 sky130_fd_sc_hd__nand3_2 _38192_ (.A(_15930_),
    .B(_15926_),
    .C(_15928_),
    .Y(_16139_));
 sky130_fd_sc_hd__a21oi_2 _38193_ (.A1(_15935_),
    .A2(_16139_),
    .B1(_15931_),
    .Y(_16140_));
 sky130_fd_sc_hd__and3_2 _38194_ (.A(_15747_),
    .B(_15735_),
    .C(_15933_),
    .X(_16141_));
 sky130_fd_sc_hd__nor2_2 _38195_ (.A(_16140_),
    .B(_16141_),
    .Y(_16142_));
 sky130_fd_sc_hd__xor2_2 _38196_ (.A(_16138_),
    .B(_16142_),
    .X(_02669_));
 sky130_fd_sc_hd__o21ai_2 _38197_ (.A1(_16140_),
    .A2(_16141_),
    .B1(_16131_),
    .Y(_16143_));
 sky130_fd_sc_hd__inv_2 _38198_ (.A(_16113_),
    .Y(_16144_));
 sky130_fd_sc_hd__a21oi_2 _38199_ (.A1(_16103_),
    .A2(_16106_),
    .B1(_16105_),
    .Y(_16145_));
 sky130_fd_sc_hd__a21oi_2 _38200_ (.A1(_16107_),
    .A2(_16144_),
    .B1(_16145_),
    .Y(_16146_));
 sky130_fd_sc_hd__a21oi_2 _38201_ (.A1(_16064_),
    .A2(_16073_),
    .B1(_16065_),
    .Y(_16147_));
 sky130_fd_sc_hd__a21oi_2 _38202_ (.A1(_16067_),
    .A2(_16063_),
    .B1(_16032_),
    .Y(_16148_));
 sky130_fd_sc_hd__nor2_2 _38203_ (.A(_15973_),
    .B(_15971_),
    .Y(_16149_));
 sky130_fd_sc_hd__nand2_2 _38204_ (.A(_10827_),
    .B(_19579_),
    .Y(_16150_));
 sky130_fd_sc_hd__and4_2 _38205_ (.A(_08946_),
    .B(_10824_),
    .C(_10823_),
    .D(_08650_),
    .X(_16151_));
 sky130_fd_sc_hd__o22a_2 _38206_ (.A1(_09933_),
    .A2(_10830_),
    .B1(_10832_),
    .B2(_09256_),
    .X(_16152_));
 sky130_fd_sc_hd__nor2_2 _38207_ (.A(_16151_),
    .B(_16152_),
    .Y(_16153_));
 sky130_fd_sc_hd__nor2_2 _38208_ (.A(_16150_),
    .B(_16153_),
    .Y(_16154_));
 sky130_fd_sc_hd__and2_2 _38209_ (.A(_16153_),
    .B(_16150_),
    .X(_16155_));
 sky130_fd_sc_hd__o22ai_2 _38210_ (.A1(_15970_),
    .A2(_16149_),
    .B1(_16154_),
    .B2(_16155_),
    .Y(_16156_));
 sky130_fd_sc_hd__nand2_2 _38211_ (.A(_16153_),
    .B(_16150_),
    .Y(_16157_));
 sky130_fd_sc_hd__nor2_2 _38212_ (.A(_15970_),
    .B(_16149_),
    .Y(_16158_));
 sky130_fd_sc_hd__nand3b_2 _38213_ (.A_N(_16154_),
    .B(_16157_),
    .C(_16158_),
    .Y(_16159_));
 sky130_fd_sc_hd__a22o_2 _38214_ (.A1(_10146_),
    .A2(_09994_),
    .B1(_09838_),
    .B2(_14112_),
    .X(_16160_));
 sky130_fd_sc_hd__o31ai_2 _38215_ (.A1(_10705_),
    .A2(_12090_),
    .A3(_14646_),
    .B1(_16160_),
    .Y(_16161_));
 sky130_fd_sc_hd__a21oi_2 _38216_ (.A1(_19325_),
    .A2(_19569_),
    .B1(_16161_),
    .Y(_16162_));
 sky130_fd_sc_hd__and3_2 _38217_ (.A(_16161_),
    .B(_15778_),
    .C(_19569_),
    .X(_16163_));
 sky130_fd_sc_hd__or2_2 _38218_ (.A(_16162_),
    .B(_16163_),
    .X(_16164_));
 sky130_fd_sc_hd__a21oi_2 _38219_ (.A1(_16156_),
    .A2(_16159_),
    .B1(_16164_),
    .Y(_16165_));
 sky130_fd_sc_hd__o211a_2 _38220_ (.A1(_16162_),
    .A2(_16163_),
    .B1(_16159_),
    .C1(_16156_),
    .X(_16166_));
 sky130_fd_sc_hd__a21boi_2 _38221_ (.A1(_15976_),
    .A2(_15986_),
    .B1_N(_15980_),
    .Y(_16167_));
 sky130_fd_sc_hd__o21ai_2 _38222_ (.A1(_16165_),
    .A2(_16166_),
    .B1(_16167_),
    .Y(_16168_));
 sky130_fd_sc_hd__nand2_2 _38223_ (.A(_15988_),
    .B(_15980_),
    .Y(_16169_));
 sky130_fd_sc_hd__a21o_2 _38224_ (.A1(_16156_),
    .A2(_16159_),
    .B1(_16164_),
    .X(_16170_));
 sky130_fd_sc_hd__nand3_2 _38225_ (.A(_16164_),
    .B(_16156_),
    .C(_16159_),
    .Y(_16171_));
 sky130_fd_sc_hd__nand3_2 _38226_ (.A(_16169_),
    .B(_16170_),
    .C(_16171_),
    .Y(_16172_));
 sky130_fd_sc_hd__o21bai_2 _38227_ (.A1(_15981_),
    .A2(_15982_),
    .B1_N(_15983_),
    .Y(_16173_));
 sky130_fd_sc_hd__nand2_2 _38228_ (.A(_19334_),
    .B(_19559_),
    .Y(_16174_));
 sky130_fd_sc_hd__nand2_2 _38229_ (.A(_11205_),
    .B(_10380_),
    .Y(_16175_));
 sky130_fd_sc_hd__nand2_2 _38230_ (.A(_10867_),
    .B(_09220_),
    .Y(_16176_));
 sky130_fd_sc_hd__nor2_2 _38231_ (.A(_16175_),
    .B(_16176_),
    .Y(_16177_));
 sky130_fd_sc_hd__nand2_2 _38232_ (.A(_16175_),
    .B(_16176_),
    .Y(_16178_));
 sky130_fd_sc_hd__or3b_2 _38233_ (.A(_16174_),
    .B(_16177_),
    .C_N(_16178_),
    .X(_16179_));
 sky130_fd_sc_hd__inv_2 _38234_ (.A(_16177_),
    .Y(_16180_));
 sky130_fd_sc_hd__nand2_2 _38235_ (.A(_16180_),
    .B(_16178_),
    .Y(_16181_));
 sky130_fd_sc_hd__nand2_2 _38236_ (.A(_16181_),
    .B(_16174_),
    .Y(_16182_));
 sky130_fd_sc_hd__nand3_2 _38237_ (.A(_16173_),
    .B(_16179_),
    .C(_16182_),
    .Y(_16183_));
 sky130_fd_sc_hd__nand2_2 _38238_ (.A(_16002_),
    .B(_15998_),
    .Y(_16184_));
 sky130_fd_sc_hd__inv_2 _38239_ (.A(_16184_),
    .Y(_16185_));
 sky130_fd_sc_hd__a21oi_2 _38240_ (.A1(_16179_),
    .A2(_16182_),
    .B1(_16173_),
    .Y(_16186_));
 sky130_fd_sc_hd__nor2_2 _38241_ (.A(_16185_),
    .B(_16186_),
    .Y(_16187_));
 sky130_fd_sc_hd__a21o_2 _38242_ (.A1(_16179_),
    .A2(_16182_),
    .B1(_16173_),
    .X(_16188_));
 sky130_fd_sc_hd__a21oi_2 _38243_ (.A1(_16188_),
    .A2(_16183_),
    .B1(_16184_),
    .Y(_16189_));
 sky130_fd_sc_hd__a21oi_2 _38244_ (.A1(_16183_),
    .A2(_16187_),
    .B1(_16189_),
    .Y(_16190_));
 sky130_fd_sc_hd__a21o_2 _38245_ (.A1(_16168_),
    .A2(_16172_),
    .B1(_16190_),
    .X(_16191_));
 sky130_fd_sc_hd__nand3_2 _38246_ (.A(_16168_),
    .B(_16172_),
    .C(_16190_),
    .Y(_16192_));
 sky130_fd_sc_hd__nor2_2 _38247_ (.A(_16022_),
    .B(_16021_),
    .Y(_16193_));
 sky130_fd_sc_hd__a21oi_2 _38248_ (.A1(_15987_),
    .A2(_15988_),
    .B1(_15968_),
    .Y(_16194_));
 sky130_fd_sc_hd__o21ai_2 _38249_ (.A1(_16193_),
    .A2(_16194_),
    .B1(_15989_),
    .Y(_16195_));
 sky130_fd_sc_hd__a21oi_2 _38250_ (.A1(_16191_),
    .A2(_16192_),
    .B1(_16195_),
    .Y(_16196_));
 sky130_fd_sc_hd__inv_2 _38251_ (.A(_15989_),
    .Y(_16197_));
 sky130_fd_sc_hd__nand2_2 _38252_ (.A(_15987_),
    .B(_15988_),
    .Y(_16198_));
 sky130_fd_sc_hd__a21oi_2 _38253_ (.A1(_15992_),
    .A2(_16198_),
    .B1(_16193_),
    .Y(_16199_));
 sky130_fd_sc_hd__o211a_2 _38254_ (.A1(_16197_),
    .A2(_16199_),
    .B1(_16192_),
    .C1(_16191_),
    .X(_16200_));
 sky130_fd_sc_hd__nand2_2 _38255_ (.A(_15947_),
    .B(_15943_),
    .Y(_16201_));
 sky130_fd_sc_hd__nand2_2 _38256_ (.A(_08382_),
    .B(_11410_),
    .Y(_16202_));
 sky130_fd_sc_hd__nand2_2 _38257_ (.A(_09617_),
    .B(_10538_),
    .Y(_16203_));
 sky130_fd_sc_hd__or2_2 _38258_ (.A(_16202_),
    .B(_16203_),
    .X(_16204_));
 sky130_fd_sc_hd__nand2_2 _38259_ (.A(_16202_),
    .B(_16203_),
    .Y(_16205_));
 sky130_fd_sc_hd__a22oi_2 _38260_ (.A1(_19344_),
    .A2(_19546_),
    .B1(_16204_),
    .B2(_16205_),
    .Y(_16206_));
 sky130_fd_sc_hd__and4_2 _38261_ (.A(_16204_),
    .B(_19343_),
    .C(_19546_),
    .D(_16205_),
    .X(_16207_));
 sky130_fd_sc_hd__nor2_2 _38262_ (.A(_16206_),
    .B(_16207_),
    .Y(_16208_));
 sky130_fd_sc_hd__nor2_2 _38263_ (.A(_16201_),
    .B(_16208_),
    .Y(_16209_));
 sky130_fd_sc_hd__and2_2 _38264_ (.A(_16208_),
    .B(_16201_),
    .X(_16210_));
 sky130_fd_sc_hd__and4_2 _38265_ (.A(_11429_),
    .B(_07481_),
    .C(_07907_),
    .D(_11427_),
    .X(_16211_));
 sky130_fd_sc_hd__nand2_2 _38266_ (.A(_11759_),
    .B(_07906_),
    .Y(_16212_));
 sky130_fd_sc_hd__o21a_2 _38267_ (.A1(_12596_),
    .A2(_10519_),
    .B1(_16212_),
    .X(_16213_));
 sky130_fd_sc_hd__nor2_2 _38268_ (.A(_16211_),
    .B(_16213_),
    .Y(_16214_));
 sky130_fd_sc_hd__xor2_2 _38269_ (.A(_15952_),
    .B(_16214_),
    .X(_16215_));
 sky130_fd_sc_hd__o21bai_2 _38270_ (.A1(_16209_),
    .A2(_16210_),
    .B1_N(_16215_),
    .Y(_16216_));
 sky130_fd_sc_hd__nand2_2 _38271_ (.A(_16208_),
    .B(_16201_),
    .Y(_16217_));
 sky130_fd_sc_hd__nand3b_2 _38272_ (.A_N(_16209_),
    .B(_16215_),
    .C(_16217_),
    .Y(_16218_));
 sky130_fd_sc_hd__a21oi_2 _38273_ (.A1(_16001_),
    .A2(_16002_),
    .B1(_16004_),
    .Y(_16219_));
 sky130_fd_sc_hd__o21ai_2 _38274_ (.A1(_16219_),
    .A2(_15995_),
    .B1(_16006_),
    .Y(_16220_));
 sky130_fd_sc_hd__a21oi_2 _38275_ (.A1(_16216_),
    .A2(_16218_),
    .B1(_16220_),
    .Y(_16221_));
 sky130_fd_sc_hd__nand3_2 _38276_ (.A(_16216_),
    .B(_16218_),
    .C(_16220_),
    .Y(_16222_));
 sky130_fd_sc_hd__nand2_2 _38277_ (.A(_15962_),
    .B(_15950_),
    .Y(_16223_));
 sky130_fd_sc_hd__nand2_2 _38278_ (.A(_16222_),
    .B(_16223_),
    .Y(_16224_));
 sky130_fd_sc_hd__nor2_2 _38279_ (.A(_16221_),
    .B(_16224_),
    .Y(_16225_));
 sky130_fd_sc_hd__nand2_2 _38280_ (.A(_16216_),
    .B(_16218_),
    .Y(_16226_));
 sky130_fd_sc_hd__inv_2 _38281_ (.A(_16220_),
    .Y(_16227_));
 sky130_fd_sc_hd__nand2_2 _38282_ (.A(_16226_),
    .B(_16227_),
    .Y(_16228_));
 sky130_fd_sc_hd__a21oi_2 _38283_ (.A1(_16228_),
    .A2(_16222_),
    .B1(_16223_),
    .Y(_16229_));
 sky130_fd_sc_hd__nor2_2 _38284_ (.A(_16225_),
    .B(_16229_),
    .Y(_16230_));
 sky130_fd_sc_hd__o21ai_2 _38285_ (.A1(_16196_),
    .A2(_16200_),
    .B1(_16230_),
    .Y(_16231_));
 sky130_fd_sc_hd__a21oi_2 _38286_ (.A1(_16024_),
    .A2(_16025_),
    .B1(_16018_),
    .Y(_16232_));
 sky130_fd_sc_hd__nand2_2 _38287_ (.A(_16191_),
    .B(_16192_),
    .Y(_16233_));
 sky130_fd_sc_hd__nor2_2 _38288_ (.A(_16197_),
    .B(_16199_),
    .Y(_16234_));
 sky130_fd_sc_hd__nand2_2 _38289_ (.A(_16233_),
    .B(_16234_),
    .Y(_16235_));
 sky130_fd_sc_hd__inv_2 _38290_ (.A(_16222_),
    .Y(_16236_));
 sky130_fd_sc_hd__inv_2 _38291_ (.A(_16223_),
    .Y(_16237_));
 sky130_fd_sc_hd__o21ai_2 _38292_ (.A1(_16221_),
    .A2(_16236_),
    .B1(_16237_),
    .Y(_16238_));
 sky130_fd_sc_hd__nand3_2 _38293_ (.A(_16228_),
    .B(_16223_),
    .C(_16222_),
    .Y(_16239_));
 sky130_fd_sc_hd__nand2_2 _38294_ (.A(_16238_),
    .B(_16239_),
    .Y(_16240_));
 sky130_fd_sc_hd__nand3_2 _38295_ (.A(_16195_),
    .B(_16191_),
    .C(_16192_),
    .Y(_16241_));
 sky130_fd_sc_hd__nand3_2 _38296_ (.A(_16235_),
    .B(_16240_),
    .C(_16241_),
    .Y(_16242_));
 sky130_fd_sc_hd__nand3_2 _38297_ (.A(_16231_),
    .B(_16232_),
    .C(_16242_),
    .Y(_16243_));
 sky130_fd_sc_hd__o22ai_2 _38298_ (.A1(_16229_),
    .A2(_16225_),
    .B1(_16196_),
    .B2(_16200_),
    .Y(_16244_));
 sky130_fd_sc_hd__a21o_2 _38299_ (.A1(_15960_),
    .A2(_15963_),
    .B1(_15965_),
    .X(_16245_));
 sky130_fd_sc_hd__nand3_2 _38300_ (.A(_15960_),
    .B(_15963_),
    .C(_15965_),
    .Y(_16246_));
 sky130_fd_sc_hd__nand2_2 _38301_ (.A(_16245_),
    .B(_16246_),
    .Y(_16247_));
 sky130_fd_sc_hd__o21ai_2 _38302_ (.A1(_16247_),
    .A2(_16016_),
    .B1(_16026_),
    .Y(_16248_));
 sky130_fd_sc_hd__nand3_2 _38303_ (.A(_16235_),
    .B(_16230_),
    .C(_16241_),
    .Y(_16249_));
 sky130_fd_sc_hd__nand3_2 _38304_ (.A(_16244_),
    .B(_16248_),
    .C(_16249_),
    .Y(_16250_));
 sky130_fd_sc_hd__nand2_2 _38305_ (.A(_16243_),
    .B(_16250_),
    .Y(_16251_));
 sky130_fd_sc_hd__inv_2 _38306_ (.A(_15965_),
    .Y(_16252_));
 sky130_fd_sc_hd__a21oi_2 _38307_ (.A1(_15961_),
    .A2(_15962_),
    .B1(_15959_),
    .Y(_16253_));
 sky130_fd_sc_hd__o21ai_2 _38308_ (.A1(_16252_),
    .A2(_16253_),
    .B1(_15963_),
    .Y(_16254_));
 sky130_fd_sc_hd__nand2_2 _38309_ (.A(_16039_),
    .B(_16045_),
    .Y(_16255_));
 sky130_fd_sc_hd__a221o_2 _38310_ (.A1(_15864_),
    .A2(_15866_),
    .B1(_15955_),
    .B2(_15952_),
    .C1(_15953_),
    .X(_16256_));
 sky130_fd_sc_hd__a21o_2 _38311_ (.A1(_15955_),
    .A2(_15952_),
    .B1(_15953_),
    .X(_16257_));
 sky130_fd_sc_hd__nand2_2 _38312_ (.A(_16257_),
    .B(_15869_),
    .Y(_16258_));
 sky130_fd_sc_hd__nand2_2 _38313_ (.A(_16256_),
    .B(_16258_),
    .Y(_16259_));
 sky130_fd_sc_hd__nand2_2 _38314_ (.A(_16259_),
    .B(_16045_),
    .Y(_16260_));
 sky130_fd_sc_hd__buf_1 _38315_ (.A(_16258_),
    .X(_16261_));
 sky130_fd_sc_hd__nand3_2 _38316_ (.A(_16256_),
    .B(_16261_),
    .C(_16038_),
    .Y(_16262_));
 sky130_fd_sc_hd__a22oi_2 _38317_ (.A1(_16041_),
    .A2(_16255_),
    .B1(_16260_),
    .B2(_16262_),
    .Y(_16263_));
 sky130_fd_sc_hd__nand3_2 _38318_ (.A(_16262_),
    .B(_16041_),
    .C(_16255_),
    .Y(_16264_));
 sky130_fd_sc_hd__a21o_2 _38319_ (.A1(_16045_),
    .A2(_16259_),
    .B1(_16264_),
    .X(_16265_));
 sky130_fd_sc_hd__nand3b_2 _38320_ (.A_N(_16263_),
    .B(_15478_),
    .C(_16265_),
    .Y(_16266_));
 sky130_fd_sc_hd__a21oi_2 _38321_ (.A1(_16045_),
    .A2(_16259_),
    .B1(_16264_),
    .Y(_16267_));
 sky130_fd_sc_hd__o21ai_2 _38322_ (.A1(_16263_),
    .A2(_16267_),
    .B1(_15886_),
    .Y(_16268_));
 sky130_fd_sc_hd__nand3_2 _38323_ (.A(_16254_),
    .B(_16266_),
    .C(_16268_),
    .Y(_16269_));
 sky130_fd_sc_hd__a21boi_2 _38324_ (.A1(_15960_),
    .A2(_15965_),
    .B1_N(_15963_),
    .Y(_16270_));
 sky130_fd_sc_hd__o21ai_2 _38325_ (.A1(_16263_),
    .A2(_16267_),
    .B1(_15478_),
    .Y(_16271_));
 sky130_fd_sc_hd__nand3b_2 _38326_ (.A_N(_16263_),
    .B(_15886_),
    .C(_16265_),
    .Y(_16272_));
 sky130_fd_sc_hd__a21boi_2 _38327_ (.A1(_16044_),
    .A2(_15476_),
    .B1_N(_16048_),
    .Y(_16273_));
 sky130_fd_sc_hd__a31oi_2 _38328_ (.A1(_16270_),
    .A2(_16271_),
    .A3(_16272_),
    .B1(_16273_),
    .Y(_16274_));
 sky130_fd_sc_hd__nand3_2 _38329_ (.A(_16270_),
    .B(_16272_),
    .C(_16271_),
    .Y(_16275_));
 sky130_fd_sc_hd__a21bo_2 _38330_ (.A1(_16044_),
    .A2(_15476_),
    .B1_N(_16048_),
    .X(_16276_));
 sky130_fd_sc_hd__a21oi_2 _38331_ (.A1(_16275_),
    .A2(_16269_),
    .B1(_16276_),
    .Y(_16277_));
 sky130_fd_sc_hd__a21oi_2 _38332_ (.A1(_16269_),
    .A2(_16274_),
    .B1(_16277_),
    .Y(_16278_));
 sky130_fd_sc_hd__nand2_2 _38333_ (.A(_16251_),
    .B(_16278_),
    .Y(_16279_));
 sky130_fd_sc_hd__nand2_2 _38334_ (.A(_16275_),
    .B(_16269_),
    .Y(_16280_));
 sky130_fd_sc_hd__nand2_2 _38335_ (.A(_16280_),
    .B(_16273_),
    .Y(_16281_));
 sky130_fd_sc_hd__nand3_2 _38336_ (.A(_16275_),
    .B(_16269_),
    .C(_16276_),
    .Y(_16282_));
 sky130_fd_sc_hd__nand2_2 _38337_ (.A(_16281_),
    .B(_16282_),
    .Y(_16283_));
 sky130_fd_sc_hd__nand3_2 _38338_ (.A(_16243_),
    .B(_16250_),
    .C(_16283_),
    .Y(_16284_));
 sky130_fd_sc_hd__nand3_2 _38339_ (.A(_16148_),
    .B(_16279_),
    .C(_16284_),
    .Y(_16285_));
 sky130_fd_sc_hd__a21oi_2 _38340_ (.A1(_16070_),
    .A2(_16061_),
    .B1(_16083_),
    .Y(_16286_));
 sky130_fd_sc_hd__and2_2 _38341_ (.A(_15752_),
    .B(_13406_),
    .X(_16287_));
 sky130_fd_sc_hd__o21a_2 _38342_ (.A1(_15753_),
    .A2(_16287_),
    .B1(_16061_),
    .X(_16288_));
 sky130_fd_sc_hd__o2bb2ai_2 _38343_ (.A1_N(_16070_),
    .A2_N(_16288_),
    .B1(_16087_),
    .B2(_15753_),
    .Y(_16289_));
 sky130_fd_sc_hd__nor2_2 _38344_ (.A(_16286_),
    .B(_16289_),
    .Y(_16290_));
 sky130_fd_sc_hd__a21o_2 _38345_ (.A1(_16070_),
    .A2(_16061_),
    .B1(_16085_),
    .X(_16291_));
 sky130_fd_sc_hd__nand2_2 _38346_ (.A(_16288_),
    .B(_16070_),
    .Y(_16292_));
 sky130_fd_sc_hd__buf_1 _38347_ (.A(_16092_),
    .X(_16293_));
 sky130_fd_sc_hd__buf_1 _38348_ (.A(_16293_),
    .X(_16294_));
 sky130_fd_sc_hd__a21oi_2 _38349_ (.A1(_16291_),
    .A2(_16292_),
    .B1(_16294_),
    .Y(_16295_));
 sky130_fd_sc_hd__nor2_2 _38350_ (.A(_16290_),
    .B(_16295_),
    .Y(_16296_));
 sky130_fd_sc_hd__o21ai_2 _38351_ (.A1(_16071_),
    .A2(_16030_),
    .B1(_16072_),
    .Y(_16297_));
 sky130_fd_sc_hd__inv_2 _38352_ (.A(_16282_),
    .Y(_16298_));
 sky130_fd_sc_hd__o2bb2ai_2 _38353_ (.A1_N(_16250_),
    .A2_N(_16243_),
    .B1(_16277_),
    .B2(_16298_),
    .Y(_16299_));
 sky130_fd_sc_hd__nand3_2 _38354_ (.A(_16243_),
    .B(_16250_),
    .C(_16278_),
    .Y(_16300_));
 sky130_fd_sc_hd__nand3_2 _38355_ (.A(_16297_),
    .B(_16299_),
    .C(_16300_),
    .Y(_16301_));
 sky130_fd_sc_hd__nand3_2 _38356_ (.A(_16285_),
    .B(_16296_),
    .C(_16301_),
    .Y(_16302_));
 sky130_fd_sc_hd__o2bb2ai_2 _38357_ (.A1_N(_16301_),
    .A2_N(_16285_),
    .B1(_16295_),
    .B2(_16290_),
    .Y(_16303_));
 sky130_fd_sc_hd__o211ai_2 _38358_ (.A1(_16147_),
    .A2(_16098_),
    .B1(_16302_),
    .C1(_16303_),
    .Y(_16304_));
 sky130_fd_sc_hd__a21o_2 _38359_ (.A1(_16291_),
    .A2(_16292_),
    .B1(_16093_),
    .X(_16305_));
 sky130_fd_sc_hd__o21ai_2 _38360_ (.A1(_16286_),
    .A2(_16289_),
    .B1(_16305_),
    .Y(_16306_));
 sky130_fd_sc_hd__a21o_2 _38361_ (.A1(_16285_),
    .A2(_16301_),
    .B1(_16306_),
    .X(_16307_));
 sky130_fd_sc_hd__a21boi_2 _38362_ (.A1(_16074_),
    .A2(_16102_),
    .B1_N(_16080_),
    .Y(_16308_));
 sky130_fd_sc_hd__nand3_2 _38363_ (.A(_16306_),
    .B(_16285_),
    .C(_16301_),
    .Y(_16309_));
 sky130_fd_sc_hd__nand3_2 _38364_ (.A(_16307_),
    .B(_16308_),
    .C(_16309_),
    .Y(_16310_));
 sky130_fd_sc_hd__nand2_2 _38365_ (.A(_16094_),
    .B(_16293_),
    .Y(_16311_));
 sky130_fd_sc_hd__nand2_2 _38366_ (.A(_16311_),
    .B(_16091_),
    .Y(_16312_));
 sky130_fd_sc_hd__inv_2 _38367_ (.A(_16312_),
    .Y(_16313_));
 sky130_fd_sc_hd__nor2_2 _38368_ (.A(_15081_),
    .B(_16313_),
    .Y(_16314_));
 sky130_fd_sc_hd__nor2_2 _38369_ (.A(_14823_),
    .B(_16312_),
    .Y(_16315_));
 sky130_fd_sc_hd__o2bb2ai_2 _38370_ (.A1_N(_16304_),
    .A2_N(_16310_),
    .B1(_16314_),
    .B2(_16315_),
    .Y(_16316_));
 sky130_fd_sc_hd__nor2_2 _38371_ (.A(_16315_),
    .B(_16314_),
    .Y(_16317_));
 sky130_fd_sc_hd__nand3_2 _38372_ (.A(_16310_),
    .B(_16304_),
    .C(_16317_),
    .Y(_16318_));
 sky130_fd_sc_hd__nand3_2 _38373_ (.A(_16146_),
    .B(_16316_),
    .C(_16318_),
    .Y(_16319_));
 sky130_fd_sc_hd__inv_2 _38374_ (.A(_16317_),
    .Y(_16320_));
 sky130_fd_sc_hd__nand3_2 _38375_ (.A(_16310_),
    .B(_16304_),
    .C(_16320_),
    .Y(_16321_));
 sky130_fd_sc_hd__nor2_2 _38376_ (.A(_16118_),
    .B(_16313_),
    .Y(_16322_));
 sky130_fd_sc_hd__nor2_2 _38377_ (.A(_16120_),
    .B(_16312_),
    .Y(_16323_));
 sky130_fd_sc_hd__o2bb2ai_2 _38378_ (.A1_N(_16304_),
    .A2_N(_16310_),
    .B1(_16322_),
    .B2(_16323_),
    .Y(_16324_));
 sky130_fd_sc_hd__o211ai_2 _38379_ (.A1(_16145_),
    .A2(_16123_),
    .B1(_16321_),
    .C1(_16324_),
    .Y(_16325_));
 sky130_fd_sc_hd__nand2_2 _38380_ (.A(_16319_),
    .B(_16325_),
    .Y(_16326_));
 sky130_fd_sc_hd__nand2_2 _38381_ (.A(_16326_),
    .B(_16119_),
    .Y(_16327_));
 sky130_fd_sc_hd__a21oi_2 _38382_ (.A1(_16115_),
    .A2(_16114_),
    .B1(_15939_),
    .Y(_16328_));
 sky130_fd_sc_hd__a21oi_2 _38383_ (.A1(_16116_),
    .A2(_15913_),
    .B1(_16328_),
    .Y(_16329_));
 sky130_fd_sc_hd__inv_2 _38384_ (.A(_16119_),
    .Y(_16330_));
 sky130_fd_sc_hd__nand3_2 _38385_ (.A(_16319_),
    .B(_16325_),
    .C(_16330_),
    .Y(_16331_));
 sky130_fd_sc_hd__nand3_2 _38386_ (.A(_16327_),
    .B(_16329_),
    .C(_16331_),
    .Y(_16332_));
 sky130_fd_sc_hd__a31oi_2 _38387_ (.A1(_15939_),
    .A2(_16115_),
    .A3(_16114_),
    .B1(_16129_),
    .Y(_16333_));
 sky130_fd_sc_hd__nand3_2 _38388_ (.A(_16319_),
    .B(_16325_),
    .C(_16119_),
    .Y(_16334_));
 sky130_fd_sc_hd__o2bb2ai_2 _38389_ (.A1_N(_16325_),
    .A2_N(_16319_),
    .B1(_15729_),
    .B2(_16111_),
    .Y(_16335_));
 sky130_fd_sc_hd__o211ai_2 _38390_ (.A1(_16328_),
    .A2(_16333_),
    .B1(_16334_),
    .C1(_16335_),
    .Y(_16336_));
 sky130_fd_sc_hd__nand2_2 _38391_ (.A(_16332_),
    .B(_16336_),
    .Y(_16337_));
 sky130_fd_sc_hd__a21oi_2 _38392_ (.A1(_16143_),
    .A2(_16137_),
    .B1(_16337_),
    .Y(_16338_));
 sky130_fd_sc_hd__and3_2 _38393_ (.A(_16143_),
    .B(_16137_),
    .C(_16337_),
    .X(_16339_));
 sky130_fd_sc_hd__nor2_2 _38394_ (.A(_16338_),
    .B(_16339_),
    .Y(_02670_));
 sky130_fd_sc_hd__inv_2 _38395_ (.A(_16321_),
    .Y(_16340_));
 sky130_fd_sc_hd__o21ai_2 _38396_ (.A1(_16145_),
    .A2(_16123_),
    .B1(_16324_),
    .Y(_16341_));
 sky130_fd_sc_hd__o2bb2ai_2 _38397_ (.A1_N(_16119_),
    .A2_N(_16319_),
    .B1(_16340_),
    .B2(_16341_),
    .Y(_16342_));
 sky130_fd_sc_hd__o21ai_2 _38398_ (.A1(_16240_),
    .A2(_16196_),
    .B1(_16241_),
    .Y(_16343_));
 sky130_fd_sc_hd__nand2_2 _38399_ (.A(_16171_),
    .B(_16156_),
    .Y(_16344_));
 sky130_fd_sc_hd__o21bai_2 _38400_ (.A1(_16150_),
    .A2(_16152_),
    .B1_N(_16151_),
    .Y(_16345_));
 sky130_fd_sc_hd__nand2_2 _38401_ (.A(_10827_),
    .B(_08910_),
    .Y(_16346_));
 sky130_fd_sc_hd__and4_2 _38402_ (.A(_09256_),
    .B(_11169_),
    .C(_13146_),
    .D(_07849_),
    .X(_16347_));
 sky130_fd_sc_hd__o22a_2 _38403_ (.A1(_08650_),
    .A2(_11509_),
    .B1(_10832_),
    .B2(_09678_),
    .X(_16348_));
 sky130_fd_sc_hd__nor2_2 _38404_ (.A(_16347_),
    .B(_16348_),
    .Y(_16349_));
 sky130_fd_sc_hd__or2_2 _38405_ (.A(_16346_),
    .B(_16349_),
    .X(_16350_));
 sky130_fd_sc_hd__nand2_2 _38406_ (.A(_16349_),
    .B(_16346_),
    .Y(_16351_));
 sky130_fd_sc_hd__nand3b_2 _38407_ (.A_N(_16345_),
    .B(_16350_),
    .C(_16351_),
    .Y(_16352_));
 sky130_fd_sc_hd__nor2_2 _38408_ (.A(_16346_),
    .B(_16349_),
    .Y(_16353_));
 sky130_fd_sc_hd__and2_2 _38409_ (.A(_16349_),
    .B(_16346_),
    .X(_16354_));
 sky130_fd_sc_hd__o21ai_2 _38410_ (.A1(_16353_),
    .A2(_16354_),
    .B1(_16345_),
    .Y(_16355_));
 sky130_fd_sc_hd__nand2_2 _38411_ (.A(_15778_),
    .B(_19566_),
    .Y(_16356_));
 sky130_fd_sc_hd__o22a_2 _38412_ (.A1(_14371_),
    .A2(_12089_),
    .B1(_14869_),
    .B2(_10485_),
    .X(_16357_));
 sky130_fd_sc_hd__and3_2 _38413_ (.A(_15781_),
    .B(_09223_),
    .C(_10966_),
    .X(_16358_));
 sky130_fd_sc_hd__nor3_2 _38414_ (.A(_16356_),
    .B(_16357_),
    .C(_16358_),
    .Y(_16359_));
 sky130_fd_sc_hd__o21a_2 _38415_ (.A1(_16357_),
    .A2(_16358_),
    .B1(_16356_),
    .X(_16360_));
 sky130_fd_sc_hd__nor2_2 _38416_ (.A(_16359_),
    .B(_16360_),
    .Y(_16361_));
 sky130_fd_sc_hd__a21o_2 _38417_ (.A1(_16352_),
    .A2(_16355_),
    .B1(_16361_),
    .X(_16362_));
 sky130_fd_sc_hd__nand3_2 _38418_ (.A(_16352_),
    .B(_16355_),
    .C(_16361_),
    .Y(_16363_));
 sky130_fd_sc_hd__nand3_2 _38419_ (.A(_16344_),
    .B(_16362_),
    .C(_16363_),
    .Y(_16364_));
 sky130_fd_sc_hd__a21oi_2 _38420_ (.A1(_16352_),
    .A2(_16355_),
    .B1(_16361_),
    .Y(_16365_));
 sky130_fd_sc_hd__and3_2 _38421_ (.A(_16352_),
    .B(_16355_),
    .C(_16361_),
    .X(_16366_));
 sky130_fd_sc_hd__a21boi_2 _38422_ (.A1(_16159_),
    .A2(_16164_),
    .B1_N(_16156_),
    .Y(_16367_));
 sky130_fd_sc_hd__o21ai_2 _38423_ (.A1(_16365_),
    .A2(_16366_),
    .B1(_16367_),
    .Y(_16368_));
 sky130_fd_sc_hd__nand2_2 _38424_ (.A(_19335_),
    .B(_19554_),
    .Y(_16369_));
 sky130_fd_sc_hd__and4_2 _38425_ (.A(_19329_),
    .B(_14068_),
    .C(_09733_),
    .D(_09216_),
    .X(_16370_));
 sky130_fd_sc_hd__nand2_2 _38426_ (.A(_19329_),
    .B(_09216_),
    .Y(_16371_));
 sky130_fd_sc_hd__o21a_2 _38427_ (.A1(_13873_),
    .A2(_13274_),
    .B1(_16371_),
    .X(_16372_));
 sky130_fd_sc_hd__or3_2 _38428_ (.A(_16369_),
    .B(_16370_),
    .C(_16372_),
    .X(_16373_));
 sky130_fd_sc_hd__o21ai_2 _38429_ (.A1(_16370_),
    .A2(_16372_),
    .B1(_16369_),
    .Y(_16374_));
 sky130_fd_sc_hd__and3_2 _38430_ (.A(_15781_),
    .B(_19572_),
    .C(_19575_),
    .X(_16375_));
 sky130_fd_sc_hd__a31o_2 _38431_ (.A1(_15778_),
    .A2(_19569_),
    .A3(_16160_),
    .B1(_16375_),
    .X(_16376_));
 sky130_fd_sc_hd__a21o_2 _38432_ (.A1(_16373_),
    .A2(_16374_),
    .B1(_16376_),
    .X(_16377_));
 sky130_fd_sc_hd__nand2_2 _38433_ (.A(_16179_),
    .B(_16180_),
    .Y(_16378_));
 sky130_fd_sc_hd__nand3_2 _38434_ (.A(_16373_),
    .B(_16376_),
    .C(_16374_),
    .Y(_16379_));
 sky130_fd_sc_hd__nand3_2 _38435_ (.A(_16377_),
    .B(_16378_),
    .C(_16379_),
    .Y(_16380_));
 sky130_fd_sc_hd__inv_2 _38436_ (.A(_16380_),
    .Y(_16381_));
 sky130_fd_sc_hd__nand2_2 _38437_ (.A(_16377_),
    .B(_16379_),
    .Y(_16382_));
 sky130_fd_sc_hd__inv_2 _38438_ (.A(_16378_),
    .Y(_16383_));
 sky130_fd_sc_hd__nand2_2 _38439_ (.A(_16382_),
    .B(_16383_),
    .Y(_16384_));
 sky130_fd_sc_hd__inv_2 _38440_ (.A(_16384_),
    .Y(_16385_));
 sky130_fd_sc_hd__o2bb2ai_2 _38441_ (.A1_N(_16364_),
    .A2_N(_16368_),
    .B1(_16381_),
    .B2(_16385_),
    .Y(_16386_));
 sky130_fd_sc_hd__nand2_2 _38442_ (.A(_16192_),
    .B(_16172_),
    .Y(_16387_));
 sky130_fd_sc_hd__nand2_2 _38443_ (.A(_16384_),
    .B(_16380_),
    .Y(_16388_));
 sky130_fd_sc_hd__nand3b_2 _38444_ (.A_N(_16388_),
    .B(_16368_),
    .C(_16364_),
    .Y(_16389_));
 sky130_fd_sc_hd__nand3_2 _38445_ (.A(_16386_),
    .B(_16387_),
    .C(_16389_),
    .Y(_16390_));
 sky130_fd_sc_hd__nor2_2 _38446_ (.A(_16378_),
    .B(_16382_),
    .Y(_16391_));
 sky130_fd_sc_hd__inv_2 _38447_ (.A(_16382_),
    .Y(_16392_));
 sky130_fd_sc_hd__nor2_2 _38448_ (.A(_16383_),
    .B(_16392_),
    .Y(_16393_));
 sky130_fd_sc_hd__o2bb2ai_2 _38449_ (.A1_N(_16364_),
    .A2_N(_16368_),
    .B1(_16391_),
    .B2(_16393_),
    .Y(_16394_));
 sky130_fd_sc_hd__a21boi_2 _38450_ (.A1(_16168_),
    .A2(_16190_),
    .B1_N(_16172_),
    .Y(_16395_));
 sky130_fd_sc_hd__nand3_2 _38451_ (.A(_16368_),
    .B(_16364_),
    .C(_16388_),
    .Y(_16396_));
 sky130_fd_sc_hd__nand3_2 _38452_ (.A(_16394_),
    .B(_16395_),
    .C(_16396_),
    .Y(_16397_));
 sky130_fd_sc_hd__nand2_2 _38453_ (.A(_16390_),
    .B(_16397_),
    .Y(_16398_));
 sky130_fd_sc_hd__o21ai_2 _38454_ (.A1(_16185_),
    .A2(_16186_),
    .B1(_16183_),
    .Y(_16399_));
 sky130_fd_sc_hd__inv_2 _38455_ (.A(_16204_),
    .Y(_16400_));
 sky130_fd_sc_hd__nand2_2 _38456_ (.A(_08790_),
    .B(_10538_),
    .Y(_16401_));
 sky130_fd_sc_hd__nand2_2 _38457_ (.A(_09617_),
    .B(_11037_),
    .Y(_16402_));
 sky130_fd_sc_hd__or2_2 _38458_ (.A(_16401_),
    .B(_16402_),
    .X(_16403_));
 sky130_fd_sc_hd__nand2_2 _38459_ (.A(_16401_),
    .B(_16402_),
    .Y(_16404_));
 sky130_fd_sc_hd__nand2_2 _38460_ (.A(_19343_),
    .B(_19541_),
    .Y(_16405_));
 sky130_fd_sc_hd__a21bo_2 _38461_ (.A1(_16403_),
    .A2(_16404_),
    .B1_N(_16405_),
    .X(_16406_));
 sky130_fd_sc_hd__nand3b_2 _38462_ (.A_N(_16405_),
    .B(_16403_),
    .C(_16404_),
    .Y(_16407_));
 sky130_fd_sc_hd__nand2_2 _38463_ (.A(_16406_),
    .B(_16407_),
    .Y(_16408_));
 sky130_fd_sc_hd__o21bai_2 _38464_ (.A1(_16400_),
    .A2(_16207_),
    .B1_N(_16408_),
    .Y(_16409_));
 sky130_fd_sc_hd__nor2_2 _38465_ (.A(_16400_),
    .B(_16207_),
    .Y(_16410_));
 sky130_fd_sc_hd__nand2_2 _38466_ (.A(_16410_),
    .B(_16408_),
    .Y(_16411_));
 sky130_fd_sc_hd__nand2_2 _38467_ (.A(_16409_),
    .B(_16411_),
    .Y(_16412_));
 sky130_fd_sc_hd__nand2_2 _38468_ (.A(_11023_),
    .B(_07483_),
    .Y(_16413_));
 sky130_fd_sc_hd__or2_2 _38469_ (.A(_16212_),
    .B(_16413_),
    .X(_16414_));
 sky130_fd_sc_hd__nand2_2 _38470_ (.A(_16212_),
    .B(_16413_),
    .Y(_16415_));
 sky130_fd_sc_hd__nand2_2 _38471_ (.A(_16414_),
    .B(_16415_),
    .Y(_16416_));
 sky130_fd_sc_hd__nor2_2 _38472_ (.A(_15951_),
    .B(_16416_),
    .Y(_16417_));
 sky130_fd_sc_hd__nand2_2 _38473_ (.A(_16416_),
    .B(_15951_),
    .Y(_16418_));
 sky130_fd_sc_hd__and2b_2 _38474_ (.A_N(_16417_),
    .B(_16418_),
    .X(_16419_));
 sky130_fd_sc_hd__buf_1 _38475_ (.A(_16419_),
    .X(_16420_));
 sky130_fd_sc_hd__nand2_2 _38476_ (.A(_16412_),
    .B(_16420_),
    .Y(_16421_));
 sky130_fd_sc_hd__and2_2 _38477_ (.A(_16414_),
    .B(_16415_),
    .X(_16422_));
 sky130_fd_sc_hd__nand2_2 _38478_ (.A(_16422_),
    .B(_15952_),
    .Y(_16423_));
 sky130_fd_sc_hd__nand2_2 _38479_ (.A(_16423_),
    .B(_16418_),
    .Y(_16424_));
 sky130_fd_sc_hd__buf_1 _38480_ (.A(_16424_),
    .X(_16425_));
 sky130_fd_sc_hd__nand3_2 _38481_ (.A(_16409_),
    .B(_16411_),
    .C(_16425_),
    .Y(_16426_));
 sky130_fd_sc_hd__nand3b_2 _38482_ (.A_N(_16399_),
    .B(_16421_),
    .C(_16426_),
    .Y(_16427_));
 sky130_fd_sc_hd__nand2_2 _38483_ (.A(_16412_),
    .B(_16425_),
    .Y(_16428_));
 sky130_fd_sc_hd__nand3_2 _38484_ (.A(_16409_),
    .B(_16411_),
    .C(_16420_),
    .Y(_16429_));
 sky130_fd_sc_hd__a32oi_2 _38485_ (.A1(_16428_),
    .A2(_16399_),
    .A3(_16429_),
    .B1(_16217_),
    .B2(_16218_),
    .Y(_16430_));
 sky130_fd_sc_hd__nand3_2 _38486_ (.A(_16428_),
    .B(_16399_),
    .C(_16429_),
    .Y(_16431_));
 sky130_fd_sc_hd__nand2_2 _38487_ (.A(_16218_),
    .B(_16217_),
    .Y(_16432_));
 sky130_fd_sc_hd__a21oi_2 _38488_ (.A1(_16427_),
    .A2(_16431_),
    .B1(_16432_),
    .Y(_16433_));
 sky130_fd_sc_hd__a21oi_2 _38489_ (.A1(_16427_),
    .A2(_16430_),
    .B1(_16433_),
    .Y(_16434_));
 sky130_fd_sc_hd__inv_2 _38490_ (.A(_16434_),
    .Y(_16435_));
 sky130_fd_sc_hd__nand2_2 _38491_ (.A(_16398_),
    .B(_16435_),
    .Y(_16436_));
 sky130_fd_sc_hd__nand3_2 _38492_ (.A(_16390_),
    .B(_16397_),
    .C(_16434_),
    .Y(_16437_));
 sky130_fd_sc_hd__nand3_2 _38493_ (.A(_16343_),
    .B(_16436_),
    .C(_16437_),
    .Y(_16438_));
 sky130_fd_sc_hd__a21oi_2 _38494_ (.A1(_16235_),
    .A2(_16230_),
    .B1(_16200_),
    .Y(_16439_));
 sky130_fd_sc_hd__nand2_2 _38495_ (.A(_16398_),
    .B(_16434_),
    .Y(_16440_));
 sky130_fd_sc_hd__nand3_2 _38496_ (.A(_16435_),
    .B(_16397_),
    .C(_16390_),
    .Y(_16441_));
 sky130_fd_sc_hd__nand3_2 _38497_ (.A(_16439_),
    .B(_16440_),
    .C(_16441_),
    .Y(_16442_));
 sky130_fd_sc_hd__nand2_2 _38498_ (.A(_15863_),
    .B(_19360_),
    .Y(_16443_));
 sky130_fd_sc_hd__nand2_2 _38499_ (.A(_15862_),
    .B(_15451_),
    .Y(_16444_));
 sky130_fd_sc_hd__nand2_2 _38500_ (.A(_16443_),
    .B(_16444_),
    .Y(_16445_));
 sky130_fd_sc_hd__o21bai_2 _38501_ (.A1(_15951_),
    .A2(_16213_),
    .B1_N(_16211_),
    .Y(_16446_));
 sky130_fd_sc_hd__xor2_2 _38502_ (.A(_16445_),
    .B(_16446_),
    .X(_16447_));
 sky130_fd_sc_hd__a21oi_2 _38503_ (.A1(_16262_),
    .A2(_16261_),
    .B1(_16447_),
    .Y(_16448_));
 sky130_fd_sc_hd__nand2_2 _38504_ (.A(_16447_),
    .B(_16261_),
    .Y(_16449_));
 sky130_fd_sc_hd__a31o_2 _38505_ (.A1(_16038_),
    .A2(_16256_),
    .A3(_16261_),
    .B1(_16449_),
    .X(_16450_));
 sky130_fd_sc_hd__nand2_2 _38506_ (.A(_16450_),
    .B(_15475_),
    .Y(_16451_));
 sky130_fd_sc_hd__and3_2 _38507_ (.A(_16262_),
    .B(_16261_),
    .C(_16447_),
    .X(_16452_));
 sky130_fd_sc_hd__o21ai_2 _38508_ (.A1(_16448_),
    .A2(_16452_),
    .B1(_15886_),
    .Y(_16453_));
 sky130_fd_sc_hd__o21ai_2 _38509_ (.A1(_16448_),
    .A2(_16451_),
    .B1(_16453_),
    .Y(_16454_));
 sky130_fd_sc_hd__nand3_2 _38510_ (.A(_16454_),
    .B(_16222_),
    .C(_16239_),
    .Y(_16455_));
 sky130_fd_sc_hd__nor2_2 _38511_ (.A(_16237_),
    .B(_16221_),
    .Y(_16456_));
 sky130_fd_sc_hd__o21ai_2 _38512_ (.A1(_16448_),
    .A2(_16452_),
    .B1(_15475_),
    .Y(_16457_));
 sky130_fd_sc_hd__a21o_2 _38513_ (.A1(_16262_),
    .A2(_16261_),
    .B1(_16447_),
    .X(_16458_));
 sky130_fd_sc_hd__nand3_2 _38514_ (.A(_16458_),
    .B(_16450_),
    .C(_15585_),
    .Y(_16459_));
 sky130_fd_sc_hd__nand2_2 _38515_ (.A(_16457_),
    .B(_16459_),
    .Y(_16460_));
 sky130_fd_sc_hd__o21ai_2 _38516_ (.A1(_16236_),
    .A2(_16456_),
    .B1(_16460_),
    .Y(_16461_));
 sky130_fd_sc_hd__o21ai_2 _38517_ (.A1(_15586_),
    .A2(_16263_),
    .B1(_16265_),
    .Y(_16462_));
 sky130_fd_sc_hd__a21oi_2 _38518_ (.A1(_16455_),
    .A2(_16461_),
    .B1(_16462_),
    .Y(_16463_));
 sky130_fd_sc_hd__nand3_2 _38519_ (.A(_16455_),
    .B(_16461_),
    .C(_16462_),
    .Y(_16464_));
 sky130_fd_sc_hd__inv_2 _38520_ (.A(_16464_),
    .Y(_16465_));
 sky130_fd_sc_hd__o2bb2ai_2 _38521_ (.A1_N(_16438_),
    .A2_N(_16442_),
    .B1(_16463_),
    .B2(_16465_),
    .Y(_16466_));
 sky130_fd_sc_hd__o31a_2 _38522_ (.A1(_16236_),
    .A2(_16456_),
    .A3(_16460_),
    .B1(_16462_),
    .X(_16467_));
 sky130_fd_sc_hd__a21oi_2 _38523_ (.A1(_16467_),
    .A2(_16461_),
    .B1(_16463_),
    .Y(_16468_));
 sky130_fd_sc_hd__nand3_2 _38524_ (.A(_16442_),
    .B(_16438_),
    .C(_16468_),
    .Y(_16469_));
 sky130_fd_sc_hd__nand2_2 _38525_ (.A(_16243_),
    .B(_16278_),
    .Y(_16470_));
 sky130_fd_sc_hd__nand2_2 _38526_ (.A(_16470_),
    .B(_16250_),
    .Y(_16471_));
 sky130_fd_sc_hd__a21oi_2 _38527_ (.A1(_16466_),
    .A2(_16469_),
    .B1(_16471_),
    .Y(_16472_));
 sky130_fd_sc_hd__and3_2 _38528_ (.A(_16244_),
    .B(_16248_),
    .C(_16249_),
    .X(_16473_));
 sky130_fd_sc_hd__a31oi_2 _38529_ (.A1(_16231_),
    .A2(_16232_),
    .A3(_16242_),
    .B1(_16283_),
    .Y(_16474_));
 sky130_fd_sc_hd__o211a_2 _38530_ (.A1(_16473_),
    .A2(_16474_),
    .B1(_16469_),
    .C1(_16466_),
    .X(_16475_));
 sky130_fd_sc_hd__a21o_2 _38531_ (.A1(_16282_),
    .A2(_16269_),
    .B1(_16085_),
    .X(_16476_));
 sky130_fd_sc_hd__nand3_2 _38532_ (.A(_16282_),
    .B(_15756_),
    .C(_16269_),
    .Y(_16477_));
 sky130_fd_sc_hd__nand2_2 _38533_ (.A(_16477_),
    .B(_16293_),
    .Y(_16478_));
 sky130_fd_sc_hd__inv_2 _38534_ (.A(_16478_),
    .Y(_16479_));
 sky130_fd_sc_hd__a21oi_2 _38535_ (.A1(_16476_),
    .A2(_16477_),
    .B1(_16093_),
    .Y(_16480_));
 sky130_fd_sc_hd__a21o_2 _38536_ (.A1(_16476_),
    .A2(_16479_),
    .B1(_16480_),
    .X(_16481_));
 sky130_fd_sc_hd__o21ai_2 _38537_ (.A1(_16472_),
    .A2(_16475_),
    .B1(_16481_),
    .Y(_16482_));
 sky130_fd_sc_hd__a21oi_2 _38538_ (.A1(_16299_),
    .A2(_16300_),
    .B1(_16297_),
    .Y(_16483_));
 sky130_fd_sc_hd__o21ai_2 _38539_ (.A1(_16306_),
    .A2(_16483_),
    .B1(_16301_),
    .Y(_16484_));
 sky130_fd_sc_hd__nand2_2 _38540_ (.A(_16466_),
    .B(_16469_),
    .Y(_16485_));
 sky130_fd_sc_hd__nor2_2 _38541_ (.A(_16473_),
    .B(_16474_),
    .Y(_16486_));
 sky130_fd_sc_hd__nand2_2 _38542_ (.A(_16485_),
    .B(_16486_),
    .Y(_16487_));
 sky130_fd_sc_hd__a21oi_2 _38543_ (.A1(_16479_),
    .A2(_16476_),
    .B1(_16480_),
    .Y(_16488_));
 sky130_fd_sc_hd__nand3_2 _38544_ (.A(_16471_),
    .B(_16469_),
    .C(_16466_),
    .Y(_16489_));
 sky130_fd_sc_hd__nand3_2 _38545_ (.A(_16487_),
    .B(_16488_),
    .C(_16489_),
    .Y(_16490_));
 sky130_fd_sc_hd__nand3_2 _38546_ (.A(_16482_),
    .B(_16484_),
    .C(_16490_),
    .Y(_16491_));
 sky130_fd_sc_hd__o21ai_2 _38547_ (.A1(_16472_),
    .A2(_16475_),
    .B1(_16488_),
    .Y(_16492_));
 sky130_fd_sc_hd__a21boi_2 _38548_ (.A1(_16285_),
    .A2(_16296_),
    .B1_N(_16301_),
    .Y(_16493_));
 sky130_fd_sc_hd__nand3_2 _38549_ (.A(_16487_),
    .B(_16481_),
    .C(_16489_),
    .Y(_16494_));
 sky130_fd_sc_hd__nand3_2 _38550_ (.A(_16492_),
    .B(_16493_),
    .C(_16494_),
    .Y(_16495_));
 sky130_fd_sc_hd__nand2_2 _38551_ (.A(_16491_),
    .B(_16495_),
    .Y(_16496_));
 sky130_fd_sc_hd__nand2_2 _38552_ (.A(_16289_),
    .B(_16291_),
    .Y(_16497_));
 sky130_fd_sc_hd__nor2_2 _38553_ (.A(_13737_),
    .B(_16497_),
    .Y(_16498_));
 sky130_fd_sc_hd__inv_2 _38554_ (.A(_16497_),
    .Y(_16499_));
 sky130_fd_sc_hd__nor2_2 _38555_ (.A(_14017_),
    .B(_16499_),
    .Y(_16500_));
 sky130_fd_sc_hd__nor2_2 _38556_ (.A(_16498_),
    .B(_16500_),
    .Y(_16501_));
 sky130_fd_sc_hd__nand2_2 _38557_ (.A(_16496_),
    .B(_16501_),
    .Y(_16502_));
 sky130_fd_sc_hd__a21boi_2 _38558_ (.A1(_16310_),
    .A2(_16320_),
    .B1_N(_16304_),
    .Y(_16503_));
 sky130_fd_sc_hd__nand3b_2 _38559_ (.A_N(_16501_),
    .B(_16491_),
    .C(_16495_),
    .Y(_16504_));
 sky130_fd_sc_hd__nand3_2 _38560_ (.A(_16502_),
    .B(_16503_),
    .C(_16504_),
    .Y(_16505_));
 sky130_fd_sc_hd__a21oi_2 _38561_ (.A1(_16307_),
    .A2(_16309_),
    .B1(_16308_),
    .Y(_16506_));
 sky130_fd_sc_hd__a31oi_2 _38562_ (.A1(_16307_),
    .A2(_16308_),
    .A3(_16309_),
    .B1(_16317_),
    .Y(_16507_));
 sky130_fd_sc_hd__nand3_2 _38563_ (.A(_16491_),
    .B(_16495_),
    .C(_16501_),
    .Y(_16508_));
 sky130_fd_sc_hd__o2bb2ai_2 _38564_ (.A1_N(_16495_),
    .A2_N(_16491_),
    .B1(_16500_),
    .B2(_16498_),
    .Y(_16509_));
 sky130_fd_sc_hd__o211ai_2 _38565_ (.A1(_16506_),
    .A2(_16507_),
    .B1(_16508_),
    .C1(_16509_),
    .Y(_16510_));
 sky130_fd_sc_hd__inv_2 _38566_ (.A(_16322_),
    .Y(_16511_));
 sky130_fd_sc_hd__a21o_2 _38567_ (.A1(_16505_),
    .A2(_16510_),
    .B1(_16511_),
    .X(_16512_));
 sky130_fd_sc_hd__nand3_2 _38568_ (.A(_16505_),
    .B(_16510_),
    .C(_16511_),
    .Y(_16513_));
 sky130_fd_sc_hd__nand3b_2 _38569_ (.A_N(_16342_),
    .B(_16512_),
    .C(_16513_),
    .Y(_16514_));
 sky130_fd_sc_hd__o2bb2ai_2 _38570_ (.A1_N(_16505_),
    .A2_N(_16510_),
    .B1(_15729_),
    .B2(_16313_),
    .Y(_16515_));
 sky130_fd_sc_hd__nand3_2 _38571_ (.A(_16505_),
    .B(_16510_),
    .C(_16322_),
    .Y(_16516_));
 sky130_fd_sc_hd__nand3_2 _38572_ (.A(_16515_),
    .B(_16342_),
    .C(_16516_),
    .Y(_16517_));
 sky130_fd_sc_hd__and2_2 _38573_ (.A(_16514_),
    .B(_16517_),
    .X(_16518_));
 sky130_fd_sc_hd__inv_2 _38574_ (.A(_16518_),
    .Y(_16519_));
 sky130_fd_sc_hd__nor2_2 _38575_ (.A(_16337_),
    .B(_16138_),
    .Y(_16520_));
 sky130_fd_sc_hd__nand3_2 _38576_ (.A(_16520_),
    .B(_15735_),
    .C(_15933_),
    .Y(_16521_));
 sky130_fd_sc_hd__inv_2 _38577_ (.A(_16521_),
    .Y(_16522_));
 sky130_fd_sc_hd__inv_2 _38578_ (.A(_16136_),
    .Y(_16523_));
 sky130_fd_sc_hd__a31oi_2 _38579_ (.A1(_15922_),
    .A2(_15923_),
    .A3(_15924_),
    .B1(_15715_),
    .Y(_16524_));
 sky130_fd_sc_hd__inv_2 _38580_ (.A(_15921_),
    .Y(_16525_));
 sky130_fd_sc_hd__o2bb2ai_2 _38581_ (.A1_N(_16129_),
    .A2_N(_16126_),
    .B1(_16524_),
    .B2(_16525_),
    .Y(_16526_));
 sky130_fd_sc_hd__o21a_2 _38582_ (.A1(_16523_),
    .A2(_16526_),
    .B1(_16131_),
    .X(_16527_));
 sky130_fd_sc_hd__inv_2 _38583_ (.A(_16334_),
    .Y(_16528_));
 sky130_fd_sc_hd__o2bb2ai_2 _38584_ (.A1_N(_16330_),
    .A2_N(_16326_),
    .B1(_16328_),
    .B2(_16333_),
    .Y(_16529_));
 sky130_fd_sc_hd__o21a_2 _38585_ (.A1(_16528_),
    .A2(_16529_),
    .B1(_16332_),
    .X(_16530_));
 sky130_fd_sc_hd__a21boi_2 _38586_ (.A1(_16335_),
    .A2(_16334_),
    .B1_N(_16329_),
    .Y(_16531_));
 sky130_fd_sc_hd__o21ai_2 _38587_ (.A1(_16137_),
    .A2(_16531_),
    .B1(_16336_),
    .Y(_16532_));
 sky130_fd_sc_hd__a31oi_2 _38588_ (.A1(_16140_),
    .A2(_16527_),
    .A3(_16530_),
    .B1(_16532_),
    .Y(_16533_));
 sky130_fd_sc_hd__a21boi_2 _38589_ (.A1(_15747_),
    .A2(_16522_),
    .B1_N(_16533_),
    .Y(_16534_));
 sky130_fd_sc_hd__or2_2 _38590_ (.A(_16519_),
    .B(_16534_),
    .X(_16535_));
 sky130_fd_sc_hd__nand2_2 _38591_ (.A(_16534_),
    .B(_16519_),
    .Y(_16536_));
 sky130_fd_sc_hd__and2_2 _38592_ (.A(_16535_),
    .B(_16536_),
    .X(_02671_));
 sky130_fd_sc_hd__nand2_2 _38593_ (.A(_16455_),
    .B(_16462_),
    .Y(_16537_));
 sky130_fd_sc_hd__a21o_2 _38594_ (.A1(_16537_),
    .A2(_16461_),
    .B1(_15755_),
    .X(_16538_));
 sky130_fd_sc_hd__nand3_2 _38595_ (.A(_15756_),
    .B(_16537_),
    .C(_16461_),
    .Y(_16539_));
 sky130_fd_sc_hd__and2_2 _38596_ (.A(_16538_),
    .B(_16539_),
    .X(_16540_));
 sky130_fd_sc_hd__nand2_2 _38597_ (.A(_16540_),
    .B(_16093_),
    .Y(_16541_));
 sky130_fd_sc_hd__inv_2 _38598_ (.A(_16541_),
    .Y(_16542_));
 sky130_fd_sc_hd__nand2_2 _38599_ (.A(_16538_),
    .B(_16539_),
    .Y(_16543_));
 sky130_fd_sc_hd__nand2_2 _38600_ (.A(_16543_),
    .B(_16089_),
    .Y(_16544_));
 sky130_fd_sc_hd__inv_2 _38601_ (.A(_16544_),
    .Y(_16545_));
 sky130_fd_sc_hd__inv_2 _38602_ (.A(_16428_),
    .Y(_16546_));
 sky130_fd_sc_hd__nand2_2 _38603_ (.A(_16429_),
    .B(_16399_),
    .Y(_16547_));
 sky130_fd_sc_hd__o2bb2ai_2 _38604_ (.A1_N(_16432_),
    .A2_N(_16427_),
    .B1(_16546_),
    .B2(_16547_),
    .Y(_16548_));
 sky130_fd_sc_hd__a21o_2 _38605_ (.A1(_15451_),
    .A2(_15862_),
    .B1(_16446_),
    .X(_16549_));
 sky130_fd_sc_hd__nand2_2 _38606_ (.A(_16549_),
    .B(_16443_),
    .Y(_16550_));
 sky130_fd_sc_hd__and2_2 _38607_ (.A(_16423_),
    .B(_16414_),
    .X(_16551_));
 sky130_fd_sc_hd__nor2_2 _38608_ (.A(_16550_),
    .B(_16551_),
    .Y(_16552_));
 sky130_fd_sc_hd__and3_2 _38609_ (.A(_16550_),
    .B(_16414_),
    .C(_16423_),
    .X(_16553_));
 sky130_fd_sc_hd__o21ai_2 _38610_ (.A1(_16552_),
    .A2(_16553_),
    .B1(_15474_),
    .Y(_16554_));
 sky130_fd_sc_hd__nand2_2 _38611_ (.A(_16551_),
    .B(_16550_),
    .Y(_16555_));
 sky130_fd_sc_hd__nand3b_2 _38612_ (.A_N(_16552_),
    .B(_15585_),
    .C(_16555_),
    .Y(_16556_));
 sky130_fd_sc_hd__and2_2 _38613_ (.A(_16554_),
    .B(_16556_),
    .X(_16557_));
 sky130_fd_sc_hd__nand2_2 _38614_ (.A(_16548_),
    .B(_16557_),
    .Y(_16558_));
 sky130_fd_sc_hd__nand3_2 _38615_ (.A(_16427_),
    .B(_16431_),
    .C(_16432_),
    .Y(_16559_));
 sky130_fd_sc_hd__nand2_2 _38616_ (.A(_16554_),
    .B(_16556_),
    .Y(_16560_));
 sky130_fd_sc_hd__nand3_2 _38617_ (.A(_16559_),
    .B(_16431_),
    .C(_16560_),
    .Y(_16561_));
 sky130_fd_sc_hd__nand2_2 _38618_ (.A(_16451_),
    .B(_16458_),
    .Y(_16562_));
 sky130_fd_sc_hd__a21oi_2 _38619_ (.A1(_16558_),
    .A2(_16561_),
    .B1(_16562_),
    .Y(_16563_));
 sky130_fd_sc_hd__a21boi_2 _38620_ (.A1(_16548_),
    .A2(_16557_),
    .B1_N(_16562_),
    .Y(_16564_));
 sky130_fd_sc_hd__nand2_2 _38621_ (.A(_16564_),
    .B(_16561_),
    .Y(_16565_));
 sky130_fd_sc_hd__inv_2 _38622_ (.A(_16565_),
    .Y(_16566_));
 sky130_fd_sc_hd__nand2_2 _38623_ (.A(_18157_),
    .B(_19343_),
    .Y(_16567_));
 sky130_fd_sc_hd__nand2_2 _38624_ (.A(_19337_),
    .B(_11037_),
    .Y(_16568_));
 sky130_fd_sc_hd__nand2_2 _38625_ (.A(_09617_),
    .B(_11901_),
    .Y(_16569_));
 sky130_fd_sc_hd__nor2_2 _38626_ (.A(_16568_),
    .B(_16569_),
    .Y(_16570_));
 sky130_fd_sc_hd__and2_2 _38627_ (.A(_16568_),
    .B(_16569_),
    .X(_16571_));
 sky130_fd_sc_hd__or3_2 _38628_ (.A(_16567_),
    .B(_16570_),
    .C(_16571_),
    .X(_16572_));
 sky130_fd_sc_hd__nand2_2 _38629_ (.A(_16407_),
    .B(_16403_),
    .Y(_16573_));
 sky130_fd_sc_hd__o21ai_2 _38630_ (.A1(_16570_),
    .A2(_16571_),
    .B1(_16567_),
    .Y(_16574_));
 sky130_fd_sc_hd__and3_2 _38631_ (.A(_16572_),
    .B(_16573_),
    .C(_16574_),
    .X(_16575_));
 sky130_fd_sc_hd__a21o_2 _38632_ (.A1(_16572_),
    .A2(_16574_),
    .B1(_16573_),
    .X(_16576_));
 sky130_fd_sc_hd__nand2_2 _38633_ (.A(_16576_),
    .B(_16419_),
    .Y(_16577_));
 sky130_fd_sc_hd__nor2_2 _38634_ (.A(_16575_),
    .B(_16577_),
    .Y(_16578_));
 sky130_fd_sc_hd__and2_2 _38635_ (.A(_16572_),
    .B(_16574_),
    .X(_16579_));
 sky130_fd_sc_hd__nand2_2 _38636_ (.A(_16579_),
    .B(_16573_),
    .Y(_16580_));
 sky130_fd_sc_hd__a21oi_2 _38637_ (.A1(_16580_),
    .A2(_16576_),
    .B1(_16420_),
    .Y(_16581_));
 sky130_fd_sc_hd__a21boi_2 _38638_ (.A1(_16377_),
    .A2(_16378_),
    .B1_N(_16379_),
    .Y(_16582_));
 sky130_fd_sc_hd__o21ai_2 _38639_ (.A1(_16578_),
    .A2(_16581_),
    .B1(_16582_),
    .Y(_16583_));
 sky130_fd_sc_hd__a21o_2 _38640_ (.A1(_16580_),
    .A2(_16576_),
    .B1(_16419_),
    .X(_16584_));
 sky130_fd_sc_hd__nand2_2 _38641_ (.A(_16380_),
    .B(_16379_),
    .Y(_16585_));
 sky130_fd_sc_hd__nand3b_2 _38642_ (.A_N(_16578_),
    .B(_16584_),
    .C(_16585_),
    .Y(_16586_));
 sky130_fd_sc_hd__inv_2 _38643_ (.A(_16409_),
    .Y(_16587_));
 sky130_fd_sc_hd__and2_2 _38644_ (.A(_16411_),
    .B(_16419_),
    .X(_16588_));
 sky130_fd_sc_hd__nor2_2 _38645_ (.A(_16587_),
    .B(_16588_),
    .Y(_16589_));
 sky130_fd_sc_hd__inv_2 _38646_ (.A(_16589_),
    .Y(_16590_));
 sky130_fd_sc_hd__a21oi_2 _38647_ (.A1(_16583_),
    .A2(_16586_),
    .B1(_16590_),
    .Y(_16591_));
 sky130_fd_sc_hd__nand3_2 _38648_ (.A(_16590_),
    .B(_16583_),
    .C(_16586_),
    .Y(_16592_));
 sky130_fd_sc_hd__inv_2 _38649_ (.A(_16592_),
    .Y(_16593_));
 sky130_fd_sc_hd__nand2_2 _38650_ (.A(_16363_),
    .B(_16355_),
    .Y(_16594_));
 sky130_fd_sc_hd__o21bai_2 _38651_ (.A1(_16346_),
    .A2(_16348_),
    .B1_N(_16347_),
    .Y(_16595_));
 sky130_fd_sc_hd__and4_2 _38652_ (.A(_09678_),
    .B(_14356_),
    .C(_10700_),
    .D(_12349_),
    .X(_16596_));
 sky130_fd_sc_hd__o22a_2 _38653_ (.A1(_07845_),
    .A2(_13848_),
    .B1(_14855_),
    .B2(_14646_),
    .X(_16597_));
 sky130_fd_sc_hd__or2_2 _38654_ (.A(_16596_),
    .B(_16597_),
    .X(_16598_));
 sky130_fd_sc_hd__nor2_2 _38655_ (.A(_10151_),
    .B(_12090_),
    .Y(_16599_));
 sky130_fd_sc_hd__nand2_2 _38656_ (.A(_16598_),
    .B(_16599_),
    .Y(_16600_));
 sky130_fd_sc_hd__nor2_2 _38657_ (.A(_16596_),
    .B(_16597_),
    .Y(_16601_));
 sky130_fd_sc_hd__inv_2 _38658_ (.A(_16599_),
    .Y(_16602_));
 sky130_fd_sc_hd__nand2_2 _38659_ (.A(_16601_),
    .B(_16602_),
    .Y(_16603_));
 sky130_fd_sc_hd__nand3b_2 _38660_ (.A_N(_16595_),
    .B(_16600_),
    .C(_16603_),
    .Y(_16604_));
 sky130_fd_sc_hd__nand2_2 _38661_ (.A(_16598_),
    .B(_16602_),
    .Y(_16605_));
 sky130_fd_sc_hd__nand2_2 _38662_ (.A(_16601_),
    .B(_16599_),
    .Y(_16606_));
 sky130_fd_sc_hd__nand3_2 _38663_ (.A(_16605_),
    .B(_16595_),
    .C(_16606_),
    .Y(_16607_));
 sky130_fd_sc_hd__nor2_2 _38664_ (.A(_09358_),
    .B(_10523_),
    .Y(_16608_));
 sky130_fd_sc_hd__a22o_2 _38665_ (.A1(_10139_),
    .A2(_08922_),
    .B1(_19320_),
    .B2(_09219_),
    .X(_16609_));
 sky130_fd_sc_hd__o21a_2 _38666_ (.A1(_10705_),
    .A2(_12104_),
    .B1(_16609_),
    .X(_16610_));
 sky130_fd_sc_hd__nor2_2 _38667_ (.A(_16608_),
    .B(_16610_),
    .Y(_16611_));
 sky130_fd_sc_hd__and2_2 _38668_ (.A(_16610_),
    .B(_16608_),
    .X(_16612_));
 sky130_fd_sc_hd__nor2_2 _38669_ (.A(_16611_),
    .B(_16612_),
    .Y(_16613_));
 sky130_fd_sc_hd__nand3_2 _38670_ (.A(_16604_),
    .B(_16607_),
    .C(_16613_),
    .Y(_16614_));
 sky130_fd_sc_hd__a21o_2 _38671_ (.A1(_16604_),
    .A2(_16607_),
    .B1(_16613_),
    .X(_16615_));
 sky130_fd_sc_hd__nand3_2 _38672_ (.A(_16594_),
    .B(_16614_),
    .C(_16615_),
    .Y(_16616_));
 sky130_fd_sc_hd__nand2_2 _38673_ (.A(_16615_),
    .B(_16614_),
    .Y(_16617_));
 sky130_fd_sc_hd__a21boi_2 _38674_ (.A1(_16352_),
    .A2(_16361_),
    .B1_N(_16355_),
    .Y(_16618_));
 sky130_fd_sc_hd__nand2_2 _38675_ (.A(_16617_),
    .B(_16618_),
    .Y(_16619_));
 sky130_fd_sc_hd__and4_2 _38676_ (.A(_14569_),
    .B(_14068_),
    .C(_10050_),
    .D(_09733_),
    .X(_16620_));
 sky130_fd_sc_hd__o22a_2 _38677_ (.A1(_14571_),
    .A2(_13274_),
    .B1(_13873_),
    .B2(_10542_),
    .X(_16621_));
 sky130_fd_sc_hd__nor2_2 _38678_ (.A(_16620_),
    .B(_16621_),
    .Y(_16622_));
 sky130_fd_sc_hd__a21o_2 _38679_ (.A1(_19335_),
    .A2(_19551_),
    .B1(_16622_),
    .X(_16623_));
 sky130_fd_sc_hd__nand3_2 _38680_ (.A(_16622_),
    .B(_19335_),
    .C(_19551_),
    .Y(_16624_));
 sky130_fd_sc_hd__o21bai_2 _38681_ (.A1(_16356_),
    .A2(_16357_),
    .B1_N(_16358_),
    .Y(_16625_));
 sky130_fd_sc_hd__a21o_2 _38682_ (.A1(_16623_),
    .A2(_16624_),
    .B1(_16625_),
    .X(_16626_));
 sky130_fd_sc_hd__or2b_2 _38683_ (.A(_16370_),
    .B_N(_16373_),
    .X(_16627_));
 sky130_fd_sc_hd__nand3_2 _38684_ (.A(_16623_),
    .B(_16625_),
    .C(_16624_),
    .Y(_16628_));
 sky130_fd_sc_hd__nand3_2 _38685_ (.A(_16626_),
    .B(_16627_),
    .C(_16628_),
    .Y(_16629_));
 sky130_fd_sc_hd__inv_2 _38686_ (.A(_16629_),
    .Y(_16630_));
 sky130_fd_sc_hd__a21oi_2 _38687_ (.A1(_16623_),
    .A2(_16624_),
    .B1(_16625_),
    .Y(_16631_));
 sky130_fd_sc_hd__and3_2 _38688_ (.A(_16623_),
    .B(_16625_),
    .C(_16624_),
    .X(_16632_));
 sky130_fd_sc_hd__and2b_2 _38689_ (.A_N(_16370_),
    .B(_16373_),
    .X(_16633_));
 sky130_fd_sc_hd__o21ai_2 _38690_ (.A1(_16631_),
    .A2(_16632_),
    .B1(_16633_),
    .Y(_16634_));
 sky130_fd_sc_hd__inv_2 _38691_ (.A(_16634_),
    .Y(_16635_));
 sky130_fd_sc_hd__o2bb2ai_2 _38692_ (.A1_N(_16616_),
    .A2_N(_16619_),
    .B1(_16630_),
    .B2(_16635_),
    .Y(_16636_));
 sky130_fd_sc_hd__and2_2 _38693_ (.A(_16634_),
    .B(_16629_),
    .X(_16637_));
 sky130_fd_sc_hd__nand3_2 _38694_ (.A(_16637_),
    .B(_16619_),
    .C(_16616_),
    .Y(_16638_));
 sky130_fd_sc_hd__a21oi_2 _38695_ (.A1(_16362_),
    .A2(_16363_),
    .B1(_16344_),
    .Y(_16639_));
 sky130_fd_sc_hd__o21ai_2 _38696_ (.A1(_16388_),
    .A2(_16639_),
    .B1(_16364_),
    .Y(_16640_));
 sky130_fd_sc_hd__a21oi_2 _38697_ (.A1(_16636_),
    .A2(_16638_),
    .B1(_16640_),
    .Y(_16641_));
 sky130_fd_sc_hd__inv_2 _38698_ (.A(_16616_),
    .Y(_16642_));
 sky130_fd_sc_hd__nand2_2 _38699_ (.A(_16637_),
    .B(_16619_),
    .Y(_16643_));
 sky130_fd_sc_hd__o211a_2 _38700_ (.A1(_16642_),
    .A2(_16643_),
    .B1(_16640_),
    .C1(_16636_),
    .X(_16644_));
 sky130_fd_sc_hd__o22ai_2 _38701_ (.A1(_16591_),
    .A2(_16593_),
    .B1(_16641_),
    .B2(_16644_),
    .Y(_16645_));
 sky130_fd_sc_hd__a21oi_2 _38702_ (.A1(_16619_),
    .A2(_16616_),
    .B1(_16637_),
    .Y(_16646_));
 sky130_fd_sc_hd__a21oi_2 _38703_ (.A1(_16604_),
    .A2(_16607_),
    .B1(_16613_),
    .Y(_16647_));
 sky130_fd_sc_hd__nor2_2 _38704_ (.A(_16647_),
    .B(_16618_),
    .Y(_16648_));
 sky130_fd_sc_hd__nand2_2 _38705_ (.A(_16634_),
    .B(_16629_),
    .Y(_16649_));
 sky130_fd_sc_hd__a21oi_2 _38706_ (.A1(_16615_),
    .A2(_16614_),
    .B1(_16594_),
    .Y(_16650_));
 sky130_fd_sc_hd__a211oi_2 _38707_ (.A1(_16648_),
    .A2(_16614_),
    .B1(_16649_),
    .C1(_16650_),
    .Y(_16651_));
 sky130_fd_sc_hd__o21a_2 _38708_ (.A1(_16388_),
    .A2(_16639_),
    .B1(_16364_),
    .X(_16652_));
 sky130_fd_sc_hd__o21ai_2 _38709_ (.A1(_16646_),
    .A2(_16651_),
    .B1(_16652_),
    .Y(_16653_));
 sky130_fd_sc_hd__o21a_2 _38710_ (.A1(_16587_),
    .A2(_16588_),
    .B1(_16586_),
    .X(_16654_));
 sky130_fd_sc_hd__a21oi_2 _38711_ (.A1(_16654_),
    .A2(_16583_),
    .B1(_16591_),
    .Y(_16655_));
 sky130_fd_sc_hd__nand3_2 _38712_ (.A(_16636_),
    .B(_16640_),
    .C(_16638_),
    .Y(_16656_));
 sky130_fd_sc_hd__nand3_2 _38713_ (.A(_16653_),
    .B(_16655_),
    .C(_16656_),
    .Y(_16657_));
 sky130_fd_sc_hd__nand2_2 _38714_ (.A(_16397_),
    .B(_16434_),
    .Y(_16658_));
 sky130_fd_sc_hd__nand2_2 _38715_ (.A(_16658_),
    .B(_16390_),
    .Y(_16659_));
 sky130_fd_sc_hd__a21oi_2 _38716_ (.A1(_16645_),
    .A2(_16657_),
    .B1(_16659_),
    .Y(_16660_));
 sky130_fd_sc_hd__nand2_2 _38717_ (.A(_16653_),
    .B(_16655_),
    .Y(_16661_));
 sky130_fd_sc_hd__o211a_2 _38718_ (.A1(_16644_),
    .A2(_16661_),
    .B1(_16659_),
    .C1(_16645_),
    .X(_16662_));
 sky130_fd_sc_hd__o22ai_2 _38719_ (.A1(_16563_),
    .A2(_16566_),
    .B1(_16660_),
    .B2(_16662_),
    .Y(_16663_));
 sky130_fd_sc_hd__nand2_2 _38720_ (.A(_16583_),
    .B(_16586_),
    .Y(_16664_));
 sky130_fd_sc_hd__nand2_2 _38721_ (.A(_16664_),
    .B(_16589_),
    .Y(_16665_));
 sky130_fd_sc_hd__a22oi_2 _38722_ (.A1(_16665_),
    .A2(_16592_),
    .B1(_16653_),
    .B2(_16656_),
    .Y(_16666_));
 sky130_fd_sc_hd__nand2_2 _38723_ (.A(_16636_),
    .B(_16640_),
    .Y(_16667_));
 sky130_fd_sc_hd__o211a_2 _38724_ (.A1(_16651_),
    .A2(_16667_),
    .B1(_16655_),
    .C1(_16653_),
    .X(_16668_));
 sky130_fd_sc_hd__o21bai_2 _38725_ (.A1(_16666_),
    .A2(_16668_),
    .B1_N(_16659_),
    .Y(_16669_));
 sky130_fd_sc_hd__nand3_2 _38726_ (.A(_16645_),
    .B(_16659_),
    .C(_16657_),
    .Y(_16670_));
 sky130_fd_sc_hd__a21oi_2 _38727_ (.A1(_16561_),
    .A2(_16564_),
    .B1(_16563_),
    .Y(_16671_));
 sky130_fd_sc_hd__nand3_2 _38728_ (.A(_16669_),
    .B(_16670_),
    .C(_16671_),
    .Y(_16672_));
 sky130_fd_sc_hd__nand2_2 _38729_ (.A(_16442_),
    .B(_16468_),
    .Y(_16673_));
 sky130_fd_sc_hd__nand2_2 _38730_ (.A(_16673_),
    .B(_16438_),
    .Y(_16674_));
 sky130_fd_sc_hd__a21oi_2 _38731_ (.A1(_16663_),
    .A2(_16672_),
    .B1(_16674_),
    .Y(_16675_));
 sky130_fd_sc_hd__nand2_2 _38732_ (.A(_16669_),
    .B(_16671_),
    .Y(_16676_));
 sky130_fd_sc_hd__o211a_2 _38733_ (.A1(_16662_),
    .A2(_16676_),
    .B1(_16674_),
    .C1(_16663_),
    .X(_16677_));
 sky130_fd_sc_hd__o22ai_2 _38734_ (.A1(_16542_),
    .A2(_16545_),
    .B1(_16675_),
    .B2(_16677_),
    .Y(_16678_));
 sky130_fd_sc_hd__o21ai_2 _38735_ (.A1(_16481_),
    .A2(_16472_),
    .B1(_16489_),
    .Y(_16679_));
 sky130_fd_sc_hd__inv_2 _38736_ (.A(_16563_),
    .Y(_16680_));
 sky130_fd_sc_hd__a22oi_2 _38737_ (.A1(_16680_),
    .A2(_16565_),
    .B1(_16669_),
    .B2(_16670_),
    .Y(_16681_));
 sky130_fd_sc_hd__nand2_2 _38738_ (.A(_16680_),
    .B(_16565_),
    .Y(_16682_));
 sky130_fd_sc_hd__nor3_2 _38739_ (.A(_16682_),
    .B(_16660_),
    .C(_16662_),
    .Y(_16683_));
 sky130_fd_sc_hd__o21bai_2 _38740_ (.A1(_16681_),
    .A2(_16683_),
    .B1_N(_16674_),
    .Y(_16684_));
 sky130_fd_sc_hd__nand3_2 _38741_ (.A(_16663_),
    .B(_16674_),
    .C(_16672_),
    .Y(_16685_));
 sky130_fd_sc_hd__nand2_2 _38742_ (.A(_16543_),
    .B(_16294_),
    .Y(_16686_));
 sky130_fd_sc_hd__nand3_2 _38743_ (.A(_16538_),
    .B(_16539_),
    .C(_16089_),
    .Y(_16687_));
 sky130_fd_sc_hd__nand2_2 _38744_ (.A(_16686_),
    .B(_16687_),
    .Y(_16688_));
 sky130_fd_sc_hd__nand3_2 _38745_ (.A(_16684_),
    .B(_16685_),
    .C(_16688_),
    .Y(_16689_));
 sky130_fd_sc_hd__nand3_2 _38746_ (.A(_16678_),
    .B(_16679_),
    .C(_16689_),
    .Y(_16690_));
 sky130_fd_sc_hd__inv_2 _38747_ (.A(_16686_),
    .Y(_16691_));
 sky130_fd_sc_hd__inv_2 _38748_ (.A(_16687_),
    .Y(_16692_));
 sky130_fd_sc_hd__o22ai_2 _38749_ (.A1(_16691_),
    .A2(_16692_),
    .B1(_16675_),
    .B2(_16677_),
    .Y(_16693_));
 sky130_fd_sc_hd__o21a_2 _38750_ (.A1(_16473_),
    .A2(_16474_),
    .B1(_16466_),
    .X(_16694_));
 sky130_fd_sc_hd__a22oi_2 _38751_ (.A1(_16694_),
    .A2(_16469_),
    .B1(_16487_),
    .B2(_16488_),
    .Y(_16695_));
 sky130_fd_sc_hd__nand2_2 _38752_ (.A(_16541_),
    .B(_16544_),
    .Y(_16696_));
 sky130_fd_sc_hd__nand3_2 _38753_ (.A(_16684_),
    .B(_16685_),
    .C(_16696_),
    .Y(_16697_));
 sky130_fd_sc_hd__nand3_2 _38754_ (.A(_16693_),
    .B(_16695_),
    .C(_16697_),
    .Y(_16698_));
 sky130_fd_sc_hd__nand2_2 _38755_ (.A(_16478_),
    .B(_16476_),
    .Y(_16699_));
 sky130_fd_sc_hd__inv_2 _38756_ (.A(_16699_),
    .Y(_16700_));
 sky130_fd_sc_hd__nor2_2 _38757_ (.A(_15081_),
    .B(_16700_),
    .Y(_16701_));
 sky130_fd_sc_hd__nor2_2 _38758_ (.A(_14017_),
    .B(_16699_),
    .Y(_16702_));
 sky130_fd_sc_hd__o2bb2ai_2 _38759_ (.A1_N(_16690_),
    .A2_N(_16698_),
    .B1(_16701_),
    .B2(_16702_),
    .Y(_16703_));
 sky130_fd_sc_hd__a21boi_2 _38760_ (.A1(_16495_),
    .A2(_16501_),
    .B1_N(_16491_),
    .Y(_16704_));
 sky130_fd_sc_hd__nor2_2 _38761_ (.A(_16702_),
    .B(_16701_),
    .Y(_16705_));
 sky130_fd_sc_hd__nand3_2 _38762_ (.A(_16690_),
    .B(_16698_),
    .C(_16705_),
    .Y(_16706_));
 sky130_fd_sc_hd__nand3_2 _38763_ (.A(_16703_),
    .B(_16704_),
    .C(_16706_),
    .Y(_16707_));
 sky130_fd_sc_hd__nor2_2 _38764_ (.A(_16118_),
    .B(_16700_),
    .Y(_16708_));
 sky130_fd_sc_hd__nor2_2 _38765_ (.A(_16120_),
    .B(_16699_),
    .Y(_16709_));
 sky130_fd_sc_hd__o2bb2ai_2 _38766_ (.A1_N(_16690_),
    .A2_N(_16698_),
    .B1(_16708_),
    .B2(_16709_),
    .Y(_16710_));
 sky130_fd_sc_hd__nand2_2 _38767_ (.A(_16495_),
    .B(_16501_),
    .Y(_16711_));
 sky130_fd_sc_hd__nand2_2 _38768_ (.A(_16711_),
    .B(_16491_),
    .Y(_16712_));
 sky130_fd_sc_hd__inv_2 _38769_ (.A(_16705_),
    .Y(_16713_));
 sky130_fd_sc_hd__nand3_2 _38770_ (.A(_16690_),
    .B(_16698_),
    .C(_16713_),
    .Y(_16714_));
 sky130_fd_sc_hd__nand3_2 _38771_ (.A(_16710_),
    .B(_16712_),
    .C(_16714_),
    .Y(_16715_));
 sky130_fd_sc_hd__a21oi_2 _38772_ (.A1(_16707_),
    .A2(_16715_),
    .B1(_16500_),
    .Y(_16716_));
 sky130_fd_sc_hd__and3_2 _38773_ (.A(_16707_),
    .B(_16715_),
    .C(_16500_),
    .X(_16717_));
 sky130_fd_sc_hd__o21ai_2 _38774_ (.A1(_16506_),
    .A2(_16507_),
    .B1(_16509_),
    .Y(_16718_));
 sky130_fd_sc_hd__inv_2 _38775_ (.A(_16508_),
    .Y(_16719_));
 sky130_fd_sc_hd__o2bb2ai_2 _38776_ (.A1_N(_16322_),
    .A2_N(_16505_),
    .B1(_16718_),
    .B2(_16719_),
    .Y(_16720_));
 sky130_fd_sc_hd__o21bai_2 _38777_ (.A1(_16716_),
    .A2(_16717_),
    .B1_N(_16720_),
    .Y(_16721_));
 sky130_fd_sc_hd__o2bb2ai_2 _38778_ (.A1_N(_16715_),
    .A2_N(_16707_),
    .B1(_15729_),
    .B2(_16499_),
    .Y(_16722_));
 sky130_fd_sc_hd__nand3_2 _38779_ (.A(_16707_),
    .B(_16715_),
    .C(_16500_),
    .Y(_16723_));
 sky130_fd_sc_hd__nand3_2 _38780_ (.A(_16722_),
    .B(_16720_),
    .C(_16723_),
    .Y(_16724_));
 sky130_fd_sc_hd__a22o_2 _38781_ (.A1(_16721_),
    .A2(_16724_),
    .B1(_16535_),
    .B2(_16517_),
    .X(_16725_));
 sky130_fd_sc_hd__o2111ai_2 _38782_ (.A1(_16519_),
    .A2(_16534_),
    .B1(_16517_),
    .C1(_16721_),
    .D1(_16724_),
    .Y(_16726_));
 sky130_fd_sc_hd__nand2_2 _38783_ (.A(_16725_),
    .B(_16726_),
    .Y(_02672_));
 sky130_fd_sc_hd__a21oi_2 _38784_ (.A1(_16678_),
    .A2(_16689_),
    .B1(_16679_),
    .Y(_16727_));
 sky130_fd_sc_hd__o21ai_2 _38785_ (.A1(_16696_),
    .A2(_16675_),
    .B1(_16685_),
    .Y(_16728_));
 sky130_fd_sc_hd__nand2_2 _38786_ (.A(_16423_),
    .B(_16414_),
    .Y(_16729_));
 sky130_fd_sc_hd__a21o_2 _38787_ (.A1(_16423_),
    .A2(_16414_),
    .B1(_16443_),
    .X(_16730_));
 sky130_fd_sc_hd__o21ai_2 _38788_ (.A1(_16444_),
    .A2(_16729_),
    .B1(_16730_),
    .Y(_16731_));
 sky130_fd_sc_hd__nor2_2 _38789_ (.A(_16731_),
    .B(_15585_),
    .Y(_16732_));
 sky130_fd_sc_hd__and2_2 _38790_ (.A(_15584_),
    .B(_16731_),
    .X(_16733_));
 sky130_fd_sc_hd__or2_2 _38791_ (.A(_16732_),
    .B(_16733_),
    .X(_16734_));
 sky130_fd_sc_hd__a21o_2 _38792_ (.A1(_16592_),
    .A2(_16586_),
    .B1(_16734_),
    .X(_16735_));
 sky130_fd_sc_hd__buf_1 _38793_ (.A(_16734_),
    .X(_16736_));
 sky130_fd_sc_hd__nand3_2 _38794_ (.A(_16736_),
    .B(_16592_),
    .C(_16586_),
    .Y(_16737_));
 sky130_fd_sc_hd__nand2_2 _38795_ (.A(_16554_),
    .B(_16730_),
    .Y(_16738_));
 sky130_fd_sc_hd__a21oi_2 _38796_ (.A1(_16735_),
    .A2(_16737_),
    .B1(_16738_),
    .Y(_16739_));
 sky130_fd_sc_hd__nand3_2 _38797_ (.A(_16735_),
    .B(_16738_),
    .C(_16737_),
    .Y(_16740_));
 sky130_fd_sc_hd__inv_2 _38798_ (.A(_16740_),
    .Y(_16741_));
 sky130_fd_sc_hd__and4_2 _38799_ (.A(_14646_),
    .B(_14350_),
    .C(_14351_),
    .D(_10966_),
    .X(_16742_));
 sky130_fd_sc_hd__o22a_2 _38800_ (.A1(_19575_),
    .A2(_18183_),
    .B1(_14353_),
    .B2(_12090_),
    .X(_16743_));
 sky130_fd_sc_hd__a211o_2 _38801_ (.A1(_19314_),
    .A2(_19569_),
    .B1(_16742_),
    .C1(_16743_),
    .X(_16744_));
 sky130_fd_sc_hd__nand2_2 _38802_ (.A(_19313_),
    .B(_09223_),
    .Y(_16745_));
 sky130_fd_sc_hd__o21bai_2 _38803_ (.A1(_16742_),
    .A2(_16743_),
    .B1_N(_16745_),
    .Y(_16746_));
 sky130_fd_sc_hd__nand2_2 _38804_ (.A(_16744_),
    .B(_16746_),
    .Y(_16747_));
 sky130_fd_sc_hd__a22o_2 _38805_ (.A1(_14351_),
    .A2(_19575_),
    .B1(_11660_),
    .B2(_14350_),
    .X(_16748_));
 sky130_fd_sc_hd__a21oi_2 _38806_ (.A1(_16748_),
    .A2(_16599_),
    .B1(_16596_),
    .Y(_16749_));
 sky130_fd_sc_hd__inv_2 _38807_ (.A(_16749_),
    .Y(_16750_));
 sky130_fd_sc_hd__nand2_2 _38808_ (.A(_16747_),
    .B(_16750_),
    .Y(_16751_));
 sky130_fd_sc_hd__inv_2 _38809_ (.A(_16751_),
    .Y(_16752_));
 sky130_fd_sc_hd__or3_2 _38810_ (.A(_11178_),
    .B(_10514_),
    .C(_15159_),
    .X(_16753_));
 sky130_fd_sc_hd__a22o_2 _38811_ (.A1(_19317_),
    .A2(_08921_),
    .B1(_14042_),
    .B2(_10055_),
    .X(_16754_));
 sky130_fd_sc_hd__a22o_2 _38812_ (.A1(_19325_),
    .A2(_19560_),
    .B1(_16753_),
    .B2(_16754_),
    .X(_16755_));
 sky130_fd_sc_hd__nand2_2 _38813_ (.A(_19324_),
    .B(_19559_),
    .Y(_16756_));
 sky130_fd_sc_hd__nand3b_2 _38814_ (.A_N(_16756_),
    .B(_16753_),
    .C(_16754_),
    .Y(_16757_));
 sky130_fd_sc_hd__and2_2 _38815_ (.A(_16755_),
    .B(_16757_),
    .X(_16758_));
 sky130_fd_sc_hd__nand3_2 _38816_ (.A(_16744_),
    .B(_16746_),
    .C(_16749_),
    .Y(_16759_));
 sky130_fd_sc_hd__nand2_2 _38817_ (.A(_16758_),
    .B(_16759_),
    .Y(_16760_));
 sky130_fd_sc_hd__nand2_2 _38818_ (.A(_16751_),
    .B(_16759_),
    .Y(_16761_));
 sky130_fd_sc_hd__nand2_2 _38819_ (.A(_16755_),
    .B(_16757_),
    .Y(_16762_));
 sky130_fd_sc_hd__nand2_2 _38820_ (.A(_16761_),
    .B(_16762_),
    .Y(_16763_));
 sky130_fd_sc_hd__nand2_2 _38821_ (.A(_16614_),
    .B(_16607_),
    .Y(_16764_));
 sky130_fd_sc_hd__o211ai_2 _38822_ (.A1(_16752_),
    .A2(_16760_),
    .B1(_16763_),
    .C1(_16764_),
    .Y(_16765_));
 sky130_fd_sc_hd__nand2_2 _38823_ (.A(_16761_),
    .B(_16758_),
    .Y(_16766_));
 sky130_fd_sc_hd__a21boi_2 _38824_ (.A1(_16604_),
    .A2(_16613_),
    .B1_N(_16607_),
    .Y(_16767_));
 sky130_fd_sc_hd__nand3_2 _38825_ (.A(_16751_),
    .B(_16759_),
    .C(_16762_),
    .Y(_16768_));
 sky130_fd_sc_hd__nand3_2 _38826_ (.A(_16766_),
    .B(_16767_),
    .C(_16768_),
    .Y(_16769_));
 sky130_fd_sc_hd__and2b_2 _38827_ (.A_N(_16620_),
    .B(_16624_),
    .X(_16770_));
 sky130_fd_sc_hd__nand2_2 _38828_ (.A(_14569_),
    .B(_10050_),
    .Y(_16771_));
 sky130_fd_sc_hd__a21o_2 _38829_ (.A1(_19332_),
    .A2(_19550_),
    .B1(_16771_),
    .X(_16772_));
 sky130_fd_sc_hd__nand2_2 _38830_ (.A(_14068_),
    .B(_19549_),
    .Y(_16773_));
 sky130_fd_sc_hd__a21o_2 _38831_ (.A1(_19329_),
    .A2(_19554_),
    .B1(_16773_),
    .X(_16774_));
 sky130_fd_sc_hd__nand2_2 _38832_ (.A(_16772_),
    .B(_16774_),
    .Y(_16775_));
 sky130_fd_sc_hd__nor2_2 _38833_ (.A(_14339_),
    .B(_11764_),
    .Y(_16776_));
 sky130_fd_sc_hd__nand2_2 _38834_ (.A(_16775_),
    .B(_16776_),
    .Y(_16777_));
 sky130_fd_sc_hd__nand3b_2 _38835_ (.A_N(_16776_),
    .B(_16772_),
    .C(_16774_),
    .Y(_16778_));
 sky130_fd_sc_hd__a2bb2o_2 _38836_ (.A1_N(_16003_),
    .A2_N(_12104_),
    .B1(_16609_),
    .B2(_16608_),
    .X(_16779_));
 sky130_fd_sc_hd__a21o_2 _38837_ (.A1(_16777_),
    .A2(_16778_),
    .B1(_16779_),
    .X(_16780_));
 sky130_fd_sc_hd__nand3_2 _38838_ (.A(_16779_),
    .B(_16777_),
    .C(_16778_),
    .Y(_16781_));
 sky130_fd_sc_hd__nand2_2 _38839_ (.A(_16780_),
    .B(_16781_),
    .Y(_16782_));
 sky130_fd_sc_hd__nor2_2 _38840_ (.A(_16770_),
    .B(_16782_),
    .Y(_16783_));
 sky130_fd_sc_hd__and2_2 _38841_ (.A(_16782_),
    .B(_16770_),
    .X(_16784_));
 sky130_fd_sc_hd__nor2_2 _38842_ (.A(_16783_),
    .B(_16784_),
    .Y(_16785_));
 sky130_fd_sc_hd__a21o_2 _38843_ (.A1(_16765_),
    .A2(_16769_),
    .B1(_16785_),
    .X(_16786_));
 sky130_fd_sc_hd__nand3_2 _38844_ (.A(_16765_),
    .B(_16769_),
    .C(_16785_),
    .Y(_16787_));
 sky130_fd_sc_hd__o21ai_2 _38845_ (.A1(_16649_),
    .A2(_16650_),
    .B1(_16616_),
    .Y(_16788_));
 sky130_fd_sc_hd__a21oi_2 _38846_ (.A1(_16786_),
    .A2(_16787_),
    .B1(_16788_),
    .Y(_16789_));
 sky130_fd_sc_hd__inv_2 _38847_ (.A(_16765_),
    .Y(_16790_));
 sky130_fd_sc_hd__nand2_2 _38848_ (.A(_16769_),
    .B(_16785_),
    .Y(_16791_));
 sky130_fd_sc_hd__o211a_2 _38849_ (.A1(_16790_),
    .A2(_16791_),
    .B1(_16786_),
    .C1(_16788_),
    .X(_16792_));
 sky130_fd_sc_hd__nand2_2 _38850_ (.A(_18157_),
    .B(_19341_),
    .Y(_16793_));
 sky130_fd_sc_hd__xor2_2 _38851_ (.A(_16567_),
    .B(_16793_),
    .X(_16794_));
 sky130_fd_sc_hd__nand3b_2 _38852_ (.A_N(_16794_),
    .B(_19338_),
    .C(_19543_),
    .Y(_16795_));
 sky130_fd_sc_hd__o21ai_2 _38853_ (.A1(_14645_),
    .A2(_15116_),
    .B1(_16794_),
    .Y(_16796_));
 sky130_fd_sc_hd__o21ba_2 _38854_ (.A1(_16567_),
    .A2(_16571_),
    .B1_N(_16570_),
    .X(_16797_));
 sky130_fd_sc_hd__a21o_2 _38855_ (.A1(_16795_),
    .A2(_16796_),
    .B1(_16797_),
    .X(_16798_));
 sky130_fd_sc_hd__nand3_2 _38856_ (.A(_16795_),
    .B(_16797_),
    .C(_16796_),
    .Y(_16799_));
 sky130_fd_sc_hd__a21o_2 _38857_ (.A1(_16798_),
    .A2(_16799_),
    .B1(_16420_),
    .X(_16800_));
 sky130_fd_sc_hd__nand3_2 _38858_ (.A(_16798_),
    .B(_16420_),
    .C(_16799_),
    .Y(_16801_));
 sky130_fd_sc_hd__o21ai_2 _38859_ (.A1(_16633_),
    .A2(_16631_),
    .B1(_16628_),
    .Y(_16802_));
 sky130_fd_sc_hd__a21oi_2 _38860_ (.A1(_16800_),
    .A2(_16801_),
    .B1(_16802_),
    .Y(_16803_));
 sky130_fd_sc_hd__and3_2 _38861_ (.A(_16800_),
    .B(_16802_),
    .C(_16801_),
    .X(_16804_));
 sky130_fd_sc_hd__nand2_2 _38862_ (.A(_16577_),
    .B(_16580_),
    .Y(_16805_));
 sky130_fd_sc_hd__o21bai_2 _38863_ (.A1(_16803_),
    .A2(_16804_),
    .B1_N(_16805_),
    .Y(_16806_));
 sky130_fd_sc_hd__a21o_2 _38864_ (.A1(_16800_),
    .A2(_16801_),
    .B1(_16802_),
    .X(_16807_));
 sky130_fd_sc_hd__nand3_2 _38865_ (.A(_16800_),
    .B(_16802_),
    .C(_16801_),
    .Y(_16808_));
 sky130_fd_sc_hd__nand3_2 _38866_ (.A(_16807_),
    .B(_16805_),
    .C(_16808_),
    .Y(_16809_));
 sky130_fd_sc_hd__nand2_2 _38867_ (.A(_16806_),
    .B(_16809_),
    .Y(_16810_));
 sky130_fd_sc_hd__o21ai_2 _38868_ (.A1(_16789_),
    .A2(_16792_),
    .B1(_16810_),
    .Y(_16811_));
 sky130_fd_sc_hd__a21o_2 _38869_ (.A1(_16786_),
    .A2(_16787_),
    .B1(_16788_),
    .X(_16812_));
 sky130_fd_sc_hd__nand3_2 _38870_ (.A(_16788_),
    .B(_16786_),
    .C(_16787_),
    .Y(_16813_));
 sky130_fd_sc_hd__nand3b_2 _38871_ (.A_N(_16810_),
    .B(_16812_),
    .C(_16813_),
    .Y(_16814_));
 sky130_fd_sc_hd__nand2_2 _38872_ (.A(_16665_),
    .B(_16592_),
    .Y(_16815_));
 sky130_fd_sc_hd__o21ai_2 _38873_ (.A1(_16815_),
    .A2(_16641_),
    .B1(_16656_),
    .Y(_16816_));
 sky130_fd_sc_hd__a21oi_2 _38874_ (.A1(_16811_),
    .A2(_16814_),
    .B1(_16816_),
    .Y(_16817_));
 sky130_fd_sc_hd__nand2_2 _38875_ (.A(_16636_),
    .B(_16638_),
    .Y(_16818_));
 sky130_fd_sc_hd__a21oi_2 _38876_ (.A1(_16818_),
    .A2(_16652_),
    .B1(_16815_),
    .Y(_16819_));
 sky130_fd_sc_hd__o211a_2 _38877_ (.A1(_16644_),
    .A2(_16819_),
    .B1(_16814_),
    .C1(_16811_),
    .X(_16820_));
 sky130_fd_sc_hd__o22ai_2 _38878_ (.A1(_16739_),
    .A2(_16741_),
    .B1(_16817_),
    .B2(_16820_),
    .Y(_16821_));
 sky130_fd_sc_hd__a31oi_2 _38879_ (.A1(_16645_),
    .A2(_16659_),
    .A3(_16657_),
    .B1(_16671_),
    .Y(_16822_));
 sky130_fd_sc_hd__nor2_2 _38880_ (.A(_16660_),
    .B(_16822_),
    .Y(_16823_));
 sky130_fd_sc_hd__nor2_2 _38881_ (.A(_16739_),
    .B(_16741_),
    .Y(_16824_));
 sky130_fd_sc_hd__nand2_2 _38882_ (.A(_16811_),
    .B(_16814_),
    .Y(_16825_));
 sky130_fd_sc_hd__nor2_2 _38883_ (.A(_16644_),
    .B(_16819_),
    .Y(_16826_));
 sky130_fd_sc_hd__nand2_2 _38884_ (.A(_16825_),
    .B(_16826_),
    .Y(_16827_));
 sky130_fd_sc_hd__nand3_2 _38885_ (.A(_16816_),
    .B(_16811_),
    .C(_16814_),
    .Y(_16828_));
 sky130_fd_sc_hd__nand3_2 _38886_ (.A(_16824_),
    .B(_16827_),
    .C(_16828_),
    .Y(_16829_));
 sky130_fd_sc_hd__nand3_2 _38887_ (.A(_16821_),
    .B(_16823_),
    .C(_16829_),
    .Y(_16830_));
 sky130_fd_sc_hd__o21ai_2 _38888_ (.A1(_16817_),
    .A2(_16820_),
    .B1(_16824_),
    .Y(_16831_));
 sky130_fd_sc_hd__nand2_2 _38889_ (.A(_16670_),
    .B(_16682_),
    .Y(_16832_));
 sky130_fd_sc_hd__nand2_2 _38890_ (.A(_16832_),
    .B(_16669_),
    .Y(_16833_));
 sky130_fd_sc_hd__a21o_2 _38891_ (.A1(_16735_),
    .A2(_16737_),
    .B1(_16738_),
    .X(_16834_));
 sky130_fd_sc_hd__nand2_2 _38892_ (.A(_16834_),
    .B(_16740_),
    .Y(_16835_));
 sky130_fd_sc_hd__nand3_2 _38893_ (.A(_16827_),
    .B(_16835_),
    .C(_16828_),
    .Y(_16836_));
 sky130_fd_sc_hd__nand3_2 _38894_ (.A(_16831_),
    .B(_16833_),
    .C(_16836_),
    .Y(_16837_));
 sky130_fd_sc_hd__nand2_2 _38895_ (.A(_16565_),
    .B(_16558_),
    .Y(_16838_));
 sky130_fd_sc_hd__nor2_2 _38896_ (.A(_15753_),
    .B(_16287_),
    .Y(_16839_));
 sky130_fd_sc_hd__nand2_2 _38897_ (.A(_16838_),
    .B(_16839_),
    .Y(_16840_));
 sky130_fd_sc_hd__nand3_2 _38898_ (.A(_16565_),
    .B(_15756_),
    .C(_16558_),
    .Y(_16841_));
 sky130_fd_sc_hd__nand2_2 _38899_ (.A(_16840_),
    .B(_16841_),
    .Y(_16842_));
 sky130_fd_sc_hd__nor2_2 _38900_ (.A(_16089_),
    .B(_16842_),
    .Y(_16843_));
 sky130_fd_sc_hd__buf_1 _38901_ (.A(_16093_),
    .X(_16844_));
 sky130_fd_sc_hd__inv_2 _38902_ (.A(_16842_),
    .Y(_16845_));
 sky130_fd_sc_hd__nor2_2 _38903_ (.A(_16844_),
    .B(_16845_),
    .Y(_16846_));
 sky130_fd_sc_hd__o2bb2ai_2 _38904_ (.A1_N(_16830_),
    .A2_N(_16837_),
    .B1(_16843_),
    .B2(_16846_),
    .Y(_16847_));
 sky130_fd_sc_hd__nand2_2 _38905_ (.A(_16842_),
    .B(_16293_),
    .Y(_16848_));
 sky130_fd_sc_hd__nand3_2 _38906_ (.A(_16840_),
    .B(_16088_),
    .C(_16841_),
    .Y(_16849_));
 sky130_fd_sc_hd__nand2_2 _38907_ (.A(_16848_),
    .B(_16849_),
    .Y(_16850_));
 sky130_fd_sc_hd__nand3_2 _38908_ (.A(_16837_),
    .B(_16830_),
    .C(_16850_),
    .Y(_16851_));
 sky130_fd_sc_hd__nand3_2 _38909_ (.A(_16728_),
    .B(_16847_),
    .C(_16851_),
    .Y(_16852_));
 sky130_fd_sc_hd__nand2_2 _38910_ (.A(_16685_),
    .B(_16696_),
    .Y(_16853_));
 sky130_fd_sc_hd__nand2_2 _38911_ (.A(_16853_),
    .B(_16684_),
    .Y(_16854_));
 sky130_fd_sc_hd__inv_2 _38912_ (.A(_16848_),
    .Y(_16855_));
 sky130_fd_sc_hd__inv_2 _38913_ (.A(_16849_),
    .Y(_16856_));
 sky130_fd_sc_hd__o2bb2ai_2 _38914_ (.A1_N(_16830_),
    .A2_N(_16837_),
    .B1(_16855_),
    .B2(_16856_),
    .Y(_16857_));
 sky130_fd_sc_hd__nand3b_2 _38915_ (.A_N(_16850_),
    .B(_16837_),
    .C(_16830_),
    .Y(_16858_));
 sky130_fd_sc_hd__nand3_2 _38916_ (.A(_16854_),
    .B(_16857_),
    .C(_16858_),
    .Y(_16859_));
 sky130_fd_sc_hd__nand2_2 _38917_ (.A(_16539_),
    .B(_16293_),
    .Y(_16860_));
 sky130_fd_sc_hd__nand2_2 _38918_ (.A(_16860_),
    .B(_16538_),
    .Y(_16861_));
 sky130_fd_sc_hd__nor2_2 _38919_ (.A(_14823_),
    .B(_16861_),
    .Y(_16862_));
 sky130_fd_sc_hd__inv_2 _38920_ (.A(_16861_),
    .Y(_16863_));
 sky130_fd_sc_hd__nor2_2 _38921_ (.A(_15081_),
    .B(_16863_),
    .Y(_16864_));
 sky130_fd_sc_hd__nor2_2 _38922_ (.A(_16862_),
    .B(_16864_),
    .Y(_16865_));
 sky130_fd_sc_hd__nand3_2 _38923_ (.A(_16852_),
    .B(_16859_),
    .C(_16865_),
    .Y(_16866_));
 sky130_fd_sc_hd__o2bb2ai_2 _38924_ (.A1_N(_16859_),
    .A2_N(_16852_),
    .B1(_16862_),
    .B2(_16864_),
    .Y(_16867_));
 sky130_fd_sc_hd__o2111ai_2 _38925_ (.A1(_16705_),
    .A2(_16727_),
    .B1(_16690_),
    .C1(_16866_),
    .D1(_16867_),
    .Y(_16868_));
 sky130_fd_sc_hd__a21oi_2 _38926_ (.A1(_16693_),
    .A2(_16697_),
    .B1(_16695_),
    .Y(_16869_));
 sky130_fd_sc_hd__a31oi_2 _38927_ (.A1(_16693_),
    .A2(_16695_),
    .A3(_16697_),
    .B1(_16705_),
    .Y(_16870_));
 sky130_fd_sc_hd__inv_2 _38928_ (.A(_16865_),
    .Y(_16871_));
 sky130_fd_sc_hd__nand3_2 _38929_ (.A(_16852_),
    .B(_16859_),
    .C(_16871_),
    .Y(_16872_));
 sky130_fd_sc_hd__nand2_2 _38930_ (.A(_16861_),
    .B(_15109_),
    .Y(_16873_));
 sky130_fd_sc_hd__inv_2 _38931_ (.A(_16873_),
    .Y(_16874_));
 sky130_fd_sc_hd__nor2_2 _38932_ (.A(_16120_),
    .B(_16861_),
    .Y(_16875_));
 sky130_fd_sc_hd__o2bb2ai_2 _38933_ (.A1_N(_16859_),
    .A2_N(_16852_),
    .B1(_16874_),
    .B2(_16875_),
    .Y(_16876_));
 sky130_fd_sc_hd__o211ai_2 _38934_ (.A1(_16869_),
    .A2(_16870_),
    .B1(_16872_),
    .C1(_16876_),
    .Y(_16877_));
 sky130_fd_sc_hd__buf_1 _38935_ (.A(_16708_),
    .X(_16878_));
 sky130_fd_sc_hd__a21oi_2 _38936_ (.A1(_16868_),
    .A2(_16877_),
    .B1(_16878_),
    .Y(_16879_));
 sky130_fd_sc_hd__and3_2 _38937_ (.A(_16868_),
    .B(_16877_),
    .C(_16878_),
    .X(_16880_));
 sky130_fd_sc_hd__a21oi_2 _38938_ (.A1(_16690_),
    .A2(_16698_),
    .B1(_16713_),
    .Y(_16881_));
 sky130_fd_sc_hd__nand2_2 _38939_ (.A(_16712_),
    .B(_16714_),
    .Y(_16882_));
 sky130_fd_sc_hd__o2bb2ai_2 _38940_ (.A1_N(_16500_),
    .A2_N(_16707_),
    .B1(_16881_),
    .B2(_16882_),
    .Y(_16883_));
 sky130_fd_sc_hd__o21bai_2 _38941_ (.A1(_16879_),
    .A2(_16880_),
    .B1_N(_16883_),
    .Y(_16884_));
 sky130_fd_sc_hd__a21o_2 _38942_ (.A1(_16868_),
    .A2(_16877_),
    .B1(_16878_),
    .X(_16885_));
 sky130_fd_sc_hd__nand3_2 _38943_ (.A(_16868_),
    .B(_16877_),
    .C(_16878_),
    .Y(_16886_));
 sky130_fd_sc_hd__nand3_2 _38944_ (.A(_16885_),
    .B(_16883_),
    .C(_16886_),
    .Y(_16887_));
 sky130_fd_sc_hd__and2_2 _38945_ (.A(_16884_),
    .B(_16887_),
    .X(_16888_));
 sky130_fd_sc_hd__nand2_2 _38946_ (.A(_16722_),
    .B(_16720_),
    .Y(_16889_));
 sky130_fd_sc_hd__o2111a_2 _38947_ (.A1(_16717_),
    .A2(_16889_),
    .B1(_16514_),
    .C1(_16517_),
    .D1(_16721_),
    .X(_16890_));
 sky130_fd_sc_hd__inv_2 _38948_ (.A(_16890_),
    .Y(_16891_));
 sky130_fd_sc_hd__nand2_2 _38949_ (.A(_16724_),
    .B(_16517_),
    .Y(_16892_));
 sky130_fd_sc_hd__nand2_2 _38950_ (.A(_16892_),
    .B(_16721_),
    .Y(_16893_));
 sky130_fd_sc_hd__o21ai_2 _38951_ (.A1(_16891_),
    .A2(_16534_),
    .B1(_16893_),
    .Y(_16894_));
 sky130_fd_sc_hd__or2_2 _38952_ (.A(_16888_),
    .B(_16894_),
    .X(_16895_));
 sky130_fd_sc_hd__nand2_2 _38953_ (.A(_16894_),
    .B(_16888_),
    .Y(_16896_));
 sky130_fd_sc_hd__and2_2 _38954_ (.A(_16895_),
    .B(_16896_),
    .X(_02673_));
 sky130_fd_sc_hd__a21o_2 _38955_ (.A1(_16809_),
    .A2(_16808_),
    .B1(_16736_),
    .X(_16897_));
 sky130_fd_sc_hd__nand3_2 _38956_ (.A(_16736_),
    .B(_16809_),
    .C(_16808_),
    .Y(_16898_));
 sky130_fd_sc_hd__nor2_2 _38957_ (.A(_16444_),
    .B(_16729_),
    .Y(_16899_));
 sky130_fd_sc_hd__and2_2 _38958_ (.A(_15886_),
    .B(_16730_),
    .X(_16900_));
 sky130_fd_sc_hd__nor2_2 _38959_ (.A(_16899_),
    .B(_16900_),
    .Y(_16901_));
 sky130_fd_sc_hd__buf_1 _38960_ (.A(_16901_),
    .X(_16902_));
 sky130_fd_sc_hd__a21oi_2 _38961_ (.A1(_16897_),
    .A2(_16898_),
    .B1(_16902_),
    .Y(_16903_));
 sky130_fd_sc_hd__and3_2 _38962_ (.A(_16897_),
    .B(_16898_),
    .C(_16901_),
    .X(_16904_));
 sky130_fd_sc_hd__a21o_2 _38963_ (.A1(_19341_),
    .A2(_19344_),
    .B1(_15116_),
    .X(_16905_));
 sky130_fd_sc_hd__nand2_2 _38964_ (.A(_14097_),
    .B(_12602_),
    .Y(_16906_));
 sky130_fd_sc_hd__a31o_2 _38965_ (.A1(_14645_),
    .A2(_14097_),
    .A3(_12602_),
    .B1(_11913_),
    .X(_16907_));
 sky130_fd_sc_hd__a31o_2 _38966_ (.A1(_19338_),
    .A2(_16905_),
    .A3(_16906_),
    .B1(_16907_),
    .X(_16908_));
 sky130_fd_sc_hd__or2_2 _38967_ (.A(_16908_),
    .B(_16425_),
    .X(_16909_));
 sky130_fd_sc_hd__nand2_2 _38968_ (.A(_16425_),
    .B(_16908_),
    .Y(_16910_));
 sky130_fd_sc_hd__a21oi_2 _38969_ (.A1(_16777_),
    .A2(_16778_),
    .B1(_16779_),
    .Y(_16911_));
 sky130_fd_sc_hd__o21ai_2 _38970_ (.A1(_16911_),
    .A2(_16770_),
    .B1(_16781_),
    .Y(_16912_));
 sky130_fd_sc_hd__a21o_2 _38971_ (.A1(_16909_),
    .A2(_16910_),
    .B1(_16912_),
    .X(_16913_));
 sky130_fd_sc_hd__nand3_2 _38972_ (.A(_16912_),
    .B(_16909_),
    .C(_16910_),
    .Y(_16914_));
 sky130_fd_sc_hd__nand2_2 _38973_ (.A(_16801_),
    .B(_16798_),
    .Y(_16915_));
 sky130_fd_sc_hd__a21oi_2 _38974_ (.A1(_16913_),
    .A2(_16914_),
    .B1(_16915_),
    .Y(_16916_));
 sky130_fd_sc_hd__and3_2 _38975_ (.A(_16913_),
    .B(_16915_),
    .C(_16914_),
    .X(_16917_));
 sky130_fd_sc_hd__nand2_2 _38976_ (.A(_16760_),
    .B(_16751_),
    .Y(_16918_));
 sky130_fd_sc_hd__inv_2 _38977_ (.A(_16742_),
    .Y(_16919_));
 sky130_fd_sc_hd__o21ai_2 _38978_ (.A1(_16745_),
    .A2(_16743_),
    .B1(_16919_),
    .Y(_16920_));
 sky130_fd_sc_hd__and4_2 _38979_ (.A(_12089_),
    .B(_11122_),
    .C(_14351_),
    .D(_19568_),
    .X(_16921_));
 sky130_fd_sc_hd__o22a_2 _38980_ (.A1(_10966_),
    .A2(_13848_),
    .B1(_14353_),
    .B2(_10485_),
    .X(_16922_));
 sky130_fd_sc_hd__or2_2 _38981_ (.A(_16921_),
    .B(_16922_),
    .X(_16923_));
 sky130_fd_sc_hd__nand2_2 _38982_ (.A(_19313_),
    .B(_08921_),
    .Y(_16924_));
 sky130_fd_sc_hd__inv_2 _38983_ (.A(_16924_),
    .Y(_16925_));
 sky130_fd_sc_hd__nand2_2 _38984_ (.A(_16923_),
    .B(_16925_),
    .Y(_16926_));
 sky130_fd_sc_hd__or3_2 _38985_ (.A(_16925_),
    .B(_16921_),
    .C(_16922_),
    .X(_16927_));
 sky130_fd_sc_hd__nand3b_2 _38986_ (.A_N(_16920_),
    .B(_16926_),
    .C(_16927_),
    .Y(_16928_));
 sky130_fd_sc_hd__nand2_2 _38987_ (.A(_16923_),
    .B(_16924_),
    .Y(_16929_));
 sky130_fd_sc_hd__or3_2 _38988_ (.A(_16924_),
    .B(_16921_),
    .C(_16922_),
    .X(_16930_));
 sky130_fd_sc_hd__nand3_2 _38989_ (.A(_16929_),
    .B(_16930_),
    .C(_16920_),
    .Y(_16931_));
 sky130_fd_sc_hd__nand2_2 _38990_ (.A(_15778_),
    .B(_19555_),
    .Y(_16932_));
 sky130_fd_sc_hd__inv_2 _38991_ (.A(_16932_),
    .Y(_16933_));
 sky130_fd_sc_hd__o22a_2 _38992_ (.A1(_14371_),
    .A2(_10514_),
    .B1(_14869_),
    .B2(_13274_),
    .X(_16934_));
 sky130_fd_sc_hd__and3_2 _38993_ (.A(_15781_),
    .B(_19559_),
    .C(_19563_),
    .X(_16935_));
 sky130_fd_sc_hd__nor2_2 _38994_ (.A(_16934_),
    .B(_16935_),
    .Y(_16936_));
 sky130_fd_sc_hd__nor2_2 _38995_ (.A(_16933_),
    .B(_16936_),
    .Y(_16937_));
 sky130_fd_sc_hd__a31o_2 _38996_ (.A1(_19560_),
    .A2(_19563_),
    .A3(_15781_),
    .B1(_16934_),
    .X(_16938_));
 sky130_fd_sc_hd__nor2_2 _38997_ (.A(_16932_),
    .B(_16938_),
    .Y(_16939_));
 sky130_fd_sc_hd__nor2_2 _38998_ (.A(_16937_),
    .B(_16939_),
    .Y(_16940_));
 sky130_fd_sc_hd__a21o_2 _38999_ (.A1(_16928_),
    .A2(_16931_),
    .B1(_16940_),
    .X(_16941_));
 sky130_fd_sc_hd__nand3_2 _39000_ (.A(_16940_),
    .B(_16928_),
    .C(_16931_),
    .Y(_16942_));
 sky130_fd_sc_hd__nand3_2 _39001_ (.A(_16918_),
    .B(_16941_),
    .C(_16942_),
    .Y(_16943_));
 sky130_fd_sc_hd__a21oi_2 _39002_ (.A1(_16928_),
    .A2(_16931_),
    .B1(_16940_),
    .Y(_16944_));
 sky130_fd_sc_hd__nor2_2 _39003_ (.A(_16933_),
    .B(_16938_),
    .Y(_16945_));
 sky130_fd_sc_hd__nor2_2 _39004_ (.A(_16932_),
    .B(_16936_),
    .Y(_16946_));
 sky130_fd_sc_hd__o211a_2 _39005_ (.A1(_16945_),
    .A2(_16946_),
    .B1(_16931_),
    .C1(_16928_),
    .X(_16947_));
 sky130_fd_sc_hd__a21oi_2 _39006_ (.A1(_16758_),
    .A2(_16759_),
    .B1(_16752_),
    .Y(_16948_));
 sky130_fd_sc_hd__o21ai_2 _39007_ (.A1(_16944_),
    .A2(_16947_),
    .B1(_16948_),
    .Y(_16949_));
 sky130_fd_sc_hd__nand2_2 _39008_ (.A(_19335_),
    .B(_19542_),
    .Y(_16950_));
 sky130_fd_sc_hd__and4_2 _39009_ (.A(_14569_),
    .B(_14068_),
    .C(_19545_),
    .D(_10371_),
    .X(_16951_));
 sky130_fd_sc_hd__a22o_2 _39010_ (.A1(_14569_),
    .A2(_10371_),
    .B1(_19332_),
    .B2(_11038_),
    .X(_16952_));
 sky130_fd_sc_hd__or3b_2 _39011_ (.A(_16950_),
    .B(_16951_),
    .C_N(_16952_),
    .X(_16953_));
 sky130_fd_sc_hd__inv_2 _39012_ (.A(_16952_),
    .Y(_16954_));
 sky130_fd_sc_hd__o21ai_2 _39013_ (.A1(_16951_),
    .A2(_16954_),
    .B1(_16950_),
    .Y(_16955_));
 sky130_fd_sc_hd__nand2_2 _39014_ (.A(_16953_),
    .B(_16955_),
    .Y(_16956_));
 sky130_fd_sc_hd__a21o_2 _39015_ (.A1(_16753_),
    .A2(_16757_),
    .B1(_16956_),
    .X(_16957_));
 sky130_fd_sc_hd__and2_2 _39016_ (.A(_16757_),
    .B(_16753_),
    .X(_16958_));
 sky130_fd_sc_hd__nand2_2 _39017_ (.A(_16958_),
    .B(_16956_),
    .Y(_16959_));
 sky130_fd_sc_hd__nor2_2 _39018_ (.A(_16771_),
    .B(_16773_),
    .Y(_16960_));
 sky130_fd_sc_hd__inv_2 _39019_ (.A(_16777_),
    .Y(_16961_));
 sky130_fd_sc_hd__nor2_2 _39020_ (.A(_16960_),
    .B(_16961_),
    .Y(_16962_));
 sky130_fd_sc_hd__inv_2 _39021_ (.A(_16962_),
    .Y(_16963_));
 sky130_fd_sc_hd__a21oi_2 _39022_ (.A1(_16957_),
    .A2(_16959_),
    .B1(_16963_),
    .Y(_16964_));
 sky130_fd_sc_hd__nand2_2 _39023_ (.A(_16957_),
    .B(_16959_),
    .Y(_16965_));
 sky130_fd_sc_hd__nor2_2 _39024_ (.A(_16962_),
    .B(_16965_),
    .Y(_16966_));
 sky130_fd_sc_hd__o2bb2ai_2 _39025_ (.A1_N(_16943_),
    .A2_N(_16949_),
    .B1(_16964_),
    .B2(_16966_),
    .Y(_16967_));
 sky130_fd_sc_hd__nand2_2 _39026_ (.A(_16965_),
    .B(_16963_),
    .Y(_16968_));
 sky130_fd_sc_hd__nand3_2 _39027_ (.A(_16957_),
    .B(_16962_),
    .C(_16959_),
    .Y(_16969_));
 sky130_fd_sc_hd__nand2_2 _39028_ (.A(_16968_),
    .B(_16969_),
    .Y(_16970_));
 sky130_fd_sc_hd__nand3_2 _39029_ (.A(_16970_),
    .B(_16943_),
    .C(_16949_),
    .Y(_16971_));
 sky130_fd_sc_hd__nand2_2 _39030_ (.A(_16791_),
    .B(_16765_),
    .Y(_16972_));
 sky130_fd_sc_hd__a21oi_2 _39031_ (.A1(_16967_),
    .A2(_16971_),
    .B1(_16972_),
    .Y(_16973_));
 sky130_fd_sc_hd__and3_2 _39032_ (.A(_16967_),
    .B(_16971_),
    .C(_16972_),
    .X(_16974_));
 sky130_fd_sc_hd__o22ai_2 _39033_ (.A1(_16916_),
    .A2(_16917_),
    .B1(_16973_),
    .B2(_16974_),
    .Y(_16975_));
 sky130_fd_sc_hd__nand2_2 _39034_ (.A(_16967_),
    .B(_16971_),
    .Y(_16976_));
 sky130_fd_sc_hd__a311oi_2 _39035_ (.A1(_16766_),
    .A2(_16767_),
    .A3(_16768_),
    .B1(_16784_),
    .C1(_16783_),
    .Y(_16977_));
 sky130_fd_sc_hd__nor2_2 _39036_ (.A(_16790_),
    .B(_16977_),
    .Y(_16978_));
 sky130_fd_sc_hd__nand2_2 _39037_ (.A(_16976_),
    .B(_16978_),
    .Y(_16979_));
 sky130_fd_sc_hd__nor2_2 _39038_ (.A(_16916_),
    .B(_16917_),
    .Y(_16980_));
 sky130_fd_sc_hd__nand3_2 _39039_ (.A(_16967_),
    .B(_16971_),
    .C(_16972_),
    .Y(_16981_));
 sky130_fd_sc_hd__nand3_2 _39040_ (.A(_16979_),
    .B(_16980_),
    .C(_16981_),
    .Y(_16982_));
 sky130_fd_sc_hd__o21ai_2 _39041_ (.A1(_16810_),
    .A2(_16789_),
    .B1(_16813_),
    .Y(_16983_));
 sky130_fd_sc_hd__a21oi_2 _39042_ (.A1(_16975_),
    .A2(_16982_),
    .B1(_16983_),
    .Y(_16984_));
 sky130_fd_sc_hd__nand2_2 _39043_ (.A(_16979_),
    .B(_16980_),
    .Y(_16985_));
 sky130_fd_sc_hd__o211a_2 _39044_ (.A1(_16974_),
    .A2(_16985_),
    .B1(_16983_),
    .C1(_16975_),
    .X(_16986_));
 sky130_fd_sc_hd__o22ai_2 _39045_ (.A1(_16903_),
    .A2(_16904_),
    .B1(_16984_),
    .B2(_16986_),
    .Y(_16987_));
 sky130_fd_sc_hd__a21o_2 _39046_ (.A1(_16975_),
    .A2(_16982_),
    .B1(_16983_),
    .X(_16988_));
 sky130_fd_sc_hd__nor2_2 _39047_ (.A(_16903_),
    .B(_16904_),
    .Y(_16989_));
 sky130_fd_sc_hd__nand3_2 _39048_ (.A(_16975_),
    .B(_16983_),
    .C(_16982_),
    .Y(_16990_));
 sky130_fd_sc_hd__nand3_2 _39049_ (.A(_16988_),
    .B(_16989_),
    .C(_16990_),
    .Y(_16991_));
 sky130_fd_sc_hd__o21ai_2 _39050_ (.A1(_16835_),
    .A2(_16817_),
    .B1(_16828_),
    .Y(_16992_));
 sky130_fd_sc_hd__a21oi_2 _39051_ (.A1(_16987_),
    .A2(_16991_),
    .B1(_16992_),
    .Y(_16993_));
 sky130_fd_sc_hd__a21oi_2 _39052_ (.A1(_16825_),
    .A2(_16826_),
    .B1(_16835_),
    .Y(_16994_));
 sky130_fd_sc_hd__o211a_2 _39053_ (.A1(_16820_),
    .A2(_16994_),
    .B1(_16991_),
    .C1(_16987_),
    .X(_16995_));
 sky130_fd_sc_hd__nand3_2 _39054_ (.A(_16740_),
    .B(_16083_),
    .C(_16735_),
    .Y(_16996_));
 sky130_fd_sc_hd__nand2_2 _39055_ (.A(_16996_),
    .B(_16093_),
    .Y(_16997_));
 sky130_fd_sc_hd__a21o_2 _39056_ (.A1(_16740_),
    .A2(_16735_),
    .B1(_16085_),
    .X(_16998_));
 sky130_fd_sc_hd__inv_2 _39057_ (.A(_16998_),
    .Y(_16999_));
 sky130_fd_sc_hd__nand2_2 _39058_ (.A(_16998_),
    .B(_16996_),
    .Y(_17000_));
 sky130_fd_sc_hd__nand2_2 _39059_ (.A(_17000_),
    .B(_16089_),
    .Y(_17001_));
 sky130_fd_sc_hd__o21ai_2 _39060_ (.A1(_16997_),
    .A2(_16999_),
    .B1(_17001_),
    .Y(_17002_));
 sky130_fd_sc_hd__o21ai_2 _39061_ (.A1(_16993_),
    .A2(_16995_),
    .B1(_17002_),
    .Y(_17003_));
 sky130_fd_sc_hd__nand2_2 _39062_ (.A(_16837_),
    .B(_16850_),
    .Y(_17004_));
 sky130_fd_sc_hd__nand2_2 _39063_ (.A(_17004_),
    .B(_16830_),
    .Y(_17005_));
 sky130_fd_sc_hd__a21o_2 _39064_ (.A1(_16987_),
    .A2(_16991_),
    .B1(_16992_),
    .X(_17006_));
 sky130_fd_sc_hd__nand3_2 _39065_ (.A(_16987_),
    .B(_16992_),
    .C(_16991_),
    .Y(_17007_));
 sky130_fd_sc_hd__nand3b_2 _39066_ (.A_N(_17002_),
    .B(_17006_),
    .C(_17007_),
    .Y(_17008_));
 sky130_fd_sc_hd__nand3_2 _39067_ (.A(_17003_),
    .B(_17005_),
    .C(_17008_),
    .Y(_17009_));
 sky130_fd_sc_hd__and2_2 _39068_ (.A(_17000_),
    .B(_16294_),
    .X(_17010_));
 sky130_fd_sc_hd__nor2_2 _39069_ (.A(_16844_),
    .B(_17000_),
    .Y(_17011_));
 sky130_fd_sc_hd__o22ai_2 _39070_ (.A1(_17010_),
    .A2(_17011_),
    .B1(_16993_),
    .B2(_16995_),
    .Y(_17012_));
 sky130_fd_sc_hd__a21boi_2 _39071_ (.A1(_16837_),
    .A2(_16850_),
    .B1_N(_16830_),
    .Y(_17013_));
 sky130_fd_sc_hd__nand3_2 _39072_ (.A(_17006_),
    .B(_17007_),
    .C(_17002_),
    .Y(_17014_));
 sky130_fd_sc_hd__nand3_2 _39073_ (.A(_17012_),
    .B(_17013_),
    .C(_17014_),
    .Y(_17015_));
 sky130_fd_sc_hd__nand2_2 _39074_ (.A(_16841_),
    .B(_16293_),
    .Y(_17016_));
 sky130_fd_sc_hd__nand2_2 _39075_ (.A(_17016_),
    .B(_16840_),
    .Y(_17017_));
 sky130_fd_sc_hd__nor2_2 _39076_ (.A(_13737_),
    .B(_17017_),
    .Y(_17018_));
 sky130_fd_sc_hd__inv_2 _39077_ (.A(_17017_),
    .Y(_17019_));
 sky130_fd_sc_hd__nor2_2 _39078_ (.A(_14823_),
    .B(_17019_),
    .Y(_17020_));
 sky130_fd_sc_hd__nor2_2 _39079_ (.A(_17018_),
    .B(_17020_),
    .Y(_17021_));
 sky130_fd_sc_hd__a21oi_2 _39080_ (.A1(_17009_),
    .A2(_17015_),
    .B1(_17021_),
    .Y(_17022_));
 sky130_fd_sc_hd__a21oi_2 _39081_ (.A1(_16857_),
    .A2(_16858_),
    .B1(_16854_),
    .Y(_17023_));
 sky130_fd_sc_hd__a31oi_2 _39082_ (.A1(_16854_),
    .A2(_16857_),
    .A3(_16858_),
    .B1(_16865_),
    .Y(_17024_));
 sky130_fd_sc_hd__nand3_2 _39083_ (.A(_17009_),
    .B(_17015_),
    .C(_17021_),
    .Y(_17025_));
 sky130_fd_sc_hd__o21ai_2 _39084_ (.A1(_17023_),
    .A2(_17024_),
    .B1(_17025_),
    .Y(_17026_));
 sky130_fd_sc_hd__nor2_2 _39085_ (.A(_16118_),
    .B(_17017_),
    .Y(_17027_));
 sky130_fd_sc_hd__nor2_2 _39086_ (.A(_16120_),
    .B(_17019_),
    .Y(_17028_));
 sky130_fd_sc_hd__o2bb2ai_2 _39087_ (.A1_N(_17015_),
    .A2_N(_17009_),
    .B1(_17027_),
    .B2(_17028_),
    .Y(_17029_));
 sky130_fd_sc_hd__a21oi_2 _39088_ (.A1(_16859_),
    .A2(_16871_),
    .B1(_17023_),
    .Y(_17030_));
 sky130_fd_sc_hd__nand3b_2 _39089_ (.A_N(_17021_),
    .B(_17009_),
    .C(_17015_),
    .Y(_17031_));
 sky130_fd_sc_hd__nand3_2 _39090_ (.A(_17029_),
    .B(_17030_),
    .C(_17031_),
    .Y(_17032_));
 sky130_fd_sc_hd__o211a_2 _39091_ (.A1(_17022_),
    .A2(_17026_),
    .B1(_16874_),
    .C1(_17032_),
    .X(_17033_));
 sky130_fd_sc_hd__o2bb2ai_2 _39092_ (.A1_N(_17015_),
    .A2_N(_17009_),
    .B1(_17020_),
    .B2(_17018_),
    .Y(_17034_));
 sky130_fd_sc_hd__o211ai_2 _39093_ (.A1(_17023_),
    .A2(_17024_),
    .B1(_17025_),
    .C1(_17034_),
    .Y(_17035_));
 sky130_fd_sc_hd__nand2_2 _39094_ (.A(_17035_),
    .B(_17032_),
    .Y(_17036_));
 sky130_fd_sc_hd__nor2_2 _39095_ (.A(_16869_),
    .B(_16870_),
    .Y(_17037_));
 sky130_fd_sc_hd__a21oi_2 _39096_ (.A1(_16867_),
    .A2(_16866_),
    .B1(_17037_),
    .Y(_17038_));
 sky130_fd_sc_hd__inv_2 _39097_ (.A(_16878_),
    .Y(_17039_));
 sky130_fd_sc_hd__a31oi_2 _39098_ (.A1(_17037_),
    .A2(_16867_),
    .A3(_16866_),
    .B1(_17039_),
    .Y(_17040_));
 sky130_fd_sc_hd__o2bb2ai_2 _39099_ (.A1_N(_16873_),
    .A2_N(_17036_),
    .B1(_17038_),
    .B2(_17040_),
    .Y(_17041_));
 sky130_fd_sc_hd__a2bb2oi_2 _39100_ (.A1_N(_15729_),
    .A2_N(_16863_),
    .B1(_17032_),
    .B2(_17035_),
    .Y(_17042_));
 sky130_fd_sc_hd__nor2_2 _39101_ (.A(_17038_),
    .B(_17040_),
    .Y(_17043_));
 sky130_fd_sc_hd__o21ai_2 _39102_ (.A1(_17042_),
    .A2(_17033_),
    .B1(_17043_),
    .Y(_17044_));
 sky130_fd_sc_hd__o21a_2 _39103_ (.A1(_17033_),
    .A2(_17041_),
    .B1(_17044_),
    .X(_17045_));
 sky130_fd_sc_hd__a21o_2 _39104_ (.A1(_16896_),
    .A2(_16887_),
    .B1(_17045_),
    .X(_17046_));
 sky130_fd_sc_hd__nand3_2 _39105_ (.A(_16896_),
    .B(_16887_),
    .C(_17045_),
    .Y(_17047_));
 sky130_fd_sc_hd__nand2_2 _39106_ (.A(_17046_),
    .B(_17047_),
    .Y(_02674_));
 sky130_fd_sc_hd__buf_1 _39107_ (.A(_14855_),
    .X(_17048_));
 sky130_fd_sc_hd__o41ai_2 _39108_ (.A1(_18184_),
    .A2(_17048_),
    .A3(_09226_),
    .A4(_19572_),
    .B1(_16930_),
    .Y(_17049_));
 sky130_fd_sc_hd__nor2_2 _39109_ (.A(_10152_),
    .B(_10523_),
    .Y(_17050_));
 sky130_fd_sc_hd__or4_2 _39110_ (.A(_09223_),
    .B(_13848_),
    .C(_14855_),
    .D(_15159_),
    .X(_17051_));
 sky130_fd_sc_hd__a22o_2 _39111_ (.A1(_19309_),
    .A2(_19566_),
    .B1(_10485_),
    .B2(_14350_),
    .X(_17052_));
 sky130_fd_sc_hd__nand2_2 _39112_ (.A(_17051_),
    .B(_17052_),
    .Y(_17053_));
 sky130_fd_sc_hd__or2_2 _39113_ (.A(_17050_),
    .B(_17053_),
    .X(_17054_));
 sky130_fd_sc_hd__nand2_2 _39114_ (.A(_17053_),
    .B(_17050_),
    .Y(_17055_));
 sky130_fd_sc_hd__nand3b_2 _39115_ (.A_N(_17049_),
    .B(_17054_),
    .C(_17055_),
    .Y(_17056_));
 sky130_fd_sc_hd__inv_2 _39116_ (.A(_17050_),
    .Y(_17057_));
 sky130_fd_sc_hd__or2_2 _39117_ (.A(_17057_),
    .B(_17053_),
    .X(_17058_));
 sky130_fd_sc_hd__nand2_2 _39118_ (.A(_17053_),
    .B(_17057_),
    .Y(_17059_));
 sky130_fd_sc_hd__nand3_2 _39119_ (.A(_17058_),
    .B(_17049_),
    .C(_17059_),
    .Y(_17060_));
 sky130_fd_sc_hd__nand2_2 _39120_ (.A(_15778_),
    .B(_19551_),
    .Y(_17061_));
 sky130_fd_sc_hd__a22o_2 _39121_ (.A1(_19317_),
    .A2(_09733_),
    .B1(_14042_),
    .B2(_19554_),
    .X(_17062_));
 sky130_fd_sc_hd__o21ai_2 _39122_ (.A1(_16003_),
    .A2(_15415_),
    .B1(_17062_),
    .Y(_17063_));
 sky130_fd_sc_hd__or2_2 _39123_ (.A(_17061_),
    .B(_17063_),
    .X(_17064_));
 sky130_fd_sc_hd__nand2_2 _39124_ (.A(_17063_),
    .B(_17061_),
    .Y(_17065_));
 sky130_fd_sc_hd__and2_2 _39125_ (.A(_17064_),
    .B(_17065_),
    .X(_17066_));
 sky130_fd_sc_hd__a21oi_2 _39126_ (.A1(_17056_),
    .A2(_17060_),
    .B1(_17066_),
    .Y(_17067_));
 sky130_fd_sc_hd__and3_2 _39127_ (.A(_17056_),
    .B(_17060_),
    .C(_17066_),
    .X(_17068_));
 sky130_fd_sc_hd__nand2_2 _39128_ (.A(_16942_),
    .B(_16931_),
    .Y(_17069_));
 sky130_fd_sc_hd__o21bai_2 _39129_ (.A1(_17067_),
    .A2(_17068_),
    .B1_N(_17069_),
    .Y(_17070_));
 sky130_fd_sc_hd__nand3_2 _39130_ (.A(_17056_),
    .B(_17060_),
    .C(_17066_),
    .Y(_17071_));
 sky130_fd_sc_hd__nand3b_2 _39131_ (.A_N(_17067_),
    .B(_17071_),
    .C(_17069_),
    .Y(_17072_));
 sky130_fd_sc_hd__inv_2 _39132_ (.A(_16953_),
    .Y(_17073_));
 sky130_fd_sc_hd__nor2_2 _39133_ (.A(_16951_),
    .B(_17073_),
    .Y(_17074_));
 sky130_fd_sc_hd__or2_2 _39134_ (.A(_16935_),
    .B(_16939_),
    .X(_17075_));
 sky130_fd_sc_hd__nand2_2 _39135_ (.A(_18157_),
    .B(_19334_),
    .Y(_17076_));
 sky130_fd_sc_hd__buf_1 _39136_ (.A(_17076_),
    .X(_17077_));
 sky130_fd_sc_hd__nand2_2 _39137_ (.A(_14569_),
    .B(_19545_),
    .Y(_17078_));
 sky130_fd_sc_hd__or3_2 _39138_ (.A(_17078_),
    .B(_13873_),
    .C(_10519_),
    .X(_17079_));
 sky130_fd_sc_hd__o21ai_2 _39139_ (.A1(_13873_),
    .A2(_10520_),
    .B1(_17078_),
    .Y(_17080_));
 sky130_fd_sc_hd__nand2_2 _39140_ (.A(_17079_),
    .B(_17080_),
    .Y(_17081_));
 sky130_fd_sc_hd__or2_2 _39141_ (.A(_17077_),
    .B(_17081_),
    .X(_17082_));
 sky130_fd_sc_hd__nand2_2 _39142_ (.A(_17081_),
    .B(_17077_),
    .Y(_17083_));
 sky130_fd_sc_hd__and2_2 _39143_ (.A(_17082_),
    .B(_17083_),
    .X(_17084_));
 sky130_fd_sc_hd__nor2_2 _39144_ (.A(_17075_),
    .B(_17084_),
    .Y(_17085_));
 sky130_fd_sc_hd__and3_2 _39145_ (.A(_17075_),
    .B(_17083_),
    .C(_17082_),
    .X(_17086_));
 sky130_fd_sc_hd__nor3_2 _39146_ (.A(_17074_),
    .B(_17085_),
    .C(_17086_),
    .Y(_17087_));
 sky130_fd_sc_hd__o21a_2 _39147_ (.A1(_17085_),
    .A2(_17086_),
    .B1(_17074_),
    .X(_17088_));
 sky130_fd_sc_hd__nor2_2 _39148_ (.A(_17087_),
    .B(_17088_),
    .Y(_17089_));
 sky130_fd_sc_hd__a21oi_2 _39149_ (.A1(_17070_),
    .A2(_17072_),
    .B1(_17089_),
    .Y(_17090_));
 sky130_fd_sc_hd__or2_2 _39150_ (.A(_17075_),
    .B(_17084_),
    .X(_17091_));
 sky130_fd_sc_hd__nand2_2 _39151_ (.A(_17084_),
    .B(_17075_),
    .Y(_17092_));
 sky130_fd_sc_hd__nand3b_2 _39152_ (.A_N(_17074_),
    .B(_17091_),
    .C(_17092_),
    .Y(_17093_));
 sky130_fd_sc_hd__o21ai_2 _39153_ (.A1(_17085_),
    .A2(_17086_),
    .B1(_17074_),
    .Y(_17094_));
 sky130_fd_sc_hd__and4_2 _39154_ (.A(_17070_),
    .B(_17072_),
    .C(_17093_),
    .D(_17094_),
    .X(_17095_));
 sky130_fd_sc_hd__nand2_2 _39155_ (.A(_16971_),
    .B(_16943_),
    .Y(_17096_));
 sky130_fd_sc_hd__o21bai_2 _39156_ (.A1(_17090_),
    .A2(_17095_),
    .B1_N(_17096_),
    .Y(_17097_));
 sky130_fd_sc_hd__a21o_2 _39157_ (.A1(_17070_),
    .A2(_17072_),
    .B1(_17089_),
    .X(_17098_));
 sky130_fd_sc_hd__nand3_2 _39158_ (.A(_17089_),
    .B(_17070_),
    .C(_17072_),
    .Y(_17099_));
 sky130_fd_sc_hd__nand3_2 _39159_ (.A(_17098_),
    .B(_17096_),
    .C(_17099_),
    .Y(_17100_));
 sky130_fd_sc_hd__nor2_2 _39160_ (.A(_16956_),
    .B(_16958_),
    .Y(_17101_));
 sky130_fd_sc_hd__nor2_2 _39161_ (.A(_17101_),
    .B(_16966_),
    .Y(_17102_));
 sky130_fd_sc_hd__and4_2 _39162_ (.A(_18158_),
    .B(_19338_),
    .C(_19341_),
    .D(_19344_),
    .X(_17103_));
 sky130_fd_sc_hd__nor2_2 _39163_ (.A(_16907_),
    .B(_16424_),
    .Y(_17104_));
 sky130_fd_sc_hd__or2_2 _39164_ (.A(_17103_),
    .B(_17104_),
    .X(_17105_));
 sky130_fd_sc_hd__buf_1 _39165_ (.A(_17105_),
    .X(_17106_));
 sky130_fd_sc_hd__nand2_2 _39166_ (.A(_16420_),
    .B(_17103_),
    .Y(_17107_));
 sky130_fd_sc_hd__and2_2 _39167_ (.A(_16425_),
    .B(_16907_),
    .X(_17108_));
 sky130_fd_sc_hd__a21o_2 _39168_ (.A1(_17106_),
    .A2(_17107_),
    .B1(_17108_),
    .X(_17109_));
 sky130_fd_sc_hd__nand2_2 _39169_ (.A(_17102_),
    .B(_17109_),
    .Y(_17110_));
 sky130_fd_sc_hd__a21oi_2 _39170_ (.A1(_17105_),
    .A2(_17107_),
    .B1(_17108_),
    .Y(_17111_));
 sky130_fd_sc_hd__o21ai_2 _39171_ (.A1(_17101_),
    .A2(_16966_),
    .B1(_17111_),
    .Y(_17112_));
 sky130_fd_sc_hd__nand2_2 _39172_ (.A(_17110_),
    .B(_17112_),
    .Y(_17113_));
 sky130_fd_sc_hd__nor2_2 _39173_ (.A(_16908_),
    .B(_16425_),
    .Y(_17114_));
 sky130_fd_sc_hd__nor2_2 _39174_ (.A(_17103_),
    .B(_17114_),
    .Y(_17115_));
 sky130_fd_sc_hd__nand2_2 _39175_ (.A(_17113_),
    .B(_17115_),
    .Y(_17116_));
 sky130_fd_sc_hd__inv_2 _39176_ (.A(_17115_),
    .Y(_17117_));
 sky130_fd_sc_hd__nand3_2 _39177_ (.A(_17110_),
    .B(_17117_),
    .C(_17112_),
    .Y(_17118_));
 sky130_fd_sc_hd__nand2_2 _39178_ (.A(_17116_),
    .B(_17118_),
    .Y(_17119_));
 sky130_fd_sc_hd__inv_2 _39179_ (.A(_17119_),
    .Y(_17120_));
 sky130_fd_sc_hd__a21oi_2 _39180_ (.A1(_17097_),
    .A2(_17100_),
    .B1(_17120_),
    .Y(_17121_));
 sky130_fd_sc_hd__and2_2 _39181_ (.A(_17113_),
    .B(_17117_),
    .X(_17122_));
 sky130_fd_sc_hd__nor2_2 _39182_ (.A(_17117_),
    .B(_17113_),
    .Y(_17123_));
 sky130_fd_sc_hd__o211a_2 _39183_ (.A1(_17122_),
    .A2(_17123_),
    .B1(_17100_),
    .C1(_17097_),
    .X(_17124_));
 sky130_fd_sc_hd__nand2_2 _39184_ (.A(_16985_),
    .B(_16981_),
    .Y(_17125_));
 sky130_fd_sc_hd__o21bai_2 _39185_ (.A1(_17121_),
    .A2(_17124_),
    .B1_N(_17125_),
    .Y(_17126_));
 sky130_fd_sc_hd__a21o_2 _39186_ (.A1(_17097_),
    .A2(_17100_),
    .B1(_17120_),
    .X(_17127_));
 sky130_fd_sc_hd__nand3_2 _39187_ (.A(_17120_),
    .B(_17097_),
    .C(_17100_),
    .Y(_17128_));
 sky130_fd_sc_hd__nand3_2 _39188_ (.A(_17127_),
    .B(_17128_),
    .C(_17125_),
    .Y(_17129_));
 sky130_fd_sc_hd__inv_2 _39189_ (.A(_16734_),
    .Y(_17130_));
 sky130_fd_sc_hd__a31o_2 _39190_ (.A1(_16909_),
    .A2(_16910_),
    .A3(_16912_),
    .B1(_16917_),
    .X(_17131_));
 sky130_fd_sc_hd__or2_2 _39191_ (.A(_17130_),
    .B(_17131_),
    .X(_17132_));
 sky130_fd_sc_hd__nand2_2 _39192_ (.A(_17131_),
    .B(_17130_),
    .Y(_17133_));
 sky130_fd_sc_hd__inv_2 _39193_ (.A(_16901_),
    .Y(_17134_));
 sky130_fd_sc_hd__buf_1 _39194_ (.A(_17134_),
    .X(_17135_));
 sky130_fd_sc_hd__a21oi_2 _39195_ (.A1(_17132_),
    .A2(_17133_),
    .B1(_17135_),
    .Y(_17136_));
 sky130_fd_sc_hd__nand3_2 _39196_ (.A(_17132_),
    .B(_17134_),
    .C(_17133_),
    .Y(_17137_));
 sky130_fd_sc_hd__nand2b_2 _39197_ (.A_N(_17136_),
    .B(_17137_),
    .Y(_17138_));
 sky130_fd_sc_hd__a21oi_2 _39198_ (.A1(_17126_),
    .A2(_17129_),
    .B1(_17138_),
    .Y(_17139_));
 sky130_fd_sc_hd__inv_2 _39199_ (.A(_17137_),
    .Y(_17140_));
 sky130_fd_sc_hd__o211a_2 _39200_ (.A1(_17136_),
    .A2(_17140_),
    .B1(_17129_),
    .C1(_17126_),
    .X(_17141_));
 sky130_fd_sc_hd__and2_2 _39201_ (.A(_16991_),
    .B(_16990_),
    .X(_17142_));
 sky130_fd_sc_hd__o21ai_2 _39202_ (.A1(_17139_),
    .A2(_17141_),
    .B1(_17142_),
    .Y(_17143_));
 sky130_fd_sc_hd__a21o_2 _39203_ (.A1(_17126_),
    .A2(_17129_),
    .B1(_17138_),
    .X(_17144_));
 sky130_fd_sc_hd__nand3_2 _39204_ (.A(_17138_),
    .B(_17126_),
    .C(_17129_),
    .Y(_17145_));
 sky130_fd_sc_hd__nand3b_2 _39205_ (.A_N(_17142_),
    .B(_17144_),
    .C(_17145_),
    .Y(_17146_));
 sky130_fd_sc_hd__buf_1 _39206_ (.A(_16089_),
    .X(_17147_));
 sky130_fd_sc_hd__a21bo_2 _39207_ (.A1(_16898_),
    .A2(_16901_),
    .B1_N(_16897_),
    .X(_17148_));
 sky130_fd_sc_hd__or2_2 _39208_ (.A(_16839_),
    .B(_17148_),
    .X(_17149_));
 sky130_fd_sc_hd__buf_1 _39209_ (.A(_16839_),
    .X(_17150_));
 sky130_fd_sc_hd__nand2_2 _39210_ (.A(_17148_),
    .B(_17150_),
    .Y(_17151_));
 sky130_fd_sc_hd__nand2_2 _39211_ (.A(_17149_),
    .B(_17151_),
    .Y(_17152_));
 sky130_fd_sc_hd__xor2_2 _39212_ (.A(_17147_),
    .B(_17152_),
    .X(_17153_));
 sky130_fd_sc_hd__a21o_2 _39213_ (.A1(_17143_),
    .A2(_17146_),
    .B1(_17153_),
    .X(_17154_));
 sky130_fd_sc_hd__o21ai_2 _39214_ (.A1(_17002_),
    .A2(_16993_),
    .B1(_17007_),
    .Y(_17155_));
 sky130_fd_sc_hd__nand3_2 _39215_ (.A(_17143_),
    .B(_17146_),
    .C(_17153_),
    .Y(_17156_));
 sky130_fd_sc_hd__nand3_2 _39216_ (.A(_17154_),
    .B(_17155_),
    .C(_17156_),
    .Y(_17157_));
 sky130_fd_sc_hd__a21oi_2 _39217_ (.A1(_17143_),
    .A2(_17146_),
    .B1(_17153_),
    .Y(_17158_));
 sky130_fd_sc_hd__and3_2 _39218_ (.A(_17143_),
    .B(_17146_),
    .C(_17153_),
    .X(_17159_));
 sky130_fd_sc_hd__o21bai_2 _39219_ (.A1(_17158_),
    .A2(_17159_),
    .B1_N(_17155_),
    .Y(_17160_));
 sky130_fd_sc_hd__nand2_2 _39220_ (.A(_16997_),
    .B(_16998_),
    .Y(_17161_));
 sky130_fd_sc_hd__inv_2 _39221_ (.A(_17161_),
    .Y(_17162_));
 sky130_fd_sc_hd__nor2_2 _39222_ (.A(_15320_),
    .B(_17162_),
    .Y(_17163_));
 sky130_fd_sc_hd__buf_1 _39223_ (.A(_15109_),
    .X(_17164_));
 sky130_fd_sc_hd__buf_1 _39224_ (.A(_17164_),
    .X(_17165_));
 sky130_fd_sc_hd__nor2_2 _39225_ (.A(_17165_),
    .B(_17161_),
    .Y(_17166_));
 sky130_fd_sc_hd__o2bb2ai_2 _39226_ (.A1_N(_17157_),
    .A2_N(_17160_),
    .B1(_17163_),
    .B2(_17166_),
    .Y(_17167_));
 sky130_fd_sc_hd__nand2_2 _39227_ (.A(_17015_),
    .B(_17021_),
    .Y(_17168_));
 sky130_fd_sc_hd__nand2_2 _39228_ (.A(_17168_),
    .B(_17009_),
    .Y(_17169_));
 sky130_fd_sc_hd__nor2_2 _39229_ (.A(_16118_),
    .B(_17161_),
    .Y(_17170_));
 sky130_fd_sc_hd__nor2_2 _39230_ (.A(_15109_),
    .B(_17162_),
    .Y(_17171_));
 sky130_fd_sc_hd__nor2_2 _39231_ (.A(_17170_),
    .B(_17171_),
    .Y(_17172_));
 sky130_fd_sc_hd__inv_2 _39232_ (.A(_17172_),
    .Y(_17173_));
 sky130_fd_sc_hd__nand3_2 _39233_ (.A(_17160_),
    .B(_17157_),
    .C(_17173_),
    .Y(_17174_));
 sky130_fd_sc_hd__nand3_2 _39234_ (.A(_17167_),
    .B(_17169_),
    .C(_17174_),
    .Y(_17175_));
 sky130_fd_sc_hd__o2bb2ai_2 _39235_ (.A1_N(_17157_),
    .A2_N(_17160_),
    .B1(_17170_),
    .B2(_17171_),
    .Y(_17176_));
 sky130_fd_sc_hd__inv_2 _39236_ (.A(_17169_),
    .Y(_17177_));
 sky130_fd_sc_hd__nand3_2 _39237_ (.A(_17160_),
    .B(_17157_),
    .C(_17172_),
    .Y(_17178_));
 sky130_fd_sc_hd__nand3_2 _39238_ (.A(_17176_),
    .B(_17177_),
    .C(_17178_),
    .Y(_17179_));
 sky130_fd_sc_hd__buf_1 _39239_ (.A(_15320_),
    .X(_17180_));
 sky130_fd_sc_hd__o2bb2ai_2 _39240_ (.A1_N(_17175_),
    .A2_N(_17179_),
    .B1(_17180_),
    .B2(_17019_),
    .Y(_17181_));
 sky130_fd_sc_hd__nand3_2 _39241_ (.A(_17175_),
    .B(_17179_),
    .C(_17020_),
    .Y(_17182_));
 sky130_fd_sc_hd__nand3_2 _39242_ (.A(_17035_),
    .B(_17032_),
    .C(_16874_),
    .Y(_17183_));
 sky130_fd_sc_hd__nand2_2 _39243_ (.A(_17183_),
    .B(_17035_),
    .Y(_17184_));
 sky130_fd_sc_hd__a21oi_2 _39244_ (.A1(_17181_),
    .A2(_17182_),
    .B1(_17184_),
    .Y(_17185_));
 sky130_fd_sc_hd__and3_2 _39245_ (.A(_17181_),
    .B(_17184_),
    .C(_17182_),
    .X(_17186_));
 sky130_fd_sc_hd__nor2_2 _39246_ (.A(_17185_),
    .B(_17186_),
    .Y(_17187_));
 sky130_fd_sc_hd__o2111a_2 _39247_ (.A1(_17033_),
    .A2(_17041_),
    .B1(_16887_),
    .C1(_17044_),
    .D1(_16884_),
    .X(_17188_));
 sky130_fd_sc_hd__nand2_2 _39248_ (.A(_16890_),
    .B(_17188_),
    .Y(_17189_));
 sky130_fd_sc_hd__nor2_2 _39249_ (.A(_16521_),
    .B(_17189_),
    .Y(_17190_));
 sky130_fd_sc_hd__o2111ai_2 _39250_ (.A1(_17033_),
    .A2(_17041_),
    .B1(_16887_),
    .C1(_17044_),
    .D1(_16884_),
    .Y(_17191_));
 sky130_fd_sc_hd__o2bb2ai_2 _39251_ (.A1_N(_17035_),
    .A2_N(_17032_),
    .B1(_17180_),
    .B2(_16863_),
    .Y(_17192_));
 sky130_fd_sc_hd__nand2_2 _39252_ (.A(_16868_),
    .B(_16878_),
    .Y(_17193_));
 sky130_fd_sc_hd__nand2_2 _39253_ (.A(_17193_),
    .B(_16877_),
    .Y(_17194_));
 sky130_fd_sc_hd__a21oi_2 _39254_ (.A1(_17192_),
    .A2(_17183_),
    .B1(_17194_),
    .Y(_17195_));
 sky130_fd_sc_hd__o22a_2 _39255_ (.A1(_17033_),
    .A2(_17041_),
    .B1(_16887_),
    .B2(_17195_),
    .X(_17196_));
 sky130_fd_sc_hd__o21ai_2 _39256_ (.A1(_16893_),
    .A2(_17191_),
    .B1(_17196_),
    .Y(_17197_));
 sky130_fd_sc_hd__o21bai_2 _39257_ (.A1(_17189_),
    .A2(_16533_),
    .B1_N(_17197_),
    .Y(_17198_));
 sky130_fd_sc_hd__a21o_2 _39258_ (.A1(_15747_),
    .A2(_17190_),
    .B1(_17198_),
    .X(_17199_));
 sky130_fd_sc_hd__or2_2 _39259_ (.A(_17187_),
    .B(_17199_),
    .X(_17200_));
 sky130_fd_sc_hd__nand2_2 _39260_ (.A(_17199_),
    .B(_17187_),
    .Y(_17201_));
 sky130_fd_sc_hd__and2_2 _39261_ (.A(_17200_),
    .B(_17201_),
    .X(_02675_));
 sky130_fd_sc_hd__a21oi_2 _39262_ (.A1(_17154_),
    .A2(_17156_),
    .B1(_17155_),
    .Y(_17202_));
 sky130_fd_sc_hd__o21ai_2 _39263_ (.A1(_17172_),
    .A2(_17202_),
    .B1(_17157_),
    .Y(_17203_));
 sky130_fd_sc_hd__nand2_2 _39264_ (.A(_17143_),
    .B(_17153_),
    .Y(_17204_));
 sky130_fd_sc_hd__nand2_2 _39265_ (.A(_17204_),
    .B(_17146_),
    .Y(_17205_));
 sky130_fd_sc_hd__nand2_2 _39266_ (.A(_17099_),
    .B(_17072_),
    .Y(_17206_));
 sky130_fd_sc_hd__nand2_2 _39267_ (.A(_17071_),
    .B(_17060_),
    .Y(_17207_));
 sky130_fd_sc_hd__nor2_2 _39268_ (.A(_10152_),
    .B(_14939_),
    .Y(_17208_));
 sky130_fd_sc_hd__or4_2 _39269_ (.A(_19566_),
    .B(_18183_),
    .C(_14353_),
    .D(_10514_),
    .X(_17209_));
 sky130_fd_sc_hd__a22o_2 _39270_ (.A1(_19309_),
    .A2(_19563_),
    .B1(_15159_),
    .B2(_11123_),
    .X(_17210_));
 sky130_fd_sc_hd__nand2_2 _39271_ (.A(_17209_),
    .B(_17210_),
    .Y(_17211_));
 sky130_fd_sc_hd__or2_2 _39272_ (.A(_17208_),
    .B(_17211_),
    .X(_17212_));
 sky130_fd_sc_hd__nand2_2 _39273_ (.A(_17211_),
    .B(_17208_),
    .Y(_17213_));
 sky130_fd_sc_hd__nand2_2 _39274_ (.A(_17212_),
    .B(_17213_),
    .Y(_17214_));
 sky130_fd_sc_hd__o21ai_2 _39275_ (.A1(_17057_),
    .A2(_17053_),
    .B1(_17051_),
    .Y(_17215_));
 sky130_fd_sc_hd__nand2_2 _39276_ (.A(_17214_),
    .B(_17215_),
    .Y(_17216_));
 sky130_fd_sc_hd__nand3b_2 _39277_ (.A_N(_17215_),
    .B(_17212_),
    .C(_17213_),
    .Y(_17217_));
 sky130_fd_sc_hd__nand2_2 _39278_ (.A(_19325_),
    .B(_19547_),
    .Y(_17218_));
 sky130_fd_sc_hd__or2_2 _39279_ (.A(_10705_),
    .B(_15656_),
    .X(_17219_));
 sky130_fd_sc_hd__a22o_2 _39280_ (.A1(_19317_),
    .A2(_19554_),
    .B1(_19321_),
    .B2(_19550_),
    .X(_17220_));
 sky130_fd_sc_hd__nand2_2 _39281_ (.A(_17219_),
    .B(_17220_),
    .Y(_17221_));
 sky130_fd_sc_hd__or2_2 _39282_ (.A(_17218_),
    .B(_17221_),
    .X(_17222_));
 sky130_fd_sc_hd__nand2_2 _39283_ (.A(_17221_),
    .B(_17218_),
    .Y(_17223_));
 sky130_fd_sc_hd__nand2_2 _39284_ (.A(_17222_),
    .B(_17223_),
    .Y(_17224_));
 sky130_fd_sc_hd__a21o_2 _39285_ (.A1(_17216_),
    .A2(_17217_),
    .B1(_17224_),
    .X(_17225_));
 sky130_fd_sc_hd__nand3_2 _39286_ (.A(_17216_),
    .B(_17217_),
    .C(_17224_),
    .Y(_17226_));
 sky130_fd_sc_hd__nand3b_2 _39287_ (.A_N(_17207_),
    .B(_17225_),
    .C(_17226_),
    .Y(_17227_));
 sky130_fd_sc_hd__inv_2 _39288_ (.A(_17224_),
    .Y(_17228_));
 sky130_fd_sc_hd__a21o_2 _39289_ (.A1(_17216_),
    .A2(_17217_),
    .B1(_17228_),
    .X(_17229_));
 sky130_fd_sc_hd__nand3_2 _39290_ (.A(_17216_),
    .B(_17217_),
    .C(_17228_),
    .Y(_17230_));
 sky130_fd_sc_hd__nand3_2 _39291_ (.A(_17229_),
    .B(_17207_),
    .C(_17230_),
    .Y(_17231_));
 sky130_fd_sc_hd__nand2_2 _39292_ (.A(_17227_),
    .B(_17231_),
    .Y(_17232_));
 sky130_fd_sc_hd__o21ai_2 _39293_ (.A1(_16003_),
    .A2(_15415_),
    .B1(_17064_),
    .Y(_17233_));
 sky130_fd_sc_hd__nand2_2 _39294_ (.A(_18156_),
    .B(_19331_),
    .Y(_17234_));
 sky130_fd_sc_hd__or3_2 _39295_ (.A(_17234_),
    .B(_14571_),
    .C(_10519_),
    .X(_17235_));
 sky130_fd_sc_hd__o21ai_2 _39296_ (.A1(_14571_),
    .A2(_10520_),
    .B1(_17234_),
    .Y(_17236_));
 sky130_fd_sc_hd__nand2_2 _39297_ (.A(_17235_),
    .B(_17236_),
    .Y(_17237_));
 sky130_fd_sc_hd__nor2_2 _39298_ (.A(_17077_),
    .B(_17237_),
    .Y(_17238_));
 sky130_fd_sc_hd__and2_2 _39299_ (.A(_17237_),
    .B(_17077_),
    .X(_17239_));
 sky130_fd_sc_hd__nor2_2 _39300_ (.A(_17238_),
    .B(_17239_),
    .Y(_17240_));
 sky130_fd_sc_hd__nor2_2 _39301_ (.A(_17233_),
    .B(_17240_),
    .Y(_17241_));
 sky130_fd_sc_hd__and2_2 _39302_ (.A(_17240_),
    .B(_17233_),
    .X(_17242_));
 sky130_fd_sc_hd__nor2_2 _39303_ (.A(_17241_),
    .B(_17242_),
    .Y(_17243_));
 sky130_fd_sc_hd__nand2_2 _39304_ (.A(_17082_),
    .B(_17079_),
    .Y(_17244_));
 sky130_fd_sc_hd__nand2_2 _39305_ (.A(_17243_),
    .B(_17244_),
    .Y(_17245_));
 sky130_fd_sc_hd__inv_2 _39306_ (.A(_17244_),
    .Y(_17246_));
 sky130_fd_sc_hd__o21ai_2 _39307_ (.A1(_17241_),
    .A2(_17242_),
    .B1(_17246_),
    .Y(_17247_));
 sky130_fd_sc_hd__nand2_2 _39308_ (.A(_17245_),
    .B(_17247_),
    .Y(_17248_));
 sky130_fd_sc_hd__nand2_2 _39309_ (.A(_17232_),
    .B(_17248_),
    .Y(_17249_));
 sky130_fd_sc_hd__inv_2 _39310_ (.A(_17248_),
    .Y(_17250_));
 sky130_fd_sc_hd__nand3_2 _39311_ (.A(_17250_),
    .B(_17227_),
    .C(_17231_),
    .Y(_17251_));
 sky130_fd_sc_hd__nand3_2 _39312_ (.A(_17206_),
    .B(_17249_),
    .C(_17251_),
    .Y(_17252_));
 sky130_fd_sc_hd__a22oi_2 _39313_ (.A1(_17247_),
    .A2(_17245_),
    .B1(_17227_),
    .B2(_17231_),
    .Y(_17253_));
 sky130_fd_sc_hd__nor2_2 _39314_ (.A(_17246_),
    .B(_17243_),
    .Y(_17254_));
 sky130_fd_sc_hd__and2_2 _39315_ (.A(_17243_),
    .B(_17246_),
    .X(_17255_));
 sky130_fd_sc_hd__o211a_2 _39316_ (.A1(_17254_),
    .A2(_17255_),
    .B1(_17231_),
    .C1(_17227_),
    .X(_17256_));
 sky130_fd_sc_hd__a21boi_2 _39317_ (.A1(_17089_),
    .A2(_17070_),
    .B1_N(_17072_),
    .Y(_17257_));
 sky130_fd_sc_hd__o21ai_2 _39318_ (.A1(_17253_),
    .A2(_17256_),
    .B1(_17257_),
    .Y(_17258_));
 sky130_fd_sc_hd__o21ai_2 _39319_ (.A1(_17086_),
    .A2(_17087_),
    .B1(_17111_),
    .Y(_17259_));
 sky130_fd_sc_hd__nand3_2 _39320_ (.A(_17093_),
    .B(_17092_),
    .C(_17109_),
    .Y(_17260_));
 sky130_fd_sc_hd__inv_2 _39321_ (.A(_17106_),
    .Y(_17261_));
 sky130_fd_sc_hd__a21o_2 _39322_ (.A1(_17259_),
    .A2(_17260_),
    .B1(_17261_),
    .X(_17262_));
 sky130_fd_sc_hd__buf_1 _39323_ (.A(_17261_),
    .X(_17263_));
 sky130_fd_sc_hd__nand3_2 _39324_ (.A(_17259_),
    .B(_17263_),
    .C(_17260_),
    .Y(_17264_));
 sky130_fd_sc_hd__nand2_2 _39325_ (.A(_17262_),
    .B(_17264_),
    .Y(_17265_));
 sky130_fd_sc_hd__a21oi_2 _39326_ (.A1(_17252_),
    .A2(_17258_),
    .B1(_17265_),
    .Y(_17266_));
 sky130_fd_sc_hd__and3_2 _39327_ (.A(_17252_),
    .B(_17258_),
    .C(_17265_),
    .X(_17267_));
 sky130_fd_sc_hd__a21oi_2 _39328_ (.A1(_17098_),
    .A2(_17099_),
    .B1(_17096_),
    .Y(_17268_));
 sky130_fd_sc_hd__o21ai_2 _39329_ (.A1(_17119_),
    .A2(_17268_),
    .B1(_17100_),
    .Y(_17269_));
 sky130_fd_sc_hd__o21bai_2 _39330_ (.A1(_17266_),
    .A2(_17267_),
    .B1_N(_17269_),
    .Y(_17270_));
 sky130_fd_sc_hd__a21o_2 _39331_ (.A1(_17252_),
    .A2(_17258_),
    .B1(_17265_),
    .X(_17271_));
 sky130_fd_sc_hd__nand3_2 _39332_ (.A(_17252_),
    .B(_17258_),
    .C(_17265_),
    .Y(_17272_));
 sky130_fd_sc_hd__nand3_2 _39333_ (.A(_17271_),
    .B(_17269_),
    .C(_17272_),
    .Y(_17273_));
 sky130_fd_sc_hd__nand2_2 _39334_ (.A(_17118_),
    .B(_17112_),
    .Y(_17274_));
 sky130_fd_sc_hd__nand2_2 _39335_ (.A(_17274_),
    .B(_17130_),
    .Y(_17275_));
 sky130_fd_sc_hd__nand3_2 _39336_ (.A(_17118_),
    .B(_16736_),
    .C(_17112_),
    .Y(_17276_));
 sky130_fd_sc_hd__nand2_2 _39337_ (.A(_17275_),
    .B(_17276_),
    .Y(_17277_));
 sky130_fd_sc_hd__nand2_2 _39338_ (.A(_17277_),
    .B(_16902_),
    .Y(_17278_));
 sky130_fd_sc_hd__nand3_2 _39339_ (.A(_17275_),
    .B(_17134_),
    .C(_17276_),
    .Y(_17279_));
 sky130_fd_sc_hd__nand2_2 _39340_ (.A(_17278_),
    .B(_17279_),
    .Y(_17280_));
 sky130_fd_sc_hd__inv_2 _39341_ (.A(_17280_),
    .Y(_17281_));
 sky130_fd_sc_hd__a21o_2 _39342_ (.A1(_17270_),
    .A2(_17273_),
    .B1(_17281_),
    .X(_17282_));
 sky130_fd_sc_hd__a21boi_2 _39343_ (.A1(_17138_),
    .A2(_17126_),
    .B1_N(_17129_),
    .Y(_17283_));
 sky130_fd_sc_hd__nand3_2 _39344_ (.A(_17270_),
    .B(_17273_),
    .C(_17281_),
    .Y(_17284_));
 sky130_fd_sc_hd__nand3_2 _39345_ (.A(_17282_),
    .B(_17283_),
    .C(_17284_),
    .Y(_17285_));
 sky130_fd_sc_hd__buf_1 _39346_ (.A(_16902_),
    .X(_17286_));
 sky130_fd_sc_hd__inv_2 _39347_ (.A(_17277_),
    .Y(_17287_));
 sky130_fd_sc_hd__nor2_2 _39348_ (.A(_17286_),
    .B(_17287_),
    .Y(_17288_));
 sky130_fd_sc_hd__nor2_2 _39349_ (.A(_17135_),
    .B(_17277_),
    .Y(_17289_));
 sky130_fd_sc_hd__o2bb2ai_2 _39350_ (.A1_N(_17273_),
    .A2_N(_17270_),
    .B1(_17288_),
    .B2(_17289_),
    .Y(_17290_));
 sky130_fd_sc_hd__nor2_2 _39351_ (.A(_17136_),
    .B(_17140_),
    .Y(_17291_));
 sky130_fd_sc_hd__a21oi_2 _39352_ (.A1(_17127_),
    .A2(_17128_),
    .B1(_17125_),
    .Y(_17292_));
 sky130_fd_sc_hd__o21ai_2 _39353_ (.A1(_17291_),
    .A2(_17292_),
    .B1(_17129_),
    .Y(_17293_));
 sky130_fd_sc_hd__nand3_2 _39354_ (.A(_17270_),
    .B(_17273_),
    .C(_17280_),
    .Y(_17294_));
 sky130_fd_sc_hd__nand3_2 _39355_ (.A(_17290_),
    .B(_17293_),
    .C(_17294_),
    .Y(_17295_));
 sky130_fd_sc_hd__nand2_2 _39356_ (.A(_17285_),
    .B(_17295_),
    .Y(_17296_));
 sky130_fd_sc_hd__nand2_2 _39357_ (.A(_17132_),
    .B(_16902_),
    .Y(_17297_));
 sky130_fd_sc_hd__a21o_2 _39358_ (.A1(_17297_),
    .A2(_17133_),
    .B1(_16083_),
    .X(_17298_));
 sky130_fd_sc_hd__nand3_2 _39359_ (.A(_17297_),
    .B(_16083_),
    .C(_17133_),
    .Y(_17299_));
 sky130_fd_sc_hd__nand2_2 _39360_ (.A(_17299_),
    .B(_16294_),
    .Y(_17300_));
 sky130_fd_sc_hd__inv_2 _39361_ (.A(_17300_),
    .Y(_17301_));
 sky130_fd_sc_hd__a21oi_2 _39362_ (.A1(_17298_),
    .A2(_17299_),
    .B1(_16844_),
    .Y(_17302_));
 sky130_fd_sc_hd__a21o_2 _39363_ (.A1(_17298_),
    .A2(_17301_),
    .B1(_17302_),
    .X(_17303_));
 sky130_fd_sc_hd__nand2_2 _39364_ (.A(_17296_),
    .B(_17303_),
    .Y(_17304_));
 sky130_fd_sc_hd__a21oi_2 _39365_ (.A1(_17301_),
    .A2(_17298_),
    .B1(_17302_),
    .Y(_17305_));
 sky130_fd_sc_hd__nand3_2 _39366_ (.A(_17285_),
    .B(_17295_),
    .C(_17305_),
    .Y(_17306_));
 sky130_fd_sc_hd__nand3_2 _39367_ (.A(_17205_),
    .B(_17304_),
    .C(_17306_),
    .Y(_17307_));
 sky130_fd_sc_hd__a21boi_2 _39368_ (.A1(_17143_),
    .A2(_17153_),
    .B1_N(_17146_),
    .Y(_17308_));
 sky130_fd_sc_hd__nand2_2 _39369_ (.A(_17296_),
    .B(_17305_),
    .Y(_17309_));
 sky130_fd_sc_hd__nand3_2 _39370_ (.A(_17285_),
    .B(_17295_),
    .C(_17303_),
    .Y(_17310_));
 sky130_fd_sc_hd__nand3_2 _39371_ (.A(_17308_),
    .B(_17309_),
    .C(_17310_),
    .Y(_17311_));
 sky130_fd_sc_hd__inv_2 _39372_ (.A(_17151_),
    .Y(_17312_));
 sky130_fd_sc_hd__and2_2 _39373_ (.A(_17149_),
    .B(_16294_),
    .X(_17313_));
 sky130_fd_sc_hd__nor2_2 _39374_ (.A(_17312_),
    .B(_17313_),
    .Y(_17314_));
 sky130_fd_sc_hd__nor2_2 _39375_ (.A(_14018_),
    .B(_17314_),
    .Y(_17315_));
 sky130_fd_sc_hd__inv_2 _39376_ (.A(_17315_),
    .Y(_17316_));
 sky130_fd_sc_hd__nand2_2 _39377_ (.A(_17314_),
    .B(_14019_),
    .Y(_17317_));
 sky130_fd_sc_hd__and2_2 _39378_ (.A(_17316_),
    .B(_17317_),
    .X(_17318_));
 sky130_fd_sc_hd__a21o_2 _39379_ (.A1(_17307_),
    .A2(_17311_),
    .B1(_17318_),
    .X(_17319_));
 sky130_fd_sc_hd__nand2_2 _39380_ (.A(_17316_),
    .B(_17317_),
    .Y(_17320_));
 sky130_fd_sc_hd__a31oi_2 _39381_ (.A1(_17308_),
    .A2(_17309_),
    .A3(_17310_),
    .B1(_17320_),
    .Y(_17321_));
 sky130_fd_sc_hd__nand2_2 _39382_ (.A(_17321_),
    .B(_17307_),
    .Y(_17322_));
 sky130_fd_sc_hd__nand3_2 _39383_ (.A(_17203_),
    .B(_17319_),
    .C(_17322_),
    .Y(_17323_));
 sky130_fd_sc_hd__a21boi_2 _39384_ (.A1(_17160_),
    .A2(_17173_),
    .B1_N(_17157_),
    .Y(_17324_));
 sky130_fd_sc_hd__a21o_2 _39385_ (.A1(_17307_),
    .A2(_17311_),
    .B1(_17320_),
    .X(_17325_));
 sky130_fd_sc_hd__nand3_2 _39386_ (.A(_17307_),
    .B(_17311_),
    .C(_17320_),
    .Y(_17326_));
 sky130_fd_sc_hd__nand3_2 _39387_ (.A(_17324_),
    .B(_17325_),
    .C(_17326_),
    .Y(_17327_));
 sky130_fd_sc_hd__o2bb2ai_2 _39388_ (.A1_N(_17323_),
    .A2_N(_17327_),
    .B1(_17180_),
    .B2(_17162_),
    .Y(_17328_));
 sky130_fd_sc_hd__nand3_2 _39389_ (.A(_17327_),
    .B(_17323_),
    .C(_17163_),
    .Y(_17329_));
 sky130_fd_sc_hd__nand2_2 _39390_ (.A(_17179_),
    .B(_17020_),
    .Y(_17330_));
 sky130_fd_sc_hd__nand2_2 _39391_ (.A(_17330_),
    .B(_17175_),
    .Y(_17331_));
 sky130_fd_sc_hd__a21oi_2 _39392_ (.A1(_17328_),
    .A2(_17329_),
    .B1(_17331_),
    .Y(_17332_));
 sky130_fd_sc_hd__and3_2 _39393_ (.A(_17331_),
    .B(_17328_),
    .C(_17329_),
    .X(_17333_));
 sky130_fd_sc_hd__nor2_2 _39394_ (.A(_17332_),
    .B(_17333_),
    .Y(_17334_));
 sky130_fd_sc_hd__nand3_2 _39395_ (.A(_17181_),
    .B(_17184_),
    .C(_17182_),
    .Y(_17335_));
 sky130_fd_sc_hd__nand2_2 _39396_ (.A(_17201_),
    .B(_17335_),
    .Y(_17336_));
 sky130_fd_sc_hd__xor2_2 _39397_ (.A(_17334_),
    .B(_17336_),
    .X(_02676_));
 sky130_fd_sc_hd__a21oi_2 _39398_ (.A1(_17309_),
    .A2(_17310_),
    .B1(_17308_),
    .Y(_17337_));
 sky130_fd_sc_hd__inv_2 _39399_ (.A(_17242_),
    .Y(_17338_));
 sky130_fd_sc_hd__a21o_2 _39400_ (.A1(_17245_),
    .A2(_17338_),
    .B1(_17109_),
    .X(_17339_));
 sky130_fd_sc_hd__nand3_2 _39401_ (.A(_17109_),
    .B(_17245_),
    .C(_17338_),
    .Y(_17340_));
 sky130_fd_sc_hd__nand2_2 _39402_ (.A(_17339_),
    .B(_17340_),
    .Y(_17341_));
 sky130_fd_sc_hd__nand2_2 _39403_ (.A(_17341_),
    .B(_17106_),
    .Y(_17342_));
 sky130_fd_sc_hd__inv_2 _39404_ (.A(_17342_),
    .Y(_17343_));
 sky130_fd_sc_hd__nand3_2 _39405_ (.A(_17339_),
    .B(_17263_),
    .C(_17340_),
    .Y(_17344_));
 sky130_fd_sc_hd__inv_2 _39406_ (.A(_17344_),
    .Y(_17345_));
 sky130_fd_sc_hd__nand2_2 _39407_ (.A(_17230_),
    .B(_17216_),
    .Y(_17346_));
 sky130_fd_sc_hd__a21bo_2 _39408_ (.A1(_17208_),
    .A2(_17210_),
    .B1_N(_17209_),
    .X(_17347_));
 sky130_fd_sc_hd__nor2_2 _39409_ (.A(_10152_),
    .B(_10543_),
    .Y(_17348_));
 sky130_fd_sc_hd__or4_2 _39410_ (.A(_19563_),
    .B(_18183_),
    .C(_17048_),
    .D(_14939_),
    .X(_17349_));
 sky130_fd_sc_hd__a22o_2 _39411_ (.A1(_19309_),
    .A2(_19560_),
    .B1(_10523_),
    .B2(_11123_),
    .X(_17350_));
 sky130_fd_sc_hd__nand2_2 _39412_ (.A(_17349_),
    .B(_17350_),
    .Y(_17351_));
 sky130_fd_sc_hd__or2_2 _39413_ (.A(_17348_),
    .B(_17351_),
    .X(_17352_));
 sky130_fd_sc_hd__nand2_2 _39414_ (.A(_17351_),
    .B(_17348_),
    .Y(_17353_));
 sky130_fd_sc_hd__nand3b_2 _39415_ (.A_N(_17347_),
    .B(_17352_),
    .C(_17353_),
    .Y(_17354_));
 sky130_fd_sc_hd__inv_2 _39416_ (.A(_17348_),
    .Y(_17355_));
 sky130_fd_sc_hd__or2_2 _39417_ (.A(_17355_),
    .B(_17351_),
    .X(_17356_));
 sky130_fd_sc_hd__nand2_2 _39418_ (.A(_17351_),
    .B(_17355_),
    .Y(_17357_));
 sky130_fd_sc_hd__nand3_2 _39419_ (.A(_17356_),
    .B(_17347_),
    .C(_17357_),
    .Y(_17358_));
 sky130_fd_sc_hd__nand2_2 _39420_ (.A(_19325_),
    .B(_19543_),
    .Y(_17359_));
 sky130_fd_sc_hd__a22o_2 _39421_ (.A1(_19318_),
    .A2(_19550_),
    .B1(_19321_),
    .B2(_19546_),
    .X(_17360_));
 sky130_fd_sc_hd__o21ai_2 _39422_ (.A1(_16003_),
    .A2(_10539_),
    .B1(_17360_),
    .Y(_17361_));
 sky130_fd_sc_hd__or2_2 _39423_ (.A(_17359_),
    .B(_17361_),
    .X(_17362_));
 sky130_fd_sc_hd__nand2_2 _39424_ (.A(_17361_),
    .B(_17359_),
    .Y(_17363_));
 sky130_fd_sc_hd__and2_2 _39425_ (.A(_17362_),
    .B(_17363_),
    .X(_17364_));
 sky130_fd_sc_hd__a21o_2 _39426_ (.A1(_17354_),
    .A2(_17358_),
    .B1(_17364_),
    .X(_17365_));
 sky130_fd_sc_hd__nand3_2 _39427_ (.A(_17354_),
    .B(_17358_),
    .C(_17364_),
    .Y(_17366_));
 sky130_fd_sc_hd__nand3_2 _39428_ (.A(_17346_),
    .B(_17365_),
    .C(_17366_),
    .Y(_17367_));
 sky130_fd_sc_hd__a21boi_2 _39429_ (.A1(_17217_),
    .A2(_17228_),
    .B1_N(_17216_),
    .Y(_17368_));
 sky130_fd_sc_hd__nand3b_2 _39430_ (.A_N(_17364_),
    .B(_17354_),
    .C(_17358_),
    .Y(_17369_));
 sky130_fd_sc_hd__a21bo_2 _39431_ (.A1(_17354_),
    .A2(_17358_),
    .B1_N(_17364_),
    .X(_17370_));
 sky130_fd_sc_hd__nand3_2 _39432_ (.A(_17368_),
    .B(_17369_),
    .C(_17370_),
    .Y(_17371_));
 sky130_fd_sc_hd__o21a_2 _39433_ (.A1(_17077_),
    .A2(_17237_),
    .B1(_17235_),
    .X(_17372_));
 sky130_fd_sc_hd__nand2_2 _39434_ (.A(_14153_),
    .B(_10166_),
    .Y(_17373_));
 sky130_fd_sc_hd__or2_2 _39435_ (.A(_17234_),
    .B(_17373_),
    .X(_17374_));
 sky130_fd_sc_hd__nand2_2 _39436_ (.A(_17234_),
    .B(_17373_),
    .Y(_17375_));
 sky130_fd_sc_hd__nand2_2 _39437_ (.A(_17374_),
    .B(_17375_),
    .Y(_17376_));
 sky130_fd_sc_hd__or2_2 _39438_ (.A(_17076_),
    .B(_17376_),
    .X(_17377_));
 sky130_fd_sc_hd__nand2_2 _39439_ (.A(_17376_),
    .B(_17077_),
    .Y(_17378_));
 sky130_fd_sc_hd__nand2_2 _39440_ (.A(_17377_),
    .B(_17378_),
    .Y(_17379_));
 sky130_fd_sc_hd__a21o_2 _39441_ (.A1(_17219_),
    .A2(_17222_),
    .B1(_17379_),
    .X(_17380_));
 sky130_fd_sc_hd__nand3_2 _39442_ (.A(_17379_),
    .B(_17219_),
    .C(_17222_),
    .Y(_17381_));
 sky130_fd_sc_hd__nand2_2 _39443_ (.A(_17380_),
    .B(_17381_),
    .Y(_17382_));
 sky130_fd_sc_hd__xor2_2 _39444_ (.A(_17372_),
    .B(_17382_),
    .X(_17383_));
 sky130_fd_sc_hd__a21o_2 _39445_ (.A1(_17367_),
    .A2(_17371_),
    .B1(_17383_),
    .X(_17384_));
 sky130_fd_sc_hd__nand3_2 _39446_ (.A(_17367_),
    .B(_17371_),
    .C(_17383_),
    .Y(_17385_));
 sky130_fd_sc_hd__o21ai_2 _39447_ (.A1(_17248_),
    .A2(_17232_),
    .B1(_17231_),
    .Y(_17386_));
 sky130_fd_sc_hd__a21oi_2 _39448_ (.A1(_17384_),
    .A2(_17385_),
    .B1(_17386_),
    .Y(_17387_));
 sky130_fd_sc_hd__a21boi_2 _39449_ (.A1(_17250_),
    .A2(_17227_),
    .B1_N(_17231_),
    .Y(_17388_));
 sky130_fd_sc_hd__nand2_2 _39450_ (.A(_17384_),
    .B(_17385_),
    .Y(_17389_));
 sky130_fd_sc_hd__nor2_2 _39451_ (.A(_17388_),
    .B(_17389_),
    .Y(_17390_));
 sky130_fd_sc_hd__o22ai_2 _39452_ (.A1(_17343_),
    .A2(_17345_),
    .B1(_17387_),
    .B2(_17390_),
    .Y(_17391_));
 sky130_fd_sc_hd__a21boi_2 _39453_ (.A1(_17258_),
    .A2(_17265_),
    .B1_N(_17252_),
    .Y(_17392_));
 sky130_fd_sc_hd__nand2_2 _39454_ (.A(_17389_),
    .B(_17388_),
    .Y(_17393_));
 sky130_fd_sc_hd__nand3_2 _39455_ (.A(_17386_),
    .B(_17384_),
    .C(_17385_),
    .Y(_17394_));
 sky130_fd_sc_hd__nand2_2 _39456_ (.A(_17341_),
    .B(_17263_),
    .Y(_17395_));
 sky130_fd_sc_hd__nand3_2 _39457_ (.A(_17339_),
    .B(_17106_),
    .C(_17340_),
    .Y(_17396_));
 sky130_fd_sc_hd__nand2_2 _39458_ (.A(_17395_),
    .B(_17396_),
    .Y(_17397_));
 sky130_fd_sc_hd__nand3_2 _39459_ (.A(_17393_),
    .B(_17394_),
    .C(_17397_),
    .Y(_17398_));
 sky130_fd_sc_hd__nand3_2 _39460_ (.A(_17391_),
    .B(_17392_),
    .C(_17398_),
    .Y(_17399_));
 sky130_fd_sc_hd__inv_2 _39461_ (.A(_17396_),
    .Y(_17400_));
 sky130_fd_sc_hd__inv_2 _39462_ (.A(_17395_),
    .Y(_17401_));
 sky130_fd_sc_hd__o2bb2ai_2 _39463_ (.A1_N(_17394_),
    .A2_N(_17393_),
    .B1(_17400_),
    .B2(_17401_),
    .Y(_17402_));
 sky130_fd_sc_hd__nand2_2 _39464_ (.A(_17206_),
    .B(_17249_),
    .Y(_17403_));
 sky130_fd_sc_hd__o2bb2ai_2 _39465_ (.A1_N(_17258_),
    .A2_N(_17265_),
    .B1(_17256_),
    .B2(_17403_),
    .Y(_17404_));
 sky130_fd_sc_hd__nand3b_2 _39466_ (.A_N(_17397_),
    .B(_17393_),
    .C(_17394_),
    .Y(_17405_));
 sky130_fd_sc_hd__nand3_2 _39467_ (.A(_17402_),
    .B(_17404_),
    .C(_17405_),
    .Y(_17406_));
 sky130_fd_sc_hd__nand3_2 _39468_ (.A(_17259_),
    .B(_17106_),
    .C(_17260_),
    .Y(_17407_));
 sky130_fd_sc_hd__buf_1 _39469_ (.A(_16736_),
    .X(_17408_));
 sky130_fd_sc_hd__nand3_2 _39470_ (.A(_17407_),
    .B(_17408_),
    .C(_17259_),
    .Y(_17409_));
 sky130_fd_sc_hd__nand2_2 _39471_ (.A(_17409_),
    .B(_16902_),
    .Y(_17410_));
 sky130_fd_sc_hd__a21o_2 _39472_ (.A1(_17407_),
    .A2(_17259_),
    .B1(_16736_),
    .X(_17411_));
 sky130_fd_sc_hd__inv_2 _39473_ (.A(_17411_),
    .Y(_17412_));
 sky130_fd_sc_hd__nand2_2 _39474_ (.A(_17411_),
    .B(_17409_),
    .Y(_17413_));
 sky130_fd_sc_hd__nand2_2 _39475_ (.A(_17413_),
    .B(_17135_),
    .Y(_17414_));
 sky130_fd_sc_hd__o21ai_2 _39476_ (.A1(_17410_),
    .A2(_17412_),
    .B1(_17414_),
    .Y(_17415_));
 sky130_fd_sc_hd__nand3_2 _39477_ (.A(_17399_),
    .B(_17406_),
    .C(_17415_),
    .Y(_17416_));
 sky130_fd_sc_hd__and2_2 _39478_ (.A(_17413_),
    .B(_17286_),
    .X(_17417_));
 sky130_fd_sc_hd__nor2_2 _39479_ (.A(_17286_),
    .B(_17413_),
    .Y(_17418_));
 sky130_fd_sc_hd__o2bb2ai_2 _39480_ (.A1_N(_17406_),
    .A2_N(_17399_),
    .B1(_17417_),
    .B2(_17418_),
    .Y(_17419_));
 sky130_fd_sc_hd__a21oi_2 _39481_ (.A1(_17271_),
    .A2(_17272_),
    .B1(_17269_),
    .Y(_17420_));
 sky130_fd_sc_hd__a21oi_2 _39482_ (.A1(_17281_),
    .A2(_17273_),
    .B1(_17420_),
    .Y(_17421_));
 sky130_fd_sc_hd__a21boi_2 _39483_ (.A1(_17416_),
    .A2(_17419_),
    .B1_N(_17421_),
    .Y(_17422_));
 sky130_fd_sc_hd__a31oi_2 _39484_ (.A1(_17271_),
    .A2(_17269_),
    .A3(_17272_),
    .B1(_17280_),
    .Y(_17423_));
 sky130_fd_sc_hd__o211ai_2 _39485_ (.A1(_17420_),
    .A2(_17423_),
    .B1(_17416_),
    .C1(_17419_),
    .Y(_17424_));
 sky130_fd_sc_hd__nand2_2 _39486_ (.A(_17276_),
    .B(_16901_),
    .Y(_17425_));
 sky130_fd_sc_hd__nand2_2 _39487_ (.A(_17425_),
    .B(_17275_),
    .Y(_17426_));
 sky130_fd_sc_hd__inv_2 _39488_ (.A(_17426_),
    .Y(_17427_));
 sky130_fd_sc_hd__nand2_2 _39489_ (.A(_17427_),
    .B(_16083_),
    .Y(_17428_));
 sky130_fd_sc_hd__nand2_2 _39490_ (.A(_17426_),
    .B(_17150_),
    .Y(_17429_));
 sky130_fd_sc_hd__a21oi_2 _39491_ (.A1(_17428_),
    .A2(_17429_),
    .B1(_16844_),
    .Y(_17430_));
 sky130_fd_sc_hd__and3_2 _39492_ (.A(_17428_),
    .B(_16294_),
    .C(_17429_),
    .X(_17431_));
 sky130_fd_sc_hd__nor2_2 _39493_ (.A(_17430_),
    .B(_17431_),
    .Y(_17432_));
 sky130_fd_sc_hd__nand2_2 _39494_ (.A(_17424_),
    .B(_17432_),
    .Y(_17433_));
 sky130_fd_sc_hd__nand2_2 _39495_ (.A(_17295_),
    .B(_17303_),
    .Y(_17434_));
 sky130_fd_sc_hd__o21a_2 _39496_ (.A1(_17412_),
    .A2(_17410_),
    .B1(_17414_),
    .X(_17435_));
 sky130_fd_sc_hd__a21o_2 _39497_ (.A1(_17399_),
    .A2(_17406_),
    .B1(_17435_),
    .X(_17436_));
 sky130_fd_sc_hd__nand3_2 _39498_ (.A(_17435_),
    .B(_17399_),
    .C(_17406_),
    .Y(_17437_));
 sky130_fd_sc_hd__nand3_2 _39499_ (.A(_17436_),
    .B(_17421_),
    .C(_17437_),
    .Y(_17438_));
 sky130_fd_sc_hd__nand2_2 _39500_ (.A(_17438_),
    .B(_17424_),
    .Y(_17439_));
 sky130_fd_sc_hd__inv_2 _39501_ (.A(_17432_),
    .Y(_17440_));
 sky130_fd_sc_hd__nand2_2 _39502_ (.A(_17439_),
    .B(_17440_),
    .Y(_17441_));
 sky130_fd_sc_hd__o2111ai_2 _39503_ (.A1(_17422_),
    .A2(_17433_),
    .B1(_17285_),
    .C1(_17434_),
    .D1(_17441_),
    .Y(_17442_));
 sky130_fd_sc_hd__nand2_2 _39504_ (.A(_17434_),
    .B(_17285_),
    .Y(_17443_));
 sky130_fd_sc_hd__nand2_2 _39505_ (.A(_17439_),
    .B(_17432_),
    .Y(_17444_));
 sky130_fd_sc_hd__nand3_2 _39506_ (.A(_17440_),
    .B(_17438_),
    .C(_17424_),
    .Y(_17445_));
 sky130_fd_sc_hd__nand3_2 _39507_ (.A(_17443_),
    .B(_17444_),
    .C(_17445_),
    .Y(_17446_));
 sky130_fd_sc_hd__nand2_2 _39508_ (.A(_17300_),
    .B(_17298_),
    .Y(_17447_));
 sky130_fd_sc_hd__nor2_2 _39509_ (.A(_16120_),
    .B(_17447_),
    .Y(_17448_));
 sky130_fd_sc_hd__inv_2 _39510_ (.A(_17447_),
    .Y(_17449_));
 sky130_fd_sc_hd__nor2_2 _39511_ (.A(_16118_),
    .B(_17449_),
    .Y(_17450_));
 sky130_fd_sc_hd__nor2_2 _39512_ (.A(_17448_),
    .B(_17450_),
    .Y(_17451_));
 sky130_fd_sc_hd__nand3_2 _39513_ (.A(_17442_),
    .B(_17446_),
    .C(_17451_),
    .Y(_17452_));
 sky130_fd_sc_hd__o2bb2ai_2 _39514_ (.A1_N(_17446_),
    .A2_N(_17442_),
    .B1(_17450_),
    .B2(_17448_),
    .Y(_17453_));
 sky130_fd_sc_hd__o211ai_2 _39515_ (.A1(_17337_),
    .A2(_17321_),
    .B1(_17452_),
    .C1(_17453_),
    .Y(_17454_));
 sky130_fd_sc_hd__a21oi_2 _39516_ (.A1(_17311_),
    .A2(_17318_),
    .B1(_17337_),
    .Y(_17455_));
 sky130_fd_sc_hd__nor2_2 _39517_ (.A(_14019_),
    .B(_17447_),
    .Y(_17456_));
 sky130_fd_sc_hd__nor2_2 _39518_ (.A(_17164_),
    .B(_17449_),
    .Y(_17457_));
 sky130_fd_sc_hd__o2bb2ai_2 _39519_ (.A1_N(_17446_),
    .A2_N(_17442_),
    .B1(_17456_),
    .B2(_17457_),
    .Y(_17458_));
 sky130_fd_sc_hd__nand3b_2 _39520_ (.A_N(_17451_),
    .B(_17442_),
    .C(_17446_),
    .Y(_17459_));
 sky130_fd_sc_hd__nand3_2 _39521_ (.A(_17455_),
    .B(_17458_),
    .C(_17459_),
    .Y(_17460_));
 sky130_fd_sc_hd__a21oi_2 _39522_ (.A1(_17454_),
    .A2(_17460_),
    .B1(_17315_),
    .Y(_17461_));
 sky130_fd_sc_hd__and3_2 _39523_ (.A(_17454_),
    .B(_17460_),
    .C(_17315_),
    .X(_17462_));
 sky130_fd_sc_hd__a21boi_2 _39524_ (.A1(_17163_),
    .A2(_17327_),
    .B1_N(_17323_),
    .Y(_17463_));
 sky130_fd_sc_hd__o21ai_2 _39525_ (.A1(_17461_),
    .A2(_17462_),
    .B1(_17463_),
    .Y(_17464_));
 sky130_fd_sc_hd__nand2_2 _39526_ (.A(_17327_),
    .B(_17163_),
    .Y(_17465_));
 sky130_fd_sc_hd__nand2_2 _39527_ (.A(_17465_),
    .B(_17323_),
    .Y(_17466_));
 sky130_fd_sc_hd__nand3_2 _39528_ (.A(_17454_),
    .B(_17460_),
    .C(_17315_),
    .Y(_17467_));
 sky130_fd_sc_hd__a21o_2 _39529_ (.A1(_17454_),
    .A2(_17460_),
    .B1(_17315_),
    .X(_17468_));
 sky130_fd_sc_hd__nand3_2 _39530_ (.A(_17466_),
    .B(_17467_),
    .C(_17468_),
    .Y(_17469_));
 sky130_fd_sc_hd__and2_2 _39531_ (.A(_17464_),
    .B(_17469_),
    .X(_17470_));
 sky130_fd_sc_hd__nand2_2 _39532_ (.A(_17334_),
    .B(_17187_),
    .Y(_17471_));
 sky130_fd_sc_hd__a21oi_2 _39533_ (.A1(_15747_),
    .A2(_17190_),
    .B1(_17198_),
    .Y(_17472_));
 sky130_fd_sc_hd__nand3_2 _39534_ (.A(_17331_),
    .B(_17328_),
    .C(_17329_),
    .Y(_17473_));
 sky130_fd_sc_hd__nand2_2 _39535_ (.A(_17473_),
    .B(_17335_),
    .Y(_17474_));
 sky130_fd_sc_hd__a21o_2 _39536_ (.A1(_17328_),
    .A2(_17329_),
    .B1(_17331_),
    .X(_17475_));
 sky130_fd_sc_hd__nand2_2 _39537_ (.A(_17474_),
    .B(_17475_),
    .Y(_17476_));
 sky130_fd_sc_hd__o21ai_2 _39538_ (.A1(_17471_),
    .A2(_17472_),
    .B1(_17476_),
    .Y(_17477_));
 sky130_fd_sc_hd__or2_2 _39539_ (.A(_17470_),
    .B(_17477_),
    .X(_17478_));
 sky130_fd_sc_hd__nand2_2 _39540_ (.A(_17477_),
    .B(_17470_),
    .Y(_17479_));
 sky130_fd_sc_hd__and2_2 _39541_ (.A(_17478_),
    .B(_17479_),
    .X(_02677_));
 sky130_fd_sc_hd__nand2_2 _39542_ (.A(_17410_),
    .B(_17411_),
    .Y(_17480_));
 sky130_fd_sc_hd__or2_2 _39543_ (.A(_17150_),
    .B(_17480_),
    .X(_17481_));
 sky130_fd_sc_hd__nand2_2 _39544_ (.A(_17480_),
    .B(_17150_),
    .Y(_17482_));
 sky130_fd_sc_hd__and3_2 _39545_ (.A(_17481_),
    .B(_16844_),
    .C(_17482_),
    .X(_17483_));
 sky130_fd_sc_hd__buf_1 _39546_ (.A(_16844_),
    .X(_17484_));
 sky130_fd_sc_hd__a21oi_2 _39547_ (.A1(_17481_),
    .A2(_17482_),
    .B1(_17484_),
    .Y(_17485_));
 sky130_fd_sc_hd__nor2_2 _39548_ (.A(_10152_),
    .B(_11036_),
    .Y(_17486_));
 sky130_fd_sc_hd__inv_2 _39549_ (.A(_17486_),
    .Y(_17487_));
 sky130_fd_sc_hd__or4_2 _39550_ (.A(_19560_),
    .B(_18183_),
    .C(_17048_),
    .D(_10543_),
    .X(_17488_));
 sky130_fd_sc_hd__a22o_2 _39551_ (.A1(_19310_),
    .A2(_19555_),
    .B1(_14939_),
    .B2(_11123_),
    .X(_17489_));
 sky130_fd_sc_hd__nand2_2 _39552_ (.A(_17488_),
    .B(_17489_),
    .Y(_17490_));
 sky130_fd_sc_hd__or2_2 _39553_ (.A(_17487_),
    .B(_17490_),
    .X(_17491_));
 sky130_fd_sc_hd__nand2_2 _39554_ (.A(_17490_),
    .B(_17487_),
    .Y(_17492_));
 sky130_fd_sc_hd__o21a_2 _39555_ (.A1(_17355_),
    .A2(_17351_),
    .B1(_17349_),
    .X(_17493_));
 sky130_fd_sc_hd__a21o_2 _39556_ (.A1(_17491_),
    .A2(_17492_),
    .B1(_17493_),
    .X(_17494_));
 sky130_fd_sc_hd__nand3_2 _39557_ (.A(_17491_),
    .B(_17493_),
    .C(_17492_),
    .Y(_17495_));
 sky130_fd_sc_hd__nand2_2 _39558_ (.A(_17494_),
    .B(_17495_),
    .Y(_17496_));
 sky130_fd_sc_hd__nand2_2 _39559_ (.A(_18158_),
    .B(_19325_),
    .Y(_17497_));
 sky130_fd_sc_hd__and4_2 _39560_ (.A(_19318_),
    .B(_19321_),
    .C(_19542_),
    .D(_19547_),
    .X(_17498_));
 sky130_fd_sc_hd__o22a_2 _39561_ (.A1(_14371_),
    .A2(_11764_),
    .B1(_14869_),
    .B2(_15116_),
    .X(_17499_));
 sky130_fd_sc_hd__or3_2 _39562_ (.A(_17497_),
    .B(_17498_),
    .C(_17499_),
    .X(_17500_));
 sky130_fd_sc_hd__buf_1 _39563_ (.A(_17497_),
    .X(_17501_));
 sky130_fd_sc_hd__o21ai_2 _39564_ (.A1(_17498_),
    .A2(_17499_),
    .B1(_17501_),
    .Y(_17502_));
 sky130_fd_sc_hd__nand2_2 _39565_ (.A(_17500_),
    .B(_17502_),
    .Y(_17503_));
 sky130_fd_sc_hd__nand2_2 _39566_ (.A(_17496_),
    .B(_17503_),
    .Y(_17504_));
 sky130_fd_sc_hd__a21boi_2 _39567_ (.A1(_17354_),
    .A2(_17364_),
    .B1_N(_17358_),
    .Y(_17505_));
 sky130_fd_sc_hd__inv_2 _39568_ (.A(_17503_),
    .Y(_17506_));
 sky130_fd_sc_hd__nand3_2 _39569_ (.A(_17494_),
    .B(_17495_),
    .C(_17506_),
    .Y(_17507_));
 sky130_fd_sc_hd__nand3_2 _39570_ (.A(_17504_),
    .B(_17505_),
    .C(_17507_),
    .Y(_17508_));
 sky130_fd_sc_hd__nand2_2 _39571_ (.A(_17496_),
    .B(_17506_),
    .Y(_17509_));
 sky130_fd_sc_hd__nand3_2 _39572_ (.A(_17494_),
    .B(_17495_),
    .C(_17503_),
    .Y(_17510_));
 sky130_fd_sc_hd__nand3b_2 _39573_ (.A_N(_17505_),
    .B(_17509_),
    .C(_17510_),
    .Y(_17511_));
 sky130_fd_sc_hd__nand2_2 _39574_ (.A(_17377_),
    .B(_17374_),
    .Y(_17512_));
 sky130_fd_sc_hd__inv_2 _39575_ (.A(_17512_),
    .Y(_17513_));
 sky130_fd_sc_hd__buf_1 _39576_ (.A(_17513_),
    .X(_17514_));
 sky130_fd_sc_hd__o21ai_2 _39577_ (.A1(_16003_),
    .A2(_10539_),
    .B1(_17362_),
    .Y(_17515_));
 sky130_fd_sc_hd__and2_2 _39578_ (.A(_17377_),
    .B(_17378_),
    .X(_17516_));
 sky130_fd_sc_hd__or2_2 _39579_ (.A(_17515_),
    .B(_17516_),
    .X(_17517_));
 sky130_fd_sc_hd__buf_1 _39580_ (.A(_17516_),
    .X(_17518_));
 sky130_fd_sc_hd__nand2_2 _39581_ (.A(_17518_),
    .B(_17515_),
    .Y(_17519_));
 sky130_fd_sc_hd__nand2_2 _39582_ (.A(_17517_),
    .B(_17519_),
    .Y(_17520_));
 sky130_fd_sc_hd__nor2_2 _39583_ (.A(_17514_),
    .B(_17520_),
    .Y(_17521_));
 sky130_fd_sc_hd__buf_1 _39584_ (.A(_17513_),
    .X(_17522_));
 sky130_fd_sc_hd__and2_2 _39585_ (.A(_17520_),
    .B(_17522_),
    .X(_17523_));
 sky130_fd_sc_hd__o2bb2ai_2 _39586_ (.A1_N(_17508_),
    .A2_N(_17511_),
    .B1(_17521_),
    .B2(_17523_),
    .Y(_17524_));
 sky130_fd_sc_hd__nand2_2 _39587_ (.A(_17520_),
    .B(_17512_),
    .Y(_17525_));
 sky130_fd_sc_hd__nand3_2 _39588_ (.A(_17517_),
    .B(_17519_),
    .C(_17514_),
    .Y(_17526_));
 sky130_fd_sc_hd__nand2_2 _39589_ (.A(_17525_),
    .B(_17526_),
    .Y(_17527_));
 sky130_fd_sc_hd__nand3_2 _39590_ (.A(_17511_),
    .B(_17508_),
    .C(_17527_),
    .Y(_17528_));
 sky130_fd_sc_hd__nand2_2 _39591_ (.A(_17385_),
    .B(_17367_),
    .Y(_17529_));
 sky130_fd_sc_hd__a21oi_2 _39592_ (.A1(_17524_),
    .A2(_17528_),
    .B1(_17529_),
    .Y(_17530_));
 sky130_fd_sc_hd__a21oi_2 _39593_ (.A1(_17370_),
    .A2(_17369_),
    .B1(_17368_),
    .Y(_17531_));
 sky130_fd_sc_hd__a21oi_2 _39594_ (.A1(_17371_),
    .A2(_17383_),
    .B1(_17531_),
    .Y(_17532_));
 sky130_fd_sc_hd__a21oi_2 _39595_ (.A1(_17511_),
    .A2(_17508_),
    .B1(_17527_),
    .Y(_17533_));
 sky130_fd_sc_hd__and3_2 _39596_ (.A(_17511_),
    .B(_17508_),
    .C(_17527_),
    .X(_17534_));
 sky130_fd_sc_hd__nor3_2 _39597_ (.A(_17532_),
    .B(_17533_),
    .C(_17534_),
    .Y(_17535_));
 sky130_fd_sc_hd__inv_2 _39598_ (.A(_17107_),
    .Y(_17536_));
 sky130_fd_sc_hd__nor2_2 _39599_ (.A(_17108_),
    .B(_17536_),
    .Y(_17537_));
 sky130_fd_sc_hd__or2_2 _39600_ (.A(_17372_),
    .B(_17382_),
    .X(_17538_));
 sky130_fd_sc_hd__nand2_2 _39601_ (.A(_17538_),
    .B(_17380_),
    .Y(_17539_));
 sky130_fd_sc_hd__nor2_2 _39602_ (.A(_17537_),
    .B(_17539_),
    .Y(_17540_));
 sky130_fd_sc_hd__and2_2 _39603_ (.A(_17539_),
    .B(_17537_),
    .X(_17541_));
 sky130_fd_sc_hd__nor2_2 _39604_ (.A(_17540_),
    .B(_17541_),
    .Y(_17542_));
 sky130_fd_sc_hd__o21bai_2 _39605_ (.A1(_17530_),
    .A2(_17535_),
    .B1_N(_17542_),
    .Y(_17543_));
 sky130_fd_sc_hd__o21ai_2 _39606_ (.A1(_17533_),
    .A2(_17534_),
    .B1(_17532_),
    .Y(_17544_));
 sky130_fd_sc_hd__nand3_2 _39607_ (.A(_17529_),
    .B(_17524_),
    .C(_17528_),
    .Y(_17545_));
 sky130_fd_sc_hd__nand3_2 _39608_ (.A(_17544_),
    .B(_17545_),
    .C(_17542_),
    .Y(_17546_));
 sky130_fd_sc_hd__o21ai_2 _39609_ (.A1(_17397_),
    .A2(_17387_),
    .B1(_17394_),
    .Y(_17547_));
 sky130_fd_sc_hd__a21oi_2 _39610_ (.A1(_17543_),
    .A2(_17546_),
    .B1(_17547_),
    .Y(_17548_));
 sky130_fd_sc_hd__a22oi_2 _39611_ (.A1(_17342_),
    .A2(_17344_),
    .B1(_17389_),
    .B2(_17388_),
    .Y(_17549_));
 sky130_fd_sc_hd__o211a_2 _39612_ (.A1(_17390_),
    .A2(_17549_),
    .B1(_17546_),
    .C1(_17543_),
    .X(_17550_));
 sky130_fd_sc_hd__a21o_2 _39613_ (.A1(_17396_),
    .A2(_17339_),
    .B1(_17408_),
    .X(_17551_));
 sky130_fd_sc_hd__nand3_2 _39614_ (.A(_17396_),
    .B(_17408_),
    .C(_17339_),
    .Y(_17552_));
 sky130_fd_sc_hd__a21o_2 _39615_ (.A1(_17551_),
    .A2(_17552_),
    .B1(_17135_),
    .X(_17553_));
 sky130_fd_sc_hd__nand3_2 _39616_ (.A(_17551_),
    .B(_17552_),
    .C(_17135_),
    .Y(_17554_));
 sky130_fd_sc_hd__nand2_2 _39617_ (.A(_17553_),
    .B(_17554_),
    .Y(_17555_));
 sky130_fd_sc_hd__o21bai_2 _39618_ (.A1(_17548_),
    .A2(_17550_),
    .B1_N(_17555_),
    .Y(_17556_));
 sky130_fd_sc_hd__a21o_2 _39619_ (.A1(_17543_),
    .A2(_17546_),
    .B1(_17547_),
    .X(_17557_));
 sky130_fd_sc_hd__nand3_2 _39620_ (.A(_17547_),
    .B(_17543_),
    .C(_17546_),
    .Y(_17558_));
 sky130_fd_sc_hd__nand3_2 _39621_ (.A(_17557_),
    .B(_17558_),
    .C(_17555_),
    .Y(_17559_));
 sky130_fd_sc_hd__nand2_2 _39622_ (.A(_17435_),
    .B(_17399_),
    .Y(_17560_));
 sky130_fd_sc_hd__nand2_2 _39623_ (.A(_17560_),
    .B(_17406_),
    .Y(_17561_));
 sky130_fd_sc_hd__a21oi_2 _39624_ (.A1(_17556_),
    .A2(_17559_),
    .B1(_17561_),
    .Y(_17562_));
 sky130_fd_sc_hd__inv_2 _39625_ (.A(_17406_),
    .Y(_17563_));
 sky130_fd_sc_hd__a31oi_2 _39626_ (.A1(_17392_),
    .A2(_17391_),
    .A3(_17398_),
    .B1(_17415_),
    .Y(_17564_));
 sky130_fd_sc_hd__o211a_2 _39627_ (.A1(_17563_),
    .A2(_17564_),
    .B1(_17559_),
    .C1(_17556_),
    .X(_17565_));
 sky130_fd_sc_hd__o22ai_2 _39628_ (.A1(_17483_),
    .A2(_17485_),
    .B1(_17562_),
    .B2(_17565_),
    .Y(_17566_));
 sky130_fd_sc_hd__a21o_2 _39629_ (.A1(_17556_),
    .A2(_17559_),
    .B1(_17561_),
    .X(_17567_));
 sky130_fd_sc_hd__nand3_2 _39630_ (.A(_17561_),
    .B(_17556_),
    .C(_17559_),
    .Y(_17568_));
 sky130_fd_sc_hd__nor2_2 _39631_ (.A(_17485_),
    .B(_17483_),
    .Y(_17569_));
 sky130_fd_sc_hd__nand3_2 _39632_ (.A(_17567_),
    .B(_17568_),
    .C(_17569_),
    .Y(_17570_));
 sky130_fd_sc_hd__nand2_2 _39633_ (.A(_17433_),
    .B(_17438_),
    .Y(_17571_));
 sky130_fd_sc_hd__a21oi_2 _39634_ (.A1(_17566_),
    .A2(_17570_),
    .B1(_17571_),
    .Y(_17572_));
 sky130_fd_sc_hd__and2_2 _39635_ (.A(_17424_),
    .B(_17432_),
    .X(_17573_));
 sky130_fd_sc_hd__o211a_2 _39636_ (.A1(_17422_),
    .A2(_17573_),
    .B1(_17570_),
    .C1(_17566_),
    .X(_17574_));
 sky130_fd_sc_hd__nand2_2 _39637_ (.A(_17428_),
    .B(_17484_),
    .Y(_17575_));
 sky130_fd_sc_hd__nand2_2 _39638_ (.A(_17575_),
    .B(_17429_),
    .Y(_17576_));
 sky130_fd_sc_hd__nor2_2 _39639_ (.A(_17164_),
    .B(_17576_),
    .Y(_17577_));
 sky130_fd_sc_hd__and2_2 _39640_ (.A(_17576_),
    .B(_15109_),
    .X(_17578_));
 sky130_fd_sc_hd__nor2_2 _39641_ (.A(_17577_),
    .B(_17578_),
    .Y(_17579_));
 sky130_fd_sc_hd__o21ai_2 _39642_ (.A1(_17572_),
    .A2(_17574_),
    .B1(_17579_),
    .Y(_17580_));
 sky130_fd_sc_hd__a21boi_2 _39643_ (.A1(_17446_),
    .A2(_17451_),
    .B1_N(_17442_),
    .Y(_17581_));
 sky130_fd_sc_hd__a21o_2 _39644_ (.A1(_17566_),
    .A2(_17570_),
    .B1(_17571_),
    .X(_17582_));
 sky130_fd_sc_hd__nand3_2 _39645_ (.A(_17566_),
    .B(_17570_),
    .C(_17571_),
    .Y(_17583_));
 sky130_fd_sc_hd__nand3b_2 _39646_ (.A_N(_17579_),
    .B(_17582_),
    .C(_17583_),
    .Y(_17584_));
 sky130_fd_sc_hd__nand3_2 _39647_ (.A(_17580_),
    .B(_17581_),
    .C(_17584_),
    .Y(_17585_));
 sky130_fd_sc_hd__o22ai_2 _39648_ (.A1(_17578_),
    .A2(_17577_),
    .B1(_17572_),
    .B2(_17574_),
    .Y(_17586_));
 sky130_fd_sc_hd__nand2_2 _39649_ (.A(_17446_),
    .B(_17451_),
    .Y(_17587_));
 sky130_fd_sc_hd__nand2_2 _39650_ (.A(_17587_),
    .B(_17442_),
    .Y(_17588_));
 sky130_fd_sc_hd__nand3_2 _39651_ (.A(_17582_),
    .B(_17583_),
    .C(_17579_),
    .Y(_17589_));
 sky130_fd_sc_hd__nand3_2 _39652_ (.A(_17586_),
    .B(_17588_),
    .C(_17589_),
    .Y(_17590_));
 sky130_fd_sc_hd__and3_2 _39653_ (.A(_17585_),
    .B(_17590_),
    .C(_17450_),
    .X(_17591_));
 sky130_fd_sc_hd__o2bb2ai_2 _39654_ (.A1_N(_17585_),
    .A2_N(_17590_),
    .B1(_17180_),
    .B2(_17449_),
    .Y(_17592_));
 sky130_fd_sc_hd__nand2_2 _39655_ (.A(_17460_),
    .B(_17315_),
    .Y(_17593_));
 sky130_fd_sc_hd__nand2_2 _39656_ (.A(_17593_),
    .B(_17454_),
    .Y(_17594_));
 sky130_fd_sc_hd__nand2_2 _39657_ (.A(_17592_),
    .B(_17594_),
    .Y(_17595_));
 sky130_fd_sc_hd__a21oi_2 _39658_ (.A1(_17585_),
    .A2(_17590_),
    .B1(_17450_),
    .Y(_17596_));
 sky130_fd_sc_hd__o21bai_2 _39659_ (.A1(_17596_),
    .A2(_17591_),
    .B1_N(_17594_),
    .Y(_17597_));
 sky130_fd_sc_hd__o21a_2 _39660_ (.A1(_17591_),
    .A2(_17595_),
    .B1(_17597_),
    .X(_17598_));
 sky130_fd_sc_hd__a21o_2 _39661_ (.A1(_17479_),
    .A2(_17469_),
    .B1(_17598_),
    .X(_17599_));
 sky130_fd_sc_hd__nand3_2 _39662_ (.A(_17479_),
    .B(_17469_),
    .C(_17598_),
    .Y(_17600_));
 sky130_fd_sc_hd__nand2_2 _39663_ (.A(_17599_),
    .B(_17600_),
    .Y(_02678_));
 sky130_fd_sc_hd__a21o_2 _39664_ (.A1(_17582_),
    .A2(_17579_),
    .B1(_17574_),
    .X(_17601_));
 sky130_fd_sc_hd__nand2_2 _39665_ (.A(_17546_),
    .B(_17545_),
    .Y(_17602_));
 sky130_fd_sc_hd__and2_2 _39666_ (.A(_17528_),
    .B(_17511_),
    .X(_17603_));
 sky130_fd_sc_hd__nor2_2 _39667_ (.A(_11913_),
    .B(_14869_),
    .Y(_17604_));
 sky130_fd_sc_hd__a21oi_2 _39668_ (.A1(_19318_),
    .A2(_19543_),
    .B1(_17604_),
    .Y(_17605_));
 sky130_fd_sc_hd__and3_2 _39669_ (.A(_17604_),
    .B(_19318_),
    .C(_19543_),
    .X(_17606_));
 sky130_fd_sc_hd__or3_2 _39670_ (.A(_17501_),
    .B(_17605_),
    .C(_17606_),
    .X(_17607_));
 sky130_fd_sc_hd__o21ai_2 _39671_ (.A1(_17605_),
    .A2(_17606_),
    .B1(_17501_),
    .Y(_17608_));
 sky130_fd_sc_hd__and2_2 _39672_ (.A(_17491_),
    .B(_17488_),
    .X(_17609_));
 sky130_fd_sc_hd__nand2_2 _39673_ (.A(_19314_),
    .B(_19547_),
    .Y(_17610_));
 sky130_fd_sc_hd__or4_2 _39674_ (.A(_19555_),
    .B(_18184_),
    .C(_17048_),
    .D(_11036_),
    .X(_17611_));
 sky130_fd_sc_hd__a22o_2 _39675_ (.A1(_19310_),
    .A2(_19551_),
    .B1(_10543_),
    .B2(_11123_),
    .X(_17612_));
 sky130_fd_sc_hd__nand2_2 _39676_ (.A(_17611_),
    .B(_17612_),
    .Y(_17613_));
 sky130_fd_sc_hd__or2_2 _39677_ (.A(_17610_),
    .B(_17613_),
    .X(_17614_));
 sky130_fd_sc_hd__nand2_2 _39678_ (.A(_17613_),
    .B(_17610_),
    .Y(_17615_));
 sky130_fd_sc_hd__nand2_2 _39679_ (.A(_17614_),
    .B(_17615_),
    .Y(_17616_));
 sky130_fd_sc_hd__nand2_2 _39680_ (.A(_17609_),
    .B(_17616_),
    .Y(_17617_));
 sky130_fd_sc_hd__a21o_2 _39681_ (.A1(_17488_),
    .A2(_17491_),
    .B1(_17616_),
    .X(_17618_));
 sky130_fd_sc_hd__nand2_2 _39682_ (.A(_17617_),
    .B(_17618_),
    .Y(_17619_));
 sky130_fd_sc_hd__a21o_2 _39683_ (.A1(_17607_),
    .A2(_17608_),
    .B1(_17619_),
    .X(_17620_));
 sky130_fd_sc_hd__nand2_2 _39684_ (.A(_17607_),
    .B(_17608_),
    .Y(_17621_));
 sky130_fd_sc_hd__inv_2 _39685_ (.A(_17621_),
    .Y(_17622_));
 sky130_fd_sc_hd__nand2_2 _39686_ (.A(_17619_),
    .B(_17622_),
    .Y(_17623_));
 sky130_fd_sc_hd__nand2_2 _39687_ (.A(_17491_),
    .B(_17492_),
    .Y(_17624_));
 sky130_fd_sc_hd__o21a_2 _39688_ (.A1(_17493_),
    .A2(_17624_),
    .B1(_17509_),
    .X(_17625_));
 sky130_fd_sc_hd__a21o_2 _39689_ (.A1(_17620_),
    .A2(_17623_),
    .B1(_17625_),
    .X(_17626_));
 sky130_fd_sc_hd__nand3_2 _39690_ (.A(_17620_),
    .B(_17625_),
    .C(_17623_),
    .Y(_17627_));
 sky130_fd_sc_hd__o21bai_2 _39691_ (.A1(_17501_),
    .A2(_17499_),
    .B1_N(_17498_),
    .Y(_17628_));
 sky130_fd_sc_hd__or2_2 _39692_ (.A(_17628_),
    .B(_17518_),
    .X(_17629_));
 sky130_fd_sc_hd__nand2_2 _39693_ (.A(_17518_),
    .B(_17628_),
    .Y(_17630_));
 sky130_fd_sc_hd__nand2_2 _39694_ (.A(_17629_),
    .B(_17630_),
    .Y(_17631_));
 sky130_fd_sc_hd__or2_2 _39695_ (.A(_17514_),
    .B(_17631_),
    .X(_17632_));
 sky130_fd_sc_hd__nand2_2 _39696_ (.A(_17631_),
    .B(_17522_),
    .Y(_17633_));
 sky130_fd_sc_hd__and2_2 _39697_ (.A(_17632_),
    .B(_17633_),
    .X(_17634_));
 sky130_fd_sc_hd__a21o_2 _39698_ (.A1(_17626_),
    .A2(_17627_),
    .B1(_17634_),
    .X(_17635_));
 sky130_fd_sc_hd__nand3_2 _39699_ (.A(_17626_),
    .B(_17634_),
    .C(_17627_),
    .Y(_17636_));
 sky130_fd_sc_hd__nand3b_2 _39700_ (.A_N(_17603_),
    .B(_17635_),
    .C(_17636_),
    .Y(_17637_));
 sky130_fd_sc_hd__nand2_2 _39701_ (.A(_17632_),
    .B(_17633_),
    .Y(_17638_));
 sky130_fd_sc_hd__a21o_2 _39702_ (.A1(_17626_),
    .A2(_17627_),
    .B1(_17638_),
    .X(_17639_));
 sky130_fd_sc_hd__nand3_2 _39703_ (.A(_17626_),
    .B(_17638_),
    .C(_17627_),
    .Y(_17640_));
 sky130_fd_sc_hd__nand3_2 _39704_ (.A(_17639_),
    .B(_17640_),
    .C(_17603_),
    .Y(_17641_));
 sky130_fd_sc_hd__or3b_2 _39705_ (.A(_17111_),
    .B(_17521_),
    .C_N(_17519_),
    .X(_17642_));
 sky130_fd_sc_hd__or2_2 _39706_ (.A(_17514_),
    .B(_17520_),
    .X(_17643_));
 sky130_fd_sc_hd__buf_1 _39707_ (.A(_17109_),
    .X(_17644_));
 sky130_fd_sc_hd__a21o_2 _39708_ (.A1(_17643_),
    .A2(_17519_),
    .B1(_17644_),
    .X(_17645_));
 sky130_fd_sc_hd__nand2_2 _39709_ (.A(_17642_),
    .B(_17645_),
    .Y(_17646_));
 sky130_fd_sc_hd__nand2_2 _39710_ (.A(_17646_),
    .B(_17263_),
    .Y(_17647_));
 sky130_fd_sc_hd__a21oi_2 _39711_ (.A1(_17643_),
    .A2(_17519_),
    .B1(_17644_),
    .Y(_17648_));
 sky130_fd_sc_hd__and3_2 _39712_ (.A(_17643_),
    .B(_17644_),
    .C(_17519_),
    .X(_17649_));
 sky130_fd_sc_hd__nor2_2 _39713_ (.A(_17648_),
    .B(_17649_),
    .Y(_17650_));
 sky130_fd_sc_hd__buf_1 _39714_ (.A(_17106_),
    .X(_17651_));
 sky130_fd_sc_hd__nand2_2 _39715_ (.A(_17650_),
    .B(_17651_),
    .Y(_17652_));
 sky130_fd_sc_hd__nand2_2 _39716_ (.A(_17647_),
    .B(_17652_),
    .Y(_17653_));
 sky130_fd_sc_hd__a21o_2 _39717_ (.A1(_17637_),
    .A2(_17641_),
    .B1(_17653_),
    .X(_17654_));
 sky130_fd_sc_hd__nand3_2 _39718_ (.A(_17637_),
    .B(_17641_),
    .C(_17653_),
    .Y(_17655_));
 sky130_fd_sc_hd__nand3b_2 _39719_ (.A_N(_17602_),
    .B(_17654_),
    .C(_17655_),
    .Y(_17656_));
 sky130_fd_sc_hd__nand2_2 _39720_ (.A(_17646_),
    .B(_17651_),
    .Y(_17657_));
 sky130_fd_sc_hd__nand2_2 _39721_ (.A(_17650_),
    .B(_17263_),
    .Y(_17658_));
 sky130_fd_sc_hd__nand2_2 _39722_ (.A(_17657_),
    .B(_17658_),
    .Y(_17659_));
 sky130_fd_sc_hd__a21o_2 _39723_ (.A1(_17637_),
    .A2(_17641_),
    .B1(_17659_),
    .X(_17660_));
 sky130_fd_sc_hd__nand3_2 _39724_ (.A(_17637_),
    .B(_17641_),
    .C(_17659_),
    .Y(_17661_));
 sky130_fd_sc_hd__nand3_2 _39725_ (.A(_17660_),
    .B(_17602_),
    .C(_17661_),
    .Y(_17662_));
 sky130_fd_sc_hd__inv_2 _39726_ (.A(_17108_),
    .Y(_17663_));
 sky130_fd_sc_hd__a21o_2 _39727_ (.A1(_17539_),
    .A2(_17663_),
    .B1(_17536_),
    .X(_17664_));
 sky130_fd_sc_hd__or2_2 _39728_ (.A(_17130_),
    .B(_17664_),
    .X(_17665_));
 sky130_fd_sc_hd__nand2_2 _39729_ (.A(_17664_),
    .B(_17130_),
    .Y(_17666_));
 sky130_fd_sc_hd__and2_2 _39730_ (.A(_17665_),
    .B(_17666_),
    .X(_17667_));
 sky130_fd_sc_hd__nor2_2 _39731_ (.A(_17286_),
    .B(_17667_),
    .Y(_17668_));
 sky130_fd_sc_hd__nand2_2 _39732_ (.A(_17667_),
    .B(_17286_),
    .Y(_17669_));
 sky130_fd_sc_hd__and2b_2 _39733_ (.A_N(_17668_),
    .B(_17669_),
    .X(_17670_));
 sky130_fd_sc_hd__a21o_2 _39734_ (.A1(_17656_),
    .A2(_17662_),
    .B1(_17670_),
    .X(_17671_));
 sky130_fd_sc_hd__nand3_2 _39735_ (.A(_17656_),
    .B(_17670_),
    .C(_17662_),
    .Y(_17672_));
 sky130_fd_sc_hd__a21o_2 _39736_ (.A1(_17557_),
    .A2(_17555_),
    .B1(_17550_),
    .X(_17673_));
 sky130_fd_sc_hd__a21o_2 _39737_ (.A1(_17671_),
    .A2(_17672_),
    .B1(_17673_),
    .X(_17674_));
 sky130_fd_sc_hd__nand3_2 _39738_ (.A(_17671_),
    .B(_17672_),
    .C(_17673_),
    .Y(_17675_));
 sky130_fd_sc_hd__a21bo_2 _39739_ (.A1(_16902_),
    .A2(_17552_),
    .B1_N(_17551_),
    .X(_17676_));
 sky130_fd_sc_hd__or2_2 _39740_ (.A(_17150_),
    .B(_17676_),
    .X(_17677_));
 sky130_fd_sc_hd__buf_1 _39741_ (.A(_17150_),
    .X(_17678_));
 sky130_fd_sc_hd__nand2_2 _39742_ (.A(_17676_),
    .B(_17678_),
    .Y(_17679_));
 sky130_fd_sc_hd__nand2_2 _39743_ (.A(_17677_),
    .B(_17679_),
    .Y(_17680_));
 sky130_fd_sc_hd__or2b_2 _39744_ (.A(_17680_),
    .B_N(_17484_),
    .X(_17681_));
 sky130_fd_sc_hd__nand2_2 _39745_ (.A(_17680_),
    .B(_17147_),
    .Y(_17682_));
 sky130_fd_sc_hd__and2_2 _39746_ (.A(_17681_),
    .B(_17682_),
    .X(_17683_));
 sky130_fd_sc_hd__a21o_2 _39747_ (.A1(_17674_),
    .A2(_17675_),
    .B1(_17683_),
    .X(_17684_));
 sky130_fd_sc_hd__nand2_2 _39748_ (.A(_17570_),
    .B(_17568_),
    .Y(_17685_));
 sky130_fd_sc_hd__nand3_2 _39749_ (.A(_17683_),
    .B(_17674_),
    .C(_17675_),
    .Y(_17686_));
 sky130_fd_sc_hd__nand3_2 _39750_ (.A(_17684_),
    .B(_17685_),
    .C(_17686_),
    .Y(_17687_));
 sky130_fd_sc_hd__a21oi_2 _39751_ (.A1(_17674_),
    .A2(_17675_),
    .B1(_17683_),
    .Y(_17688_));
 sky130_fd_sc_hd__nand2_2 _39752_ (.A(_17681_),
    .B(_17682_),
    .Y(_17689_));
 sky130_fd_sc_hd__a21oi_2 _39753_ (.A1(_17671_),
    .A2(_17672_),
    .B1(_17673_),
    .Y(_17690_));
 sky130_fd_sc_hd__nor3b_2 _39754_ (.A(_17689_),
    .B(_17690_),
    .C_N(_17675_),
    .Y(_17691_));
 sky130_fd_sc_hd__o21bai_2 _39755_ (.A1(_17688_),
    .A2(_17691_),
    .B1_N(_17685_),
    .Y(_17692_));
 sky130_fd_sc_hd__nand2_2 _39756_ (.A(_17481_),
    .B(_17484_),
    .Y(_17693_));
 sky130_fd_sc_hd__nand2_2 _39757_ (.A(_17693_),
    .B(_17482_),
    .Y(_17694_));
 sky130_fd_sc_hd__nor2_2 _39758_ (.A(_15320_),
    .B(_17694_),
    .Y(_17695_));
 sky130_fd_sc_hd__inv_2 _39759_ (.A(_17694_),
    .Y(_17696_));
 sky130_fd_sc_hd__nor2_2 _39760_ (.A(_17165_),
    .B(_17696_),
    .Y(_17697_));
 sky130_fd_sc_hd__o2bb2ai_2 _39761_ (.A1_N(_17687_),
    .A2_N(_17692_),
    .B1(_17695_),
    .B2(_17697_),
    .Y(_17698_));
 sky130_fd_sc_hd__nor2_2 _39762_ (.A(_17695_),
    .B(_17697_),
    .Y(_17699_));
 sky130_fd_sc_hd__nand3_2 _39763_ (.A(_17692_),
    .B(_17687_),
    .C(_17699_),
    .Y(_17700_));
 sky130_fd_sc_hd__nand3b_2 _39764_ (.A_N(_17601_),
    .B(_17698_),
    .C(_17700_),
    .Y(_17701_));
 sky130_fd_sc_hd__nor2_2 _39765_ (.A(_15729_),
    .B(_17696_),
    .Y(_17702_));
 sky130_fd_sc_hd__nor2_2 _39766_ (.A(_17165_),
    .B(_17694_),
    .Y(_17703_));
 sky130_fd_sc_hd__o2bb2ai_2 _39767_ (.A1_N(_17687_),
    .A2_N(_17692_),
    .B1(_17702_),
    .B2(_17703_),
    .Y(_17704_));
 sky130_fd_sc_hd__nand3b_2 _39768_ (.A_N(_17699_),
    .B(_17692_),
    .C(_17687_),
    .Y(_17705_));
 sky130_fd_sc_hd__nand3_2 _39769_ (.A(_17704_),
    .B(_17601_),
    .C(_17705_),
    .Y(_17706_));
 sky130_fd_sc_hd__a21oi_2 _39770_ (.A1(_17701_),
    .A2(_17706_),
    .B1(_17578_),
    .Y(_17707_));
 sky130_fd_sc_hd__and3_2 _39771_ (.A(_17701_),
    .B(_17706_),
    .C(_17578_),
    .X(_17708_));
 sky130_fd_sc_hd__nand3_2 _39772_ (.A(_17585_),
    .B(_17590_),
    .C(_17450_),
    .Y(_17709_));
 sky130_fd_sc_hd__nand2_2 _39773_ (.A(_17709_),
    .B(_17590_),
    .Y(_17710_));
 sky130_fd_sc_hd__o21bai_2 _39774_ (.A1(_17707_),
    .A2(_17708_),
    .B1_N(_17710_),
    .Y(_17711_));
 sky130_fd_sc_hd__nand3_2 _39775_ (.A(_17701_),
    .B(_17706_),
    .C(_17578_),
    .Y(_17712_));
 sky130_fd_sc_hd__nand3b_2 _39776_ (.A_N(_17707_),
    .B(_17710_),
    .C(_17712_),
    .Y(_17713_));
 sky130_fd_sc_hd__nand2_2 _39777_ (.A(_17711_),
    .B(_17713_),
    .Y(_17714_));
 sky130_fd_sc_hd__nand2_2 _39778_ (.A(_17594_),
    .B(_17709_),
    .Y(_17715_));
 sky130_fd_sc_hd__o2111a_2 _39779_ (.A1(_17596_),
    .A2(_17715_),
    .B1(_17469_),
    .C1(_17464_),
    .D1(_17597_),
    .X(_17716_));
 sky130_fd_sc_hd__nand3_2 _39780_ (.A(_17716_),
    .B(_17334_),
    .C(_17187_),
    .Y(_17717_));
 sky130_fd_sc_hd__o2111ai_2 _39781_ (.A1(_17596_),
    .A2(_17715_),
    .B1(_17469_),
    .C1(_17464_),
    .D1(_17597_),
    .Y(_17718_));
 sky130_fd_sc_hd__a21oi_2 _39782_ (.A1(_17592_),
    .A2(_17709_),
    .B1(_17594_),
    .Y(_17719_));
 sky130_fd_sc_hd__o22ai_2 _39783_ (.A1(_17591_),
    .A2(_17595_),
    .B1(_17469_),
    .B2(_17719_),
    .Y(_17720_));
 sky130_fd_sc_hd__o21bai_2 _39784_ (.A1(_17718_),
    .A2(_17476_),
    .B1_N(_17720_),
    .Y(_17721_));
 sky130_fd_sc_hd__o21bai_2 _39785_ (.A1(_17717_),
    .A2(_17472_),
    .B1_N(_17721_),
    .Y(_17722_));
 sky130_fd_sc_hd__xnor2_2 _39786_ (.A(_17714_),
    .B(_17722_),
    .Y(_02679_));
 sky130_fd_sc_hd__nand2_2 _39787_ (.A(_17722_),
    .B(_17711_),
    .Y(_17723_));
 sky130_fd_sc_hd__nand2_2 _39788_ (.A(_17694_),
    .B(_17165_),
    .Y(_17724_));
 sky130_fd_sc_hd__nand2_2 _39789_ (.A(_17669_),
    .B(_17666_),
    .Y(_17725_));
 sky130_fd_sc_hd__or2_2 _39790_ (.A(_17678_),
    .B(_17725_),
    .X(_17726_));
 sky130_fd_sc_hd__nand2_2 _39791_ (.A(_17725_),
    .B(_17678_),
    .Y(_17727_));
 sky130_fd_sc_hd__nand2_2 _39792_ (.A(_17726_),
    .B(_17727_),
    .Y(_17728_));
 sky130_fd_sc_hd__nor2_2 _39793_ (.A(_17147_),
    .B(_17728_),
    .Y(_17729_));
 sky130_fd_sc_hd__nor2_2 _39794_ (.A(_17678_),
    .B(_17725_),
    .Y(_17730_));
 sky130_fd_sc_hd__inv_2 _39795_ (.A(_17727_),
    .Y(_17731_));
 sky130_fd_sc_hd__o21ai_2 _39796_ (.A1(_17730_),
    .A2(_17731_),
    .B1(_17147_),
    .Y(_17732_));
 sky130_fd_sc_hd__inv_2 _39797_ (.A(_17732_),
    .Y(_17733_));
 sky130_fd_sc_hd__a21oi_2 _39798_ (.A1(_17642_),
    .A2(_17651_),
    .B1(_17648_),
    .Y(_17734_));
 sky130_fd_sc_hd__nor2_2 _39799_ (.A(_17408_),
    .B(_17734_),
    .Y(_17735_));
 sky130_fd_sc_hd__nand2_2 _39800_ (.A(_17734_),
    .B(_17408_),
    .Y(_17736_));
 sky130_fd_sc_hd__nand2_2 _39801_ (.A(_17736_),
    .B(_17286_),
    .Y(_17737_));
 sky130_fd_sc_hd__nor2_2 _39802_ (.A(_17735_),
    .B(_17737_),
    .Y(_17738_));
 sky130_fd_sc_hd__inv_2 _39803_ (.A(_17736_),
    .Y(_17739_));
 sky130_fd_sc_hd__o21ai_2 _39804_ (.A1(_17735_),
    .A2(_17739_),
    .B1(_17135_),
    .Y(_17740_));
 sky130_fd_sc_hd__inv_2 _39805_ (.A(_17740_),
    .Y(_17741_));
 sky130_fd_sc_hd__and2_2 _39806_ (.A(_17614_),
    .B(_17611_),
    .X(_17742_));
 sky130_fd_sc_hd__nand2_2 _39807_ (.A(_19314_),
    .B(_19543_),
    .Y(_17743_));
 sky130_fd_sc_hd__or4_2 _39808_ (.A(_19551_),
    .B(_18184_),
    .C(_17048_),
    .D(_11764_),
    .X(_17744_));
 sky130_fd_sc_hd__a22o_2 _39809_ (.A1(_19310_),
    .A2(_19547_),
    .B1(_11036_),
    .B2(_11124_),
    .X(_17745_));
 sky130_fd_sc_hd__nand2_2 _39810_ (.A(_17744_),
    .B(_17745_),
    .Y(_17746_));
 sky130_fd_sc_hd__or2_2 _39811_ (.A(_17743_),
    .B(_17746_),
    .X(_17747_));
 sky130_fd_sc_hd__nand2_2 _39812_ (.A(_17746_),
    .B(_17743_),
    .Y(_17748_));
 sky130_fd_sc_hd__nand2_2 _39813_ (.A(_17747_),
    .B(_17748_),
    .Y(_17749_));
 sky130_fd_sc_hd__nand2_2 _39814_ (.A(_17742_),
    .B(_17749_),
    .Y(_17750_));
 sky130_fd_sc_hd__a21o_2 _39815_ (.A1(_17611_),
    .A2(_17614_),
    .B1(_17749_),
    .X(_17751_));
 sky130_fd_sc_hd__nand2_2 _39816_ (.A(_17750_),
    .B(_17751_),
    .Y(_17752_));
 sky130_fd_sc_hd__o21ai_2 _39817_ (.A1(_19318_),
    .A2(_19321_),
    .B1(_18158_),
    .Y(_17753_));
 sky130_fd_sc_hd__and3_2 _39818_ (.A(_18157_),
    .B(_19317_),
    .C(_19321_),
    .X(_17754_));
 sky130_fd_sc_hd__or2_2 _39819_ (.A(_17753_),
    .B(_17754_),
    .X(_17755_));
 sky130_fd_sc_hd__nor2_2 _39820_ (.A(_09358_),
    .B(_17755_),
    .Y(_17756_));
 sky130_fd_sc_hd__and2_2 _39821_ (.A(_17755_),
    .B(_17501_),
    .X(_17757_));
 sky130_fd_sc_hd__nor2_2 _39822_ (.A(_17756_),
    .B(_17757_),
    .Y(_17758_));
 sky130_fd_sc_hd__nand2_2 _39823_ (.A(_17752_),
    .B(_17758_),
    .Y(_17759_));
 sky130_fd_sc_hd__inv_2 _39824_ (.A(_17758_),
    .Y(_17760_));
 sky130_fd_sc_hd__nand3_2 _39825_ (.A(_17750_),
    .B(_17751_),
    .C(_17760_),
    .Y(_17761_));
 sky130_fd_sc_hd__a21boi_2 _39826_ (.A1(_17617_),
    .A2(_17622_),
    .B1_N(_17618_),
    .Y(_17762_));
 sky130_fd_sc_hd__a21o_2 _39827_ (.A1(_17759_),
    .A2(_17761_),
    .B1(_17762_),
    .X(_17763_));
 sky130_fd_sc_hd__nand3_2 _39828_ (.A(_17759_),
    .B(_17762_),
    .C(_17761_),
    .Y(_17764_));
 sky130_fd_sc_hd__o21bai_2 _39829_ (.A1(_17501_),
    .A2(_17605_),
    .B1_N(_17606_),
    .Y(_17765_));
 sky130_fd_sc_hd__or2_2 _39830_ (.A(_17765_),
    .B(_17518_),
    .X(_17766_));
 sky130_fd_sc_hd__nand2_2 _39831_ (.A(_17518_),
    .B(_17765_),
    .Y(_17767_));
 sky130_fd_sc_hd__nand2_2 _39832_ (.A(_17766_),
    .B(_17767_),
    .Y(_17768_));
 sky130_fd_sc_hd__nor2_2 _39833_ (.A(_17522_),
    .B(_17768_),
    .Y(_17769_));
 sky130_fd_sc_hd__and2_2 _39834_ (.A(_17768_),
    .B(_17514_),
    .X(_17770_));
 sky130_fd_sc_hd__nor2_2 _39835_ (.A(_17769_),
    .B(_17770_),
    .Y(_17771_));
 sky130_fd_sc_hd__a21o_2 _39836_ (.A1(_17763_),
    .A2(_17764_),
    .B1(_17771_),
    .X(_17772_));
 sky130_fd_sc_hd__nand3_2 _39837_ (.A(_17763_),
    .B(_17764_),
    .C(_17771_),
    .Y(_17773_));
 sky130_fd_sc_hd__a21oi_2 _39838_ (.A1(_17620_),
    .A2(_17623_),
    .B1(_17625_),
    .Y(_17774_));
 sky130_fd_sc_hd__a21o_2 _39839_ (.A1(_17634_),
    .A2(_17627_),
    .B1(_17774_),
    .X(_17775_));
 sky130_fd_sc_hd__a21oi_2 _39840_ (.A1(_17772_),
    .A2(_17773_),
    .B1(_17775_),
    .Y(_17776_));
 sky130_fd_sc_hd__and3_2 _39841_ (.A(_17775_),
    .B(_17772_),
    .C(_17773_),
    .X(_17777_));
 sky130_fd_sc_hd__a21o_2 _39842_ (.A1(_17632_),
    .A2(_17630_),
    .B1(_17644_),
    .X(_17778_));
 sky130_fd_sc_hd__nand3_2 _39843_ (.A(_17632_),
    .B(_17644_),
    .C(_17630_),
    .Y(_17779_));
 sky130_fd_sc_hd__nand2_2 _39844_ (.A(_17778_),
    .B(_17779_),
    .Y(_17780_));
 sky130_fd_sc_hd__nand2_2 _39845_ (.A(_17780_),
    .B(_17263_),
    .Y(_17781_));
 sky130_fd_sc_hd__nand3_2 _39846_ (.A(_17778_),
    .B(_17651_),
    .C(_17779_),
    .Y(_17782_));
 sky130_fd_sc_hd__nand2_2 _39847_ (.A(_17781_),
    .B(_17782_),
    .Y(_17783_));
 sky130_fd_sc_hd__o21ai_2 _39848_ (.A1(_17776_),
    .A2(_17777_),
    .B1(_17783_),
    .Y(_17784_));
 sky130_fd_sc_hd__a21o_2 _39849_ (.A1(_17772_),
    .A2(_17773_),
    .B1(_17775_),
    .X(_17785_));
 sky130_fd_sc_hd__nand3_2 _39850_ (.A(_17775_),
    .B(_17772_),
    .C(_17773_),
    .Y(_17786_));
 sky130_fd_sc_hd__nand3b_2 _39851_ (.A_N(_17783_),
    .B(_17785_),
    .C(_17786_),
    .Y(_17787_));
 sky130_fd_sc_hd__nand2_2 _39852_ (.A(_17641_),
    .B(_17659_),
    .Y(_17788_));
 sky130_fd_sc_hd__nand2_2 _39853_ (.A(_17788_),
    .B(_17637_),
    .Y(_17789_));
 sky130_fd_sc_hd__a21oi_2 _39854_ (.A1(_17784_),
    .A2(_17787_),
    .B1(_17789_),
    .Y(_17790_));
 sky130_fd_sc_hd__a21oi_2 _39855_ (.A1(_17639_),
    .A2(_17640_),
    .B1(_17603_),
    .Y(_17791_));
 sky130_fd_sc_hd__a31oi_2 _39856_ (.A1(_17639_),
    .A2(_17640_),
    .A3(_17603_),
    .B1(_17653_),
    .Y(_17792_));
 sky130_fd_sc_hd__o211a_2 _39857_ (.A1(_17791_),
    .A2(_17792_),
    .B1(_17787_),
    .C1(_17784_),
    .X(_17793_));
 sky130_fd_sc_hd__o22ai_2 _39858_ (.A1(_17738_),
    .A2(_17741_),
    .B1(_17790_),
    .B2(_17793_),
    .Y(_17794_));
 sky130_fd_sc_hd__inv_2 _39859_ (.A(_17787_),
    .Y(_17795_));
 sky130_fd_sc_hd__nand2_2 _39860_ (.A(_17784_),
    .B(_17789_),
    .Y(_17796_));
 sky130_fd_sc_hd__o21a_2 _39861_ (.A1(_17735_),
    .A2(_17737_),
    .B1(_17740_),
    .X(_17797_));
 sky130_fd_sc_hd__a21o_2 _39862_ (.A1(_17784_),
    .A2(_17787_),
    .B1(_17789_),
    .X(_17798_));
 sky130_fd_sc_hd__o211ai_2 _39863_ (.A1(_17795_),
    .A2(_17796_),
    .B1(_17797_),
    .C1(_17798_),
    .Y(_17799_));
 sky130_fd_sc_hd__nand2_2 _39864_ (.A(_17672_),
    .B(_17662_),
    .Y(_17800_));
 sky130_fd_sc_hd__a21oi_2 _39865_ (.A1(_17794_),
    .A2(_17799_),
    .B1(_17800_),
    .Y(_17801_));
 sky130_fd_sc_hd__nand2_2 _39866_ (.A(_17798_),
    .B(_17797_),
    .Y(_17802_));
 sky130_fd_sc_hd__o211a_2 _39867_ (.A1(_17793_),
    .A2(_17802_),
    .B1(_17794_),
    .C1(_17800_),
    .X(_17803_));
 sky130_fd_sc_hd__o22ai_2 _39868_ (.A1(_17729_),
    .A2(_17733_),
    .B1(_17801_),
    .B2(_17803_),
    .Y(_17804_));
 sky130_fd_sc_hd__a21o_2 _39869_ (.A1(_17794_),
    .A2(_17799_),
    .B1(_17800_),
    .X(_17805_));
 sky130_fd_sc_hd__nand2_2 _39870_ (.A(_17726_),
    .B(_17484_),
    .Y(_17806_));
 sky130_fd_sc_hd__o21a_2 _39871_ (.A1(_17731_),
    .A2(_17806_),
    .B1(_17732_),
    .X(_17807_));
 sky130_fd_sc_hd__nand3_2 _39872_ (.A(_17800_),
    .B(_17794_),
    .C(_17799_),
    .Y(_17808_));
 sky130_fd_sc_hd__nand3_2 _39873_ (.A(_17805_),
    .B(_17807_),
    .C(_17808_),
    .Y(_17809_));
 sky130_fd_sc_hd__o21ai_2 _39874_ (.A1(_17689_),
    .A2(_17690_),
    .B1(_17675_),
    .Y(_17810_));
 sky130_fd_sc_hd__a21oi_2 _39875_ (.A1(_17804_),
    .A2(_17809_),
    .B1(_17810_),
    .Y(_17811_));
 sky130_fd_sc_hd__a21oi_2 _39876_ (.A1(_17805_),
    .A2(_17808_),
    .B1(_17807_),
    .Y(_17812_));
 sky130_fd_sc_hd__nand2_2 _39877_ (.A(_17810_),
    .B(_17809_),
    .Y(_17813_));
 sky130_fd_sc_hd__nor2_2 _39878_ (.A(_17812_),
    .B(_17813_),
    .Y(_17814_));
 sky130_fd_sc_hd__nand2_2 _39879_ (.A(_17681_),
    .B(_17679_),
    .Y(_17815_));
 sky130_fd_sc_hd__nor2_2 _39880_ (.A(_17164_),
    .B(_17815_),
    .Y(_17816_));
 sky130_fd_sc_hd__nand2_2 _39881_ (.A(_17815_),
    .B(_17164_),
    .Y(_17817_));
 sky130_fd_sc_hd__or2b_2 _39882_ (.A(_17816_),
    .B_N(_17817_),
    .X(_17818_));
 sky130_fd_sc_hd__o21ai_2 _39883_ (.A1(_17811_),
    .A2(_17814_),
    .B1(_17818_),
    .Y(_17819_));
 sky130_fd_sc_hd__nor2b_2 _39884_ (.A(_17816_),
    .B_N(_17817_),
    .Y(_17820_));
 sky130_fd_sc_hd__a21o_2 _39885_ (.A1(_17804_),
    .A2(_17809_),
    .B1(_17810_),
    .X(_17821_));
 sky130_fd_sc_hd__o211ai_2 _39886_ (.A1(_17812_),
    .A2(_17813_),
    .B1(_17820_),
    .C1(_17821_),
    .Y(_17822_));
 sky130_fd_sc_hd__a21oi_2 _39887_ (.A1(_17684_),
    .A2(_17686_),
    .B1(_17685_),
    .Y(_17823_));
 sky130_fd_sc_hd__o21ai_2 _39888_ (.A1(_17699_),
    .A2(_17823_),
    .B1(_17687_),
    .Y(_17824_));
 sky130_fd_sc_hd__a21oi_2 _39889_ (.A1(_17819_),
    .A2(_17822_),
    .B1(_17824_),
    .Y(_17825_));
 sky130_fd_sc_hd__nand2_2 _39890_ (.A(_17821_),
    .B(_17820_),
    .Y(_17826_));
 sky130_fd_sc_hd__o211a_2 _39891_ (.A1(_17814_),
    .A2(_17826_),
    .B1(_17819_),
    .C1(_17824_),
    .X(_17827_));
 sky130_fd_sc_hd__nor3_2 _39892_ (.A(_17724_),
    .B(_17825_),
    .C(_17827_),
    .Y(_17828_));
 sky130_fd_sc_hd__o22a_2 _39893_ (.A1(_17180_),
    .A2(_17696_),
    .B1(_17825_),
    .B2(_17827_),
    .X(_17829_));
 sky130_fd_sc_hd__a211o_2 _39894_ (.A1(_17706_),
    .A2(_17712_),
    .B1(_17828_),
    .C1(_17829_),
    .X(_17830_));
 sky130_fd_sc_hd__nand2_2 _39895_ (.A(_17712_),
    .B(_17706_),
    .Y(_17831_));
 sky130_fd_sc_hd__o21bai_2 _39896_ (.A1(_17828_),
    .A2(_17829_),
    .B1_N(_17831_),
    .Y(_17832_));
 sky130_fd_sc_hd__nand2_2 _39897_ (.A(_17830_),
    .B(_17832_),
    .Y(_17833_));
 sky130_fd_sc_hd__a21bo_2 _39898_ (.A1(_17723_),
    .A2(_17713_),
    .B1_N(_17833_),
    .X(_17834_));
 sky130_fd_sc_hd__nand3b_2 _39899_ (.A_N(_17833_),
    .B(_17723_),
    .C(_17713_),
    .Y(_17835_));
 sky130_fd_sc_hd__nand2_2 _39900_ (.A(_17834_),
    .B(_17835_),
    .Y(_02680_));
 sky130_fd_sc_hd__o21bai_2 _39901_ (.A1(_17825_),
    .A2(_17827_),
    .B1_N(_17702_),
    .Y(_17836_));
 sky130_fd_sc_hd__nand2_2 _39902_ (.A(_17836_),
    .B(_17831_),
    .Y(_17837_));
 sky130_fd_sc_hd__o2111a_2 _39903_ (.A1(_17828_),
    .A2(_17837_),
    .B1(_17711_),
    .C1(_17713_),
    .D1(_17832_),
    .X(_17838_));
 sky130_fd_sc_hd__nand2_2 _39904_ (.A(_17722_),
    .B(_17838_),
    .Y(_17839_));
 sky130_fd_sc_hd__a21bo_2 _39905_ (.A1(_17830_),
    .A2(_17713_),
    .B1_N(_17832_),
    .X(_17840_));
 sky130_fd_sc_hd__nand2_2 _39906_ (.A(_18158_),
    .B(_19314_),
    .Y(_17841_));
 sky130_fd_sc_hd__or4_2 _39907_ (.A(_19547_),
    .B(_18184_),
    .C(_17048_),
    .D(_15116_),
    .X(_17842_));
 sky130_fd_sc_hd__a22o_2 _39908_ (.A1(_19310_),
    .A2(_19542_),
    .B1(_11764_),
    .B2(_11124_),
    .X(_17843_));
 sky130_fd_sc_hd__nand2_2 _39909_ (.A(_17842_),
    .B(_17843_),
    .Y(_17844_));
 sky130_fd_sc_hd__or2_2 _39910_ (.A(_17841_),
    .B(_17844_),
    .X(_17845_));
 sky130_fd_sc_hd__nand2_2 _39911_ (.A(_17844_),
    .B(_17841_),
    .Y(_17846_));
 sky130_fd_sc_hd__nand2_2 _39912_ (.A(_17845_),
    .B(_17846_),
    .Y(_17847_));
 sky130_fd_sc_hd__a21o_2 _39913_ (.A1(_17744_),
    .A2(_17747_),
    .B1(_17847_),
    .X(_17848_));
 sky130_fd_sc_hd__nand3_2 _39914_ (.A(_17847_),
    .B(_17744_),
    .C(_17747_),
    .Y(_17849_));
 sky130_fd_sc_hd__nand2_2 _39915_ (.A(_17848_),
    .B(_17849_),
    .Y(_17850_));
 sky130_fd_sc_hd__nand2_2 _39916_ (.A(_17850_),
    .B(_17758_),
    .Y(_17851_));
 sky130_fd_sc_hd__nand3_2 _39917_ (.A(_17848_),
    .B(_17760_),
    .C(_17849_),
    .Y(_17852_));
 sky130_fd_sc_hd__nor2_2 _39918_ (.A(_17749_),
    .B(_17742_),
    .Y(_17853_));
 sky130_fd_sc_hd__a21oi_2 _39919_ (.A1(_17750_),
    .A2(_17758_),
    .B1(_17853_),
    .Y(_17854_));
 sky130_fd_sc_hd__a21oi_2 _39920_ (.A1(_17851_),
    .A2(_17852_),
    .B1(_17854_),
    .Y(_17855_));
 sky130_fd_sc_hd__and3_2 _39921_ (.A(_17851_),
    .B(_17854_),
    .C(_17852_),
    .X(_17856_));
 sky130_fd_sc_hd__nor2_2 _39922_ (.A(_17855_),
    .B(_17856_),
    .Y(_17857_));
 sky130_fd_sc_hd__or2_2 _39923_ (.A(_17754_),
    .B(_17756_),
    .X(_17858_));
 sky130_fd_sc_hd__or2_2 _39924_ (.A(_17858_),
    .B(_17516_),
    .X(_17859_));
 sky130_fd_sc_hd__nand2_2 _39925_ (.A(_17518_),
    .B(_17858_),
    .Y(_17860_));
 sky130_fd_sc_hd__nand2_2 _39926_ (.A(_17859_),
    .B(_17860_),
    .Y(_17861_));
 sky130_fd_sc_hd__nor2_2 _39927_ (.A(_17522_),
    .B(_17861_),
    .Y(_17862_));
 sky130_fd_sc_hd__and2_2 _39928_ (.A(_17861_),
    .B(_17514_),
    .X(_17863_));
 sky130_fd_sc_hd__nor2_2 _39929_ (.A(_17862_),
    .B(_17863_),
    .Y(_17864_));
 sky130_fd_sc_hd__inv_2 _39930_ (.A(_17864_),
    .Y(_17865_));
 sky130_fd_sc_hd__nand2_2 _39931_ (.A(_17857_),
    .B(_17865_),
    .Y(_17866_));
 sky130_fd_sc_hd__a21boi_2 _39932_ (.A1(_17764_),
    .A2(_17771_),
    .B1_N(_17763_),
    .Y(_17867_));
 sky130_fd_sc_hd__o21ai_2 _39933_ (.A1(_17855_),
    .A2(_17856_),
    .B1(_17864_),
    .Y(_17868_));
 sky130_fd_sc_hd__nand3_2 _39934_ (.A(_17866_),
    .B(_17867_),
    .C(_17868_),
    .Y(_17869_));
 sky130_fd_sc_hd__nand2_2 _39935_ (.A(_17857_),
    .B(_17864_),
    .Y(_17870_));
 sky130_fd_sc_hd__nand2_2 _39936_ (.A(_17773_),
    .B(_17763_),
    .Y(_17871_));
 sky130_fd_sc_hd__o21ai_2 _39937_ (.A1(_17855_),
    .A2(_17856_),
    .B1(_17865_),
    .Y(_17872_));
 sky130_fd_sc_hd__nand3_2 _39938_ (.A(_17870_),
    .B(_17871_),
    .C(_17872_),
    .Y(_17873_));
 sky130_fd_sc_hd__o21ai_2 _39939_ (.A1(_17522_),
    .A2(_17768_),
    .B1(_17767_),
    .Y(_17874_));
 sky130_fd_sc_hd__and2_2 _39940_ (.A(_17874_),
    .B(_17537_),
    .X(_17875_));
 sky130_fd_sc_hd__nor2_2 _39941_ (.A(_17537_),
    .B(_17874_),
    .Y(_17876_));
 sky130_fd_sc_hd__o2bb2ai_2 _39942_ (.A1_N(_17869_),
    .A2_N(_17873_),
    .B1(_17875_),
    .B2(_17876_),
    .Y(_17877_));
 sky130_fd_sc_hd__nor2_2 _39943_ (.A(_17876_),
    .B(_17875_),
    .Y(_17878_));
 sky130_fd_sc_hd__nand3_2 _39944_ (.A(_17873_),
    .B(_17869_),
    .C(_17878_),
    .Y(_17879_));
 sky130_fd_sc_hd__o21ai_2 _39945_ (.A1(_17783_),
    .A2(_17776_),
    .B1(_17786_),
    .Y(_17880_));
 sky130_fd_sc_hd__a21o_2 _39946_ (.A1(_17877_),
    .A2(_17879_),
    .B1(_17880_),
    .X(_17881_));
 sky130_fd_sc_hd__nand3_2 _39947_ (.A(_17880_),
    .B(_17877_),
    .C(_17879_),
    .Y(_17882_));
 sky130_fd_sc_hd__a21oi_2 _39948_ (.A1(_17632_),
    .A2(_17630_),
    .B1(_17644_),
    .Y(_17883_));
 sky130_fd_sc_hd__a211o_2 _39949_ (.A1(_17779_),
    .A2(_17651_),
    .B1(_16899_),
    .C1(_17883_),
    .X(_17884_));
 sky130_fd_sc_hd__nand2_2 _39950_ (.A(_17782_),
    .B(_17778_),
    .Y(_17885_));
 sky130_fd_sc_hd__a22oi_2 _39951_ (.A1(_17884_),
    .A2(_15586_),
    .B1(_16730_),
    .B2(_17885_),
    .Y(_17886_));
 sky130_fd_sc_hd__a211o_2 _39952_ (.A1(_17779_),
    .A2(_17651_),
    .B1(_16730_),
    .C1(_17883_),
    .X(_17887_));
 sky130_fd_sc_hd__nand2_2 _39953_ (.A(_17885_),
    .B(_16730_),
    .Y(_17888_));
 sky130_fd_sc_hd__nand2_2 _39954_ (.A(_17888_),
    .B(_17887_),
    .Y(_17889_));
 sky130_fd_sc_hd__a22o_2 _39955_ (.A1(_17886_),
    .A2(_17887_),
    .B1(_16733_),
    .B2(_17889_),
    .X(_17890_));
 sky130_fd_sc_hd__a21oi_2 _39956_ (.A1(_17881_),
    .A2(_17882_),
    .B1(_17890_),
    .Y(_17891_));
 sky130_fd_sc_hd__and3_2 _39957_ (.A(_17881_),
    .B(_17882_),
    .C(_17890_),
    .X(_17892_));
 sky130_fd_sc_hd__o21ai_2 _39958_ (.A1(_17735_),
    .A2(_17737_),
    .B1(_17740_),
    .Y(_17893_));
 sky130_fd_sc_hd__o22ai_2 _39959_ (.A1(_17795_),
    .A2(_17796_),
    .B1(_17893_),
    .B2(_17790_),
    .Y(_17894_));
 sky130_fd_sc_hd__o21bai_2 _39960_ (.A1(_17891_),
    .A2(_17892_),
    .B1_N(_17894_),
    .Y(_17895_));
 sky130_fd_sc_hd__nand3_2 _39961_ (.A(_17881_),
    .B(_17882_),
    .C(_17890_),
    .Y(_17896_));
 sky130_fd_sc_hd__nand3b_2 _39962_ (.A_N(_17891_),
    .B(_17896_),
    .C(_17894_),
    .Y(_17897_));
 sky130_fd_sc_hd__o21ai_2 _39963_ (.A1(_17408_),
    .A2(_17734_),
    .B1(_17737_),
    .Y(_17898_));
 sky130_fd_sc_hd__or2_2 _39964_ (.A(_17678_),
    .B(_17898_),
    .X(_17899_));
 sky130_fd_sc_hd__nand2_2 _39965_ (.A(_17898_),
    .B(_17678_),
    .Y(_17900_));
 sky130_fd_sc_hd__a21oi_2 _39966_ (.A1(_17899_),
    .A2(_17900_),
    .B1(_17147_),
    .Y(_17901_));
 sky130_fd_sc_hd__nand3_2 _39967_ (.A(_17899_),
    .B(_17147_),
    .C(_17900_),
    .Y(_17902_));
 sky130_fd_sc_hd__or2b_2 _39968_ (.A(_17901_),
    .B_N(_17902_),
    .X(_17903_));
 sky130_fd_sc_hd__a21o_2 _39969_ (.A1(_17895_),
    .A2(_17897_),
    .B1(_17903_),
    .X(_17904_));
 sky130_fd_sc_hd__nand3_2 _39970_ (.A(_17903_),
    .B(_17895_),
    .C(_17897_),
    .Y(_17905_));
 sky130_fd_sc_hd__o21ai_2 _39971_ (.A1(_17731_),
    .A2(_17806_),
    .B1(_17732_),
    .Y(_17906_));
 sky130_fd_sc_hd__o21ai_2 _39972_ (.A1(_17906_),
    .A2(_17801_),
    .B1(_17808_),
    .Y(_17907_));
 sky130_fd_sc_hd__nand3_2 _39973_ (.A(_17904_),
    .B(_17905_),
    .C(_17907_),
    .Y(_17908_));
 sky130_fd_sc_hd__a21oi_2 _39974_ (.A1(_17895_),
    .A2(_17897_),
    .B1(_17903_),
    .Y(_17909_));
 sky130_fd_sc_hd__inv_2 _39975_ (.A(_17902_),
    .Y(_17910_));
 sky130_fd_sc_hd__o211a_2 _39976_ (.A1(_17901_),
    .A2(_17910_),
    .B1(_17897_),
    .C1(_17895_),
    .X(_17911_));
 sky130_fd_sc_hd__o21bai_2 _39977_ (.A1(_17909_),
    .A2(_17911_),
    .B1_N(_17907_),
    .Y(_17912_));
 sky130_fd_sc_hd__nand2_2 _39978_ (.A(_17806_),
    .B(_17727_),
    .Y(_17913_));
 sky130_fd_sc_hd__nor2_2 _39979_ (.A(_17165_),
    .B(_17913_),
    .Y(_17914_));
 sky130_fd_sc_hd__and2_2 _39980_ (.A(_17913_),
    .B(_17164_),
    .X(_17915_));
 sky130_fd_sc_hd__o2bb2ai_2 _39981_ (.A1_N(_17908_),
    .A2_N(_17912_),
    .B1(_17914_),
    .B2(_17915_),
    .Y(_17916_));
 sky130_fd_sc_hd__nor2_2 _39982_ (.A(_17914_),
    .B(_17915_),
    .Y(_17917_));
 sky130_fd_sc_hd__nand3_2 _39983_ (.A(_17912_),
    .B(_17908_),
    .C(_17917_),
    .Y(_17918_));
 sky130_fd_sc_hd__buf_1 _39984_ (.A(_17918_),
    .X(_17919_));
 sky130_fd_sc_hd__nor2_2 _39985_ (.A(_17820_),
    .B(_17814_),
    .Y(_17920_));
 sky130_fd_sc_hd__o2bb2ai_2 _39986_ (.A1_N(_17916_),
    .A2_N(_17919_),
    .B1(_17811_),
    .B2(_17920_),
    .Y(_17921_));
 sky130_fd_sc_hd__o22ai_2 _39987_ (.A1(_17812_),
    .A2(_17813_),
    .B1(_17818_),
    .B2(_17811_),
    .Y(_17922_));
 sky130_fd_sc_hd__nand3_2 _39988_ (.A(_17916_),
    .B(_17922_),
    .C(_17918_),
    .Y(_17923_));
 sky130_fd_sc_hd__a22o_2 _39989_ (.A1(_17165_),
    .A2(_17815_),
    .B1(_17921_),
    .B2(_17923_),
    .X(_17924_));
 sky130_fd_sc_hd__nand2_2 _39990_ (.A(_17916_),
    .B(_17919_),
    .Y(_17925_));
 sky130_fd_sc_hd__a21oi_2 _39991_ (.A1(_17821_),
    .A2(_17820_),
    .B1(_17814_),
    .Y(_17926_));
 sky130_fd_sc_hd__a21oi_2 _39992_ (.A1(_17925_),
    .A2(_17926_),
    .B1(_17817_),
    .Y(_17927_));
 sky130_fd_sc_hd__nand2_2 _39993_ (.A(_17927_),
    .B(_17923_),
    .Y(_17928_));
 sky130_fd_sc_hd__nand2_2 _39994_ (.A(_17924_),
    .B(_17928_),
    .Y(_17929_));
 sky130_fd_sc_hd__nor2_2 _39995_ (.A(_17827_),
    .B(_17828_),
    .Y(_17930_));
 sky130_fd_sc_hd__or2_2 _39996_ (.A(_17929_),
    .B(_17930_),
    .X(_17931_));
 sky130_fd_sc_hd__nand2_2 _39997_ (.A(_17930_),
    .B(_17929_),
    .Y(_17932_));
 sky130_fd_sc_hd__nand2_2 _39998_ (.A(_17931_),
    .B(_17932_),
    .Y(_17933_));
 sky130_fd_sc_hd__a21bo_2 _39999_ (.A1(_17839_),
    .A2(_17840_),
    .B1_N(_17933_),
    .X(_17934_));
 sky130_fd_sc_hd__nand3b_2 _40000_ (.A_N(_17933_),
    .B(_17839_),
    .C(_17840_),
    .Y(_17935_));
 sky130_fd_sc_hd__nand2_2 _40001_ (.A(_17934_),
    .B(_17935_),
    .Y(_02681_));
 sky130_fd_sc_hd__a21oi_2 _40002_ (.A1(_17916_),
    .A2(_17919_),
    .B1(_17922_),
    .Y(_17936_));
 sky130_fd_sc_hd__o21a_2 _40003_ (.A1(_17108_),
    .A2(_17874_),
    .B1(_17107_),
    .X(_17937_));
 sky130_fd_sc_hd__nand2_2 _40004_ (.A(_18158_),
    .B(_19310_),
    .Y(_17938_));
 sky130_fd_sc_hd__xor2_2 _40005_ (.A(_17758_),
    .B(_17864_),
    .X(_17939_));
 sky130_fd_sc_hd__xor2_2 _40006_ (.A(_17841_),
    .B(_17939_),
    .X(_17940_));
 sky130_fd_sc_hd__xor2_2 _40007_ (.A(_17938_),
    .B(_17940_),
    .X(_17941_));
 sky130_fd_sc_hd__xnor2_2 _40008_ (.A(_17937_),
    .B(_17941_),
    .Y(_17942_));
 sky130_fd_sc_hd__inv_2 _40009_ (.A(_17942_),
    .Y(_17943_));
 sky130_fd_sc_hd__a31oi_2 _40010_ (.A1(_17916_),
    .A2(_17922_),
    .A3(_17919_),
    .B1(_17943_),
    .Y(_17944_));
 sky130_fd_sc_hd__o21ai_2 _40011_ (.A1(_17817_),
    .A2(_17936_),
    .B1(_17944_),
    .Y(_17945_));
 sky130_fd_sc_hd__nand2_2 _40012_ (.A(_17923_),
    .B(_17817_),
    .Y(_17946_));
 sky130_fd_sc_hd__nand3_2 _40013_ (.A(_17946_),
    .B(_17921_),
    .C(_17943_),
    .Y(_17947_));
 sky130_fd_sc_hd__nand2_2 _40014_ (.A(_16087_),
    .B(_14794_),
    .Y(_17948_));
 sky130_fd_sc_hd__o21a_2 _40015_ (.A1(_14794_),
    .A2(_15749_),
    .B1(_17948_),
    .X(_17949_));
 sky130_fd_sc_hd__inv_2 _40016_ (.A(_17949_),
    .Y(_17950_));
 sky130_fd_sc_hd__a21oi_2 _40017_ (.A1(_17945_),
    .A2(_17947_),
    .B1(_17950_),
    .Y(_17951_));
 sky130_fd_sc_hd__nand2_2 _40018_ (.A(_17923_),
    .B(_17942_),
    .Y(_17952_));
 sky130_fd_sc_hd__o211a_2 _40019_ (.A1(_17952_),
    .A2(_17927_),
    .B1(_17950_),
    .C1(_17947_),
    .X(_17953_));
 sky130_fd_sc_hd__and2_2 _40020_ (.A(_17879_),
    .B(_17873_),
    .X(_17954_));
 sky130_fd_sc_hd__nand2_2 _40021_ (.A(_17905_),
    .B(_17897_),
    .Y(_17955_));
 sky130_fd_sc_hd__or2_2 _40022_ (.A(_17954_),
    .B(_17955_),
    .X(_17956_));
 sky130_fd_sc_hd__nand2_2 _40023_ (.A(_17955_),
    .B(_17954_),
    .Y(_17957_));
 sky130_fd_sc_hd__o21a_2 _40024_ (.A1(_17522_),
    .A2(_17861_),
    .B1(_17860_),
    .X(_17958_));
 sky130_fd_sc_hd__a21oi_2 _40025_ (.A1(_17956_),
    .A2(_17957_),
    .B1(_17958_),
    .Y(_17959_));
 sky130_fd_sc_hd__and3_2 _40026_ (.A(_17956_),
    .B(_17957_),
    .C(_17958_),
    .X(_17960_));
 sky130_fd_sc_hd__nor2_2 _40027_ (.A(_17959_),
    .B(_17960_),
    .Y(_17961_));
 sky130_fd_sc_hd__o21ai_2 _40028_ (.A1(_17951_),
    .A2(_17953_),
    .B1(_17961_),
    .Y(_17962_));
 sky130_fd_sc_hd__nor2_2 _40029_ (.A(_17952_),
    .B(_17927_),
    .Y(_17963_));
 sky130_fd_sc_hd__nand2_2 _40030_ (.A(_17947_),
    .B(_17950_),
    .Y(_17964_));
 sky130_fd_sc_hd__nand2_2 _40031_ (.A(_17945_),
    .B(_17947_),
    .Y(_17965_));
 sky130_fd_sc_hd__nand2_2 _40032_ (.A(_17965_),
    .B(_17949_),
    .Y(_17966_));
 sky130_fd_sc_hd__o221ai_2 _40033_ (.A1(_17963_),
    .A2(_17964_),
    .B1(_17960_),
    .B2(_17959_),
    .C1(_17966_),
    .Y(_17967_));
 sky130_fd_sc_hd__o21ai_2 _40034_ (.A1(_17760_),
    .A2(_17850_),
    .B1(_17848_),
    .Y(_17968_));
 sky130_fd_sc_hd__xor2_2 _40035_ (.A(_17968_),
    .B(_17886_),
    .X(_17969_));
 sky130_fd_sc_hd__inv_2 _40036_ (.A(_17969_),
    .Y(_17970_));
 sky130_fd_sc_hd__a21o_2 _40037_ (.A1(_17919_),
    .A2(_17908_),
    .B1(_17970_),
    .X(_17971_));
 sky130_fd_sc_hd__nand3_2 _40038_ (.A(_17919_),
    .B(_17908_),
    .C(_17970_),
    .Y(_17972_));
 sky130_fd_sc_hd__a21bo_2 _40039_ (.A1(_17899_),
    .A2(_17484_),
    .B1_N(_17900_),
    .X(_17973_));
 sky130_fd_sc_hd__nor2_2 _40040_ (.A(_17180_),
    .B(_17913_),
    .Y(_17974_));
 sky130_fd_sc_hd__xor2_2 _40041_ (.A(_17973_),
    .B(_17974_),
    .X(_17975_));
 sky130_fd_sc_hd__a21o_2 _40042_ (.A1(_17971_),
    .A2(_17972_),
    .B1(_17975_),
    .X(_17976_));
 sky130_fd_sc_hd__nand3_2 _40043_ (.A(_17971_),
    .B(_17975_),
    .C(_17972_),
    .Y(_17977_));
 sky130_fd_sc_hd__nand2_2 _40044_ (.A(_15116_),
    .B(_11124_),
    .Y(_17978_));
 sky130_fd_sc_hd__nand2_2 _40045_ (.A(_17845_),
    .B(_17842_),
    .Y(_17979_));
 sky130_fd_sc_hd__xor2_2 _40046_ (.A(_17978_),
    .B(_17979_),
    .X(_17980_));
 sky130_fd_sc_hd__a21oi_2 _40047_ (.A1(_17857_),
    .A2(_17864_),
    .B1(_17855_),
    .Y(_17981_));
 sky130_fd_sc_hd__nand2_2 _40048_ (.A(_17896_),
    .B(_17882_),
    .Y(_17982_));
 sky130_fd_sc_hd__or2_2 _40049_ (.A(_17981_),
    .B(_17982_),
    .X(_17983_));
 sky130_fd_sc_hd__nand2_2 _40050_ (.A(_17982_),
    .B(_17981_),
    .Y(_17984_));
 sky130_fd_sc_hd__nand2_2 _40051_ (.A(_17983_),
    .B(_17984_),
    .Y(_17985_));
 sky130_fd_sc_hd__xor2_2 _40052_ (.A(_17980_),
    .B(_17985_),
    .X(_17986_));
 sky130_fd_sc_hd__a21o_2 _40053_ (.A1(_17976_),
    .A2(_17977_),
    .B1(_17986_),
    .X(_17987_));
 sky130_fd_sc_hd__nand3_2 _40054_ (.A(_17976_),
    .B(_17986_),
    .C(_17977_),
    .Y(_17988_));
 sky130_fd_sc_hd__nand2_2 _40055_ (.A(_17987_),
    .B(_17988_),
    .Y(_17989_));
 sky130_fd_sc_hd__a21oi_2 _40056_ (.A1(_17962_),
    .A2(_17967_),
    .B1(_17989_),
    .Y(_17990_));
 sky130_fd_sc_hd__a21oi_2 _40057_ (.A1(_17976_),
    .A2(_17977_),
    .B1(_17986_),
    .Y(_17991_));
 sky130_fd_sc_hd__inv_2 _40058_ (.A(_17988_),
    .Y(_17992_));
 sky130_fd_sc_hd__o211a_2 _40059_ (.A1(_17991_),
    .A2(_17992_),
    .B1(_17967_),
    .C1(_17962_),
    .X(_17993_));
 sky130_fd_sc_hd__o22ai_2 _40060_ (.A1(_17930_),
    .A2(_17929_),
    .B1(_17990_),
    .B2(_17993_),
    .Y(_17994_));
 sky130_fd_sc_hd__a21oi_2 _40061_ (.A1(_17839_),
    .A2(_17840_),
    .B1(_17933_),
    .Y(_17995_));
 sky130_fd_sc_hd__nand3_2 _40062_ (.A(_17839_),
    .B(_17931_),
    .C(_17840_),
    .Y(_17996_));
 sky130_fd_sc_hd__o2bb2ai_2 _40063_ (.A1_N(_17949_),
    .A2_N(_17965_),
    .B1(_17964_),
    .B2(_17963_),
    .Y(_17997_));
 sky130_fd_sc_hd__a22oi_2 _40064_ (.A1(_17987_),
    .A2(_17988_),
    .B1(_17997_),
    .B2(_17961_),
    .Y(_17998_));
 sky130_fd_sc_hd__nand2_2 _40065_ (.A(_17962_),
    .B(_17967_),
    .Y(_17999_));
 sky130_fd_sc_hd__inv_2 _40066_ (.A(_17989_),
    .Y(_18000_));
 sky130_fd_sc_hd__a22oi_2 _40067_ (.A1(_17998_),
    .A2(_17967_),
    .B1(_17999_),
    .B2(_18000_),
    .Y(_18001_));
 sky130_fd_sc_hd__nand3_2 _40068_ (.A(_17996_),
    .B(_17932_),
    .C(_18001_),
    .Y(_18002_));
 sky130_fd_sc_hd__o21ai_2 _40069_ (.A1(_17994_),
    .A2(_17995_),
    .B1(_18002_),
    .Y(_02682_));
 sky130_fd_sc_hd__xnor2_2 _40070_ (.A(_05314_),
    .B(_05178_),
    .Y(_02628_));
 sky130_fd_sc_hd__nor2_2 _40071_ (.A(_19790_),
    .B(_04846_),
    .Y(_00050_));
 sky130_fd_sc_hd__and3_2 _40072_ (.A(_02321_),
    .B(_02318_),
    .C(_00066_),
    .X(_00068_));
 sky130_fd_sc_hd__and2_2 _40073_ (.A(_02321_),
    .B(_00084_),
    .X(_00085_));
 sky130_fd_sc_hd__and2_2 _40074_ (.A(_02321_),
    .B(_00094_),
    .X(_00095_));
 sky130_fd_sc_hd__o21a_2 _40075_ (.A1(instr_sra),
    .A2(instr_srai),
    .B1(pcpi_rs1[31]),
    .X(_00216_));
 sky130_fd_sc_hd__o21a_2 _40076_ (.A1(_18240_),
    .A2(_18241_),
    .B1(_00321_),
    .X(_18003_));
 sky130_fd_sc_hd__nand2_2 _40077_ (.A(_18003_),
    .B(_18250_),
    .Y(_18004_));
 sky130_fd_sc_hd__o211a_2 _40078_ (.A1(irq_active),
    .A2(_18003_),
    .B1(_18660_),
    .C1(_18004_),
    .X(_04072_));
 sky130_fd_sc_hd__conb_1 _40079_ (.LO(mem_addr[0]));
 sky130_fd_sc_hd__conb_1 _40080_ (.LO(mem_addr[1]));
 sky130_fd_sc_hd__conb_1 _40081_ (.LO(mem_la_addr[0]));
 sky130_fd_sc_hd__conb_1 _40082_ (.LO(mem_la_addr[1]));
 sky130_fd_sc_hd__conb_1 _40083_ (.LO(trace_data[0]));
 sky130_fd_sc_hd__conb_1 _40084_ (.LO(trace_data[1]));
 sky130_fd_sc_hd__conb_1 _40085_ (.LO(trace_data[2]));
 sky130_fd_sc_hd__conb_1 _40086_ (.LO(trace_data[3]));
 sky130_fd_sc_hd__conb_1 _40087_ (.LO(trace_data[4]));
 sky130_fd_sc_hd__conb_1 _40088_ (.LO(trace_data[5]));
 sky130_fd_sc_hd__conb_1 _40089_ (.LO(trace_data[6]));
 sky130_fd_sc_hd__conb_1 _40090_ (.LO(trace_data[7]));
 sky130_fd_sc_hd__conb_1 _40091_ (.LO(trace_data[8]));
 sky130_fd_sc_hd__conb_1 _40092_ (.LO(trace_data[9]));
 sky130_fd_sc_hd__conb_1 _40093_ (.LO(trace_data[10]));
 sky130_fd_sc_hd__conb_1 _40094_ (.LO(trace_data[11]));
 sky130_fd_sc_hd__conb_1 _40095_ (.LO(trace_data[12]));
 sky130_fd_sc_hd__conb_1 _40096_ (.LO(trace_data[13]));
 sky130_fd_sc_hd__conb_1 _40097_ (.LO(trace_data[14]));
 sky130_fd_sc_hd__conb_1 _40098_ (.LO(trace_data[15]));
 sky130_fd_sc_hd__conb_1 _40099_ (.LO(trace_data[16]));
 sky130_fd_sc_hd__conb_1 _40100_ (.LO(trace_data[17]));
 sky130_fd_sc_hd__conb_1 _40101_ (.LO(trace_data[18]));
 sky130_fd_sc_hd__conb_1 _40102_ (.LO(trace_data[19]));
 sky130_fd_sc_hd__conb_1 _40103_ (.LO(trace_data[20]));
 sky130_fd_sc_hd__conb_1 _40104_ (.LO(trace_data[21]));
 sky130_fd_sc_hd__conb_1 _40105_ (.LO(trace_data[22]));
 sky130_fd_sc_hd__conb_1 _40106_ (.LO(trace_data[23]));
 sky130_fd_sc_hd__conb_1 _40107_ (.LO(trace_data[24]));
 sky130_fd_sc_hd__conb_1 _40108_ (.LO(trace_data[25]));
 sky130_fd_sc_hd__conb_1 _40109_ (.LO(trace_data[26]));
 sky130_fd_sc_hd__conb_1 _40110_ (.LO(trace_data[27]));
 sky130_fd_sc_hd__conb_1 _40111_ (.LO(trace_data[28]));
 sky130_fd_sc_hd__conb_1 _40112_ (.LO(trace_data[29]));
 sky130_fd_sc_hd__conb_1 _40113_ (.LO(trace_data[30]));
 sky130_fd_sc_hd__conb_1 _40114_ (.LO(trace_data[31]));
 sky130_fd_sc_hd__conb_1 _40115_ (.LO(trace_data[32]));
 sky130_fd_sc_hd__conb_1 _40116_ (.LO(trace_data[33]));
 sky130_fd_sc_hd__conb_1 _40117_ (.LO(trace_data[34]));
 sky130_fd_sc_hd__conb_1 _40118_ (.LO(trace_data[35]));
 sky130_fd_sc_hd__conb_1 _40119_ (.LO(trace_valid));
 sky130_fd_sc_hd__conb_1 _40120_ (.LO(_00313_));
 sky130_fd_sc_hd__buf_2 _40121_ (.A(mem_la_wdata[0]),
    .X(pcpi_rs2[0]));
 sky130_fd_sc_hd__buf_2 _40122_ (.A(mem_la_wdata[1]),
    .X(pcpi_rs2[1]));
 sky130_fd_sc_hd__buf_2 _40123_ (.A(mem_la_wdata[2]),
    .X(pcpi_rs2[2]));
 sky130_fd_sc_hd__buf_2 _40124_ (.A(mem_la_wdata[3]),
    .X(pcpi_rs2[3]));
 sky130_fd_sc_hd__buf_2 _40125_ (.A(mem_la_wdata[4]),
    .X(pcpi_rs2[4]));
 sky130_fd_sc_hd__buf_2 _40126_ (.A(mem_la_wdata[5]),
    .X(pcpi_rs2[5]));
 sky130_fd_sc_hd__buf_2 _40127_ (.A(mem_la_wdata[6]),
    .X(pcpi_rs2[6]));
 sky130_fd_sc_hd__buf_2 _40128_ (.A(mem_la_wdata[7]),
    .X(pcpi_rs2[7]));
 sky130_fd_sc_hd__mux2_1 _40129_ (.A0(decoder_trigger),
    .A1(_02410_),
    .S(_00309_),
    .X(_20586_));
 sky130_fd_sc_hd__mux2_1 _40130_ (.A0(\reg_out[2] ),
    .A1(\reg_next_pc[2] ),
    .S(_02183_),
    .X(_02184_));
 sky130_fd_sc_hd__mux2_1 _40131_ (.A0(_02184_),
    .A1(pcpi_rs1[2]),
    .S(_00301_),
    .X(mem_la_addr[2]));
 sky130_fd_sc_hd__mux2_1 _40132_ (.A0(\reg_out[3] ),
    .A1(\reg_next_pc[3] ),
    .S(_02183_),
    .X(_02185_));
 sky130_fd_sc_hd__mux2_1 _40133_ (.A0(_02185_),
    .A1(pcpi_rs1[3]),
    .S(_00301_),
    .X(mem_la_addr[3]));
 sky130_fd_sc_hd__mux2_1 _40134_ (.A0(\reg_out[4] ),
    .A1(\reg_next_pc[4] ),
    .S(_02183_),
    .X(_02186_));
 sky130_fd_sc_hd__mux2_1 _40135_ (.A0(_02186_),
    .A1(pcpi_rs1[4]),
    .S(_00301_),
    .X(mem_la_addr[4]));
 sky130_fd_sc_hd__mux2_1 _40136_ (.A0(\reg_out[5] ),
    .A1(\reg_next_pc[5] ),
    .S(_02183_),
    .X(_02187_));
 sky130_fd_sc_hd__mux2_1 _40137_ (.A0(_02187_),
    .A1(pcpi_rs1[5]),
    .S(_00301_),
    .X(mem_la_addr[5]));
 sky130_fd_sc_hd__mux2_1 _40138_ (.A0(\reg_out[6] ),
    .A1(\reg_next_pc[6] ),
    .S(_02183_),
    .X(_02188_));
 sky130_fd_sc_hd__mux2_1 _40139_ (.A0(_02188_),
    .A1(pcpi_rs1[6]),
    .S(_00301_),
    .X(mem_la_addr[6]));
 sky130_fd_sc_hd__mux2_1 _40140_ (.A0(\reg_out[7] ),
    .A1(\reg_next_pc[7] ),
    .S(_02183_),
    .X(_02189_));
 sky130_fd_sc_hd__mux2_1 _40141_ (.A0(_02189_),
    .A1(pcpi_rs1[7]),
    .S(_00301_),
    .X(mem_la_addr[7]));
 sky130_fd_sc_hd__mux2_1 _40142_ (.A0(\reg_out[8] ),
    .A1(\reg_next_pc[8] ),
    .S(_02183_),
    .X(_02190_));
 sky130_fd_sc_hd__mux2_1 _40143_ (.A0(_02190_),
    .A1(pcpi_rs1[8]),
    .S(_00301_),
    .X(mem_la_addr[8]));
 sky130_fd_sc_hd__mux2_1 _40144_ (.A0(\reg_out[9] ),
    .A1(\reg_next_pc[9] ),
    .S(_02183_),
    .X(_02191_));
 sky130_fd_sc_hd__mux2_1 _40145_ (.A0(_02191_),
    .A1(pcpi_rs1[9]),
    .S(_00301_),
    .X(mem_la_addr[9]));
 sky130_fd_sc_hd__mux2_1 _40146_ (.A0(\reg_out[10] ),
    .A1(\reg_next_pc[10] ),
    .S(_02183_),
    .X(_02192_));
 sky130_fd_sc_hd__mux2_1 _40147_ (.A0(_02192_),
    .A1(pcpi_rs1[10]),
    .S(_00301_),
    .X(mem_la_addr[10]));
 sky130_fd_sc_hd__mux2_1 _40148_ (.A0(\reg_out[11] ),
    .A1(\reg_next_pc[11] ),
    .S(_02183_),
    .X(_02193_));
 sky130_fd_sc_hd__mux2_1 _40149_ (.A0(_02193_),
    .A1(pcpi_rs1[11]),
    .S(_00301_),
    .X(mem_la_addr[11]));
 sky130_fd_sc_hd__mux2_1 _40150_ (.A0(\reg_out[12] ),
    .A1(\reg_next_pc[12] ),
    .S(_02183_),
    .X(_02194_));
 sky130_fd_sc_hd__mux2_1 _40151_ (.A0(_02194_),
    .A1(pcpi_rs1[12]),
    .S(_00301_),
    .X(mem_la_addr[12]));
 sky130_fd_sc_hd__mux2_1 _40152_ (.A0(\reg_out[13] ),
    .A1(\reg_next_pc[13] ),
    .S(_02183_),
    .X(_02195_));
 sky130_fd_sc_hd__mux2_1 _40153_ (.A0(_02195_),
    .A1(pcpi_rs1[13]),
    .S(_00301_),
    .X(mem_la_addr[13]));
 sky130_fd_sc_hd__mux2_1 _40154_ (.A0(\reg_out[14] ),
    .A1(\reg_next_pc[14] ),
    .S(_02183_),
    .X(_02196_));
 sky130_fd_sc_hd__mux2_1 _40155_ (.A0(_02196_),
    .A1(pcpi_rs1[14]),
    .S(_00301_),
    .X(mem_la_addr[14]));
 sky130_fd_sc_hd__mux2_1 _40156_ (.A0(\reg_out[15] ),
    .A1(\reg_next_pc[15] ),
    .S(_02183_),
    .X(_02197_));
 sky130_fd_sc_hd__mux2_1 _40157_ (.A0(_02197_),
    .A1(pcpi_rs1[15]),
    .S(_00301_),
    .X(mem_la_addr[15]));
 sky130_fd_sc_hd__mux2_1 _40158_ (.A0(\reg_out[16] ),
    .A1(\reg_next_pc[16] ),
    .S(_02183_),
    .X(_02198_));
 sky130_fd_sc_hd__mux2_1 _40159_ (.A0(_02198_),
    .A1(pcpi_rs1[16]),
    .S(_00301_),
    .X(mem_la_addr[16]));
 sky130_fd_sc_hd__mux2_1 _40160_ (.A0(\reg_out[17] ),
    .A1(\reg_next_pc[17] ),
    .S(_02183_),
    .X(_02199_));
 sky130_fd_sc_hd__mux2_1 _40161_ (.A0(_02199_),
    .A1(pcpi_rs1[17]),
    .S(_00301_),
    .X(mem_la_addr[17]));
 sky130_fd_sc_hd__mux2_1 _40162_ (.A0(\reg_out[18] ),
    .A1(\reg_next_pc[18] ),
    .S(_02183_),
    .X(_02200_));
 sky130_fd_sc_hd__mux2_1 _40163_ (.A0(_02200_),
    .A1(pcpi_rs1[18]),
    .S(_00301_),
    .X(mem_la_addr[18]));
 sky130_fd_sc_hd__mux2_1 _40164_ (.A0(\reg_out[19] ),
    .A1(\reg_next_pc[19] ),
    .S(_02183_),
    .X(_02201_));
 sky130_fd_sc_hd__mux2_1 _40165_ (.A0(_02201_),
    .A1(pcpi_rs1[19]),
    .S(_00301_),
    .X(mem_la_addr[19]));
 sky130_fd_sc_hd__mux2_1 _40166_ (.A0(\reg_out[20] ),
    .A1(\reg_next_pc[20] ),
    .S(_02183_),
    .X(_02202_));
 sky130_fd_sc_hd__mux2_1 _40167_ (.A0(_02202_),
    .A1(pcpi_rs1[20]),
    .S(_00301_),
    .X(mem_la_addr[20]));
 sky130_fd_sc_hd__mux2_1 _40168_ (.A0(\reg_out[21] ),
    .A1(\reg_next_pc[21] ),
    .S(_02183_),
    .X(_02203_));
 sky130_fd_sc_hd__mux2_1 _40169_ (.A0(_02203_),
    .A1(pcpi_rs1[21]),
    .S(_00301_),
    .X(mem_la_addr[21]));
 sky130_fd_sc_hd__mux2_1 _40170_ (.A0(\reg_out[22] ),
    .A1(\reg_next_pc[22] ),
    .S(_02183_),
    .X(_02204_));
 sky130_fd_sc_hd__mux2_1 _40171_ (.A0(_02204_),
    .A1(pcpi_rs1[22]),
    .S(_00301_),
    .X(mem_la_addr[22]));
 sky130_fd_sc_hd__mux2_1 _40172_ (.A0(\reg_out[23] ),
    .A1(\reg_next_pc[23] ),
    .S(_02183_),
    .X(_02205_));
 sky130_fd_sc_hd__mux2_1 _40173_ (.A0(_02205_),
    .A1(pcpi_rs1[23]),
    .S(_00301_),
    .X(mem_la_addr[23]));
 sky130_fd_sc_hd__mux2_1 _40174_ (.A0(\reg_out[24] ),
    .A1(\reg_next_pc[24] ),
    .S(_02183_),
    .X(_02206_));
 sky130_fd_sc_hd__mux2_1 _40175_ (.A0(_02206_),
    .A1(pcpi_rs1[24]),
    .S(_00301_),
    .X(mem_la_addr[24]));
 sky130_fd_sc_hd__mux2_1 _40176_ (.A0(\reg_out[25] ),
    .A1(\reg_next_pc[25] ),
    .S(_02183_),
    .X(_02207_));
 sky130_fd_sc_hd__mux2_1 _40177_ (.A0(_02207_),
    .A1(pcpi_rs1[25]),
    .S(_00301_),
    .X(mem_la_addr[25]));
 sky130_fd_sc_hd__mux2_1 _40178_ (.A0(\reg_out[26] ),
    .A1(\reg_next_pc[26] ),
    .S(_02183_),
    .X(_02208_));
 sky130_fd_sc_hd__mux2_1 _40179_ (.A0(_02208_),
    .A1(pcpi_rs1[26]),
    .S(_00301_),
    .X(mem_la_addr[26]));
 sky130_fd_sc_hd__mux2_1 _40180_ (.A0(\reg_out[27] ),
    .A1(\reg_next_pc[27] ),
    .S(_02183_),
    .X(_02209_));
 sky130_fd_sc_hd__mux2_1 _40181_ (.A0(_02209_),
    .A1(pcpi_rs1[27]),
    .S(_00301_),
    .X(mem_la_addr[27]));
 sky130_fd_sc_hd__mux2_1 _40182_ (.A0(\reg_out[28] ),
    .A1(\reg_next_pc[28] ),
    .S(_02183_),
    .X(_02210_));
 sky130_fd_sc_hd__mux2_1 _40183_ (.A0(_02210_),
    .A1(pcpi_rs1[28]),
    .S(_00301_),
    .X(mem_la_addr[28]));
 sky130_fd_sc_hd__mux2_1 _40184_ (.A0(\reg_out[29] ),
    .A1(\reg_next_pc[29] ),
    .S(_02183_),
    .X(_02211_));
 sky130_fd_sc_hd__mux2_1 _40185_ (.A0(_02211_),
    .A1(pcpi_rs1[29]),
    .S(_00301_),
    .X(mem_la_addr[29]));
 sky130_fd_sc_hd__mux2_1 _40186_ (.A0(\reg_out[30] ),
    .A1(\reg_next_pc[30] ),
    .S(_02183_),
    .X(_02212_));
 sky130_fd_sc_hd__mux2_1 _40187_ (.A0(_02212_),
    .A1(pcpi_rs1[30]),
    .S(_00301_),
    .X(mem_la_addr[30]));
 sky130_fd_sc_hd__mux2_1 _40188_ (.A0(\reg_out[31] ),
    .A1(\reg_next_pc[31] ),
    .S(_02183_),
    .X(_02213_));
 sky130_fd_sc_hd__mux2_1 _40189_ (.A0(_02213_),
    .A1(pcpi_rs1[31]),
    .S(_00301_),
    .X(mem_la_addr[31]));
 sky130_fd_sc_hd__mux2_1 _40190_ (.A0(_02167_),
    .A1(pcpi_rs2[8]),
    .S(_01683_),
    .X(mem_la_wdata[8]));
 sky130_fd_sc_hd__mux2_1 _40191_ (.A0(_02168_),
    .A1(pcpi_rs2[9]),
    .S(_01683_),
    .X(mem_la_wdata[9]));
 sky130_fd_sc_hd__mux2_1 _40192_ (.A0(_02169_),
    .A1(pcpi_rs2[10]),
    .S(_01683_),
    .X(mem_la_wdata[10]));
 sky130_fd_sc_hd__mux2_1 _40193_ (.A0(_02170_),
    .A1(pcpi_rs2[11]),
    .S(_01683_),
    .X(mem_la_wdata[11]));
 sky130_fd_sc_hd__mux2_1 _40194_ (.A0(_02171_),
    .A1(pcpi_rs2[12]),
    .S(_01683_),
    .X(mem_la_wdata[12]));
 sky130_fd_sc_hd__mux2_1 _40195_ (.A0(_02172_),
    .A1(pcpi_rs2[13]),
    .S(_01683_),
    .X(mem_la_wdata[13]));
 sky130_fd_sc_hd__mux2_1 _40196_ (.A0(_02173_),
    .A1(pcpi_rs2[14]),
    .S(_01683_),
    .X(mem_la_wdata[14]));
 sky130_fd_sc_hd__mux2_1 _40197_ (.A0(_02174_),
    .A1(pcpi_rs2[15]),
    .S(_01683_),
    .X(mem_la_wdata[15]));
 sky130_fd_sc_hd__mux2_1 _40198_ (.A0(_02175_),
    .A1(pcpi_rs2[16]),
    .S(_01683_),
    .X(mem_la_wdata[16]));
 sky130_fd_sc_hd__mux2_1 _40199_ (.A0(_02176_),
    .A1(pcpi_rs2[17]),
    .S(_01683_),
    .X(mem_la_wdata[17]));
 sky130_fd_sc_hd__mux2_1 _40200_ (.A0(_02177_),
    .A1(pcpi_rs2[18]),
    .S(_01683_),
    .X(mem_la_wdata[18]));
 sky130_fd_sc_hd__mux2_1 _40201_ (.A0(_02178_),
    .A1(pcpi_rs2[19]),
    .S(_01683_),
    .X(mem_la_wdata[19]));
 sky130_fd_sc_hd__mux2_1 _40202_ (.A0(_02179_),
    .A1(pcpi_rs2[20]),
    .S(_01683_),
    .X(mem_la_wdata[20]));
 sky130_fd_sc_hd__mux2_1 _40203_ (.A0(_02180_),
    .A1(pcpi_rs2[21]),
    .S(_01683_),
    .X(mem_la_wdata[21]));
 sky130_fd_sc_hd__mux2_1 _40204_ (.A0(_02181_),
    .A1(pcpi_rs2[22]),
    .S(_01683_),
    .X(mem_la_wdata[22]));
 sky130_fd_sc_hd__mux2_1 _40205_ (.A0(_02182_),
    .A1(pcpi_rs2[23]),
    .S(_01683_),
    .X(mem_la_wdata[23]));
 sky130_fd_sc_hd__mux2_1 _40206_ (.A0(_02167_),
    .A1(pcpi_rs2[24]),
    .S(_01683_),
    .X(mem_la_wdata[24]));
 sky130_fd_sc_hd__mux2_1 _40207_ (.A0(_02168_),
    .A1(pcpi_rs2[25]),
    .S(_01683_),
    .X(mem_la_wdata[25]));
 sky130_fd_sc_hd__mux2_1 _40208_ (.A0(_02169_),
    .A1(pcpi_rs2[26]),
    .S(_01683_),
    .X(mem_la_wdata[26]));
 sky130_fd_sc_hd__mux2_1 _40209_ (.A0(_02170_),
    .A1(pcpi_rs2[27]),
    .S(_01683_),
    .X(mem_la_wdata[27]));
 sky130_fd_sc_hd__mux2_1 _40210_ (.A0(_02171_),
    .A1(pcpi_rs2[28]),
    .S(_01683_),
    .X(mem_la_wdata[28]));
 sky130_fd_sc_hd__mux2_1 _40211_ (.A0(_02172_),
    .A1(pcpi_rs2[29]),
    .S(_01683_),
    .X(mem_la_wdata[29]));
 sky130_fd_sc_hd__mux2_1 _40212_ (.A0(_02173_),
    .A1(pcpi_rs2[30]),
    .S(_01683_),
    .X(mem_la_wdata[30]));
 sky130_fd_sc_hd__mux2_1 _40213_ (.A0(_02174_),
    .A1(pcpi_rs2[31]),
    .S(_01683_),
    .X(mem_la_wdata[31]));
 sky130_fd_sc_hd__mux2_1 _40214_ (.A0(\mem_rdata_q[7] ),
    .A1(mem_rdata[7]),
    .S(mem_xfer),
    .X(\mem_rdata_latched[7] ));
 sky130_fd_sc_hd__mux2_1 _40215_ (.A0(\mem_rdata_q[8] ),
    .A1(mem_rdata[8]),
    .S(mem_xfer),
    .X(\mem_rdata_latched[8] ));
 sky130_fd_sc_hd__mux2_1 _40216_ (.A0(\mem_rdata_q[9] ),
    .A1(mem_rdata[9]),
    .S(mem_xfer),
    .X(\mem_rdata_latched[9] ));
 sky130_fd_sc_hd__mux2_1 _40217_ (.A0(\mem_rdata_q[10] ),
    .A1(mem_rdata[10]),
    .S(mem_xfer),
    .X(\mem_rdata_latched[10] ));
 sky130_fd_sc_hd__mux2_1 _40218_ (.A0(\mem_rdata_q[11] ),
    .A1(mem_rdata[11]),
    .S(mem_xfer),
    .X(\mem_rdata_latched[11] ));
 sky130_fd_sc_hd__mux2_1 _40219_ (.A0(\mem_rdata_q[12] ),
    .A1(mem_rdata[12]),
    .S(mem_xfer),
    .X(\mem_rdata_latched[12] ));
 sky130_fd_sc_hd__mux2_1 _40220_ (.A0(\mem_rdata_q[13] ),
    .A1(mem_rdata[13]),
    .S(mem_xfer),
    .X(\mem_rdata_latched[13] ));
 sky130_fd_sc_hd__mux2_1 _40221_ (.A0(\mem_rdata_q[14] ),
    .A1(mem_rdata[14]),
    .S(mem_xfer),
    .X(\mem_rdata_latched[14] ));
 sky130_fd_sc_hd__mux2_1 _40222_ (.A0(\mem_rdata_q[15] ),
    .A1(mem_rdata[15]),
    .S(mem_xfer),
    .X(\mem_rdata_latched[15] ));
 sky130_fd_sc_hd__mux2_1 _40223_ (.A0(\mem_rdata_q[16] ),
    .A1(mem_rdata[16]),
    .S(mem_xfer),
    .X(\mem_rdata_latched[16] ));
 sky130_fd_sc_hd__mux2_1 _40224_ (.A0(\mem_rdata_q[17] ),
    .A1(mem_rdata[17]),
    .S(mem_xfer),
    .X(\mem_rdata_latched[17] ));
 sky130_fd_sc_hd__mux2_1 _40225_ (.A0(\mem_rdata_q[18] ),
    .A1(mem_rdata[18]),
    .S(mem_xfer),
    .X(\mem_rdata_latched[18] ));
 sky130_fd_sc_hd__mux2_1 _40226_ (.A0(\mem_rdata_q[19] ),
    .A1(mem_rdata[19]),
    .S(mem_xfer),
    .X(\mem_rdata_latched[19] ));
 sky130_fd_sc_hd__mux2_1 _40227_ (.A0(\mem_rdata_q[20] ),
    .A1(mem_rdata[20]),
    .S(mem_xfer),
    .X(\mem_rdata_latched[20] ));
 sky130_fd_sc_hd__mux2_1 _40228_ (.A0(\mem_rdata_q[21] ),
    .A1(mem_rdata[21]),
    .S(mem_xfer),
    .X(\mem_rdata_latched[21] ));
 sky130_fd_sc_hd__mux2_1 _40229_ (.A0(\mem_rdata_q[22] ),
    .A1(mem_rdata[22]),
    .S(mem_xfer),
    .X(\mem_rdata_latched[22] ));
 sky130_fd_sc_hd__mux2_1 _40230_ (.A0(\mem_rdata_q[23] ),
    .A1(mem_rdata[23]),
    .S(mem_xfer),
    .X(\mem_rdata_latched[23] ));
 sky130_fd_sc_hd__mux2_1 _40231_ (.A0(\mem_rdata_q[24] ),
    .A1(mem_rdata[24]),
    .S(mem_xfer),
    .X(\mem_rdata_latched[24] ));
 sky130_fd_sc_hd__mux2_1 _40232_ (.A0(\mem_rdata_q[25] ),
    .A1(mem_rdata[25]),
    .S(mem_xfer),
    .X(\mem_rdata_latched[25] ));
 sky130_fd_sc_hd__mux2_1 _40233_ (.A0(\mem_rdata_q[26] ),
    .A1(mem_rdata[26]),
    .S(mem_xfer),
    .X(\mem_rdata_latched[26] ));
 sky130_fd_sc_hd__mux2_1 _40234_ (.A0(\mem_rdata_q[27] ),
    .A1(mem_rdata[27]),
    .S(mem_xfer),
    .X(\mem_rdata_latched[27] ));
 sky130_fd_sc_hd__mux2_1 _40235_ (.A0(\mem_rdata_q[28] ),
    .A1(mem_rdata[28]),
    .S(mem_xfer),
    .X(\mem_rdata_latched[28] ));
 sky130_fd_sc_hd__mux2_1 _40236_ (.A0(\mem_rdata_q[29] ),
    .A1(mem_rdata[29]),
    .S(mem_xfer),
    .X(\mem_rdata_latched[29] ));
 sky130_fd_sc_hd__mux2_1 _40237_ (.A0(\mem_rdata_q[30] ),
    .A1(mem_rdata[30]),
    .S(mem_xfer),
    .X(\mem_rdata_latched[30] ));
 sky130_fd_sc_hd__mux2_1 _40238_ (.A0(\mem_rdata_q[31] ),
    .A1(mem_rdata[31]),
    .S(mem_xfer),
    .X(\mem_rdata_latched[31] ));
 sky130_fd_sc_hd__mux2_1 _40239_ (.A0(_02134_),
    .A1(\alu_add_sub[0] ),
    .S(_02133_),
    .X(\alu_out[0] ));
 sky130_fd_sc_hd__mux2_1 _40240_ (.A0(_02135_),
    .A1(\alu_add_sub[1] ),
    .S(_02133_),
    .X(\alu_out[1] ));
 sky130_fd_sc_hd__mux2_1 _40241_ (.A0(_02136_),
    .A1(\alu_add_sub[2] ),
    .S(_02133_),
    .X(\alu_out[2] ));
 sky130_fd_sc_hd__mux2_1 _40242_ (.A0(_02137_),
    .A1(\alu_add_sub[3] ),
    .S(_02133_),
    .X(\alu_out[3] ));
 sky130_fd_sc_hd__mux2_1 _40243_ (.A0(_02138_),
    .A1(\alu_add_sub[4] ),
    .S(_02133_),
    .X(\alu_out[4] ));
 sky130_fd_sc_hd__mux2_1 _40244_ (.A0(_02139_),
    .A1(\alu_add_sub[5] ),
    .S(_02133_),
    .X(\alu_out[5] ));
 sky130_fd_sc_hd__mux2_1 _40245_ (.A0(_02140_),
    .A1(\alu_add_sub[6] ),
    .S(_02133_),
    .X(\alu_out[6] ));
 sky130_fd_sc_hd__mux2_1 _40246_ (.A0(_02141_),
    .A1(\alu_add_sub[7] ),
    .S(_02133_),
    .X(\alu_out[7] ));
 sky130_fd_sc_hd__mux2_1 _40247_ (.A0(_02142_),
    .A1(\alu_add_sub[8] ),
    .S(_02133_),
    .X(\alu_out[8] ));
 sky130_fd_sc_hd__mux2_1 _40248_ (.A0(_02143_),
    .A1(\alu_add_sub[9] ),
    .S(_02133_),
    .X(\alu_out[9] ));
 sky130_fd_sc_hd__mux2_1 _40249_ (.A0(_02144_),
    .A1(\alu_add_sub[10] ),
    .S(_02133_),
    .X(\alu_out[10] ));
 sky130_fd_sc_hd__mux2_1 _40250_ (.A0(_02145_),
    .A1(\alu_add_sub[11] ),
    .S(_02133_),
    .X(\alu_out[11] ));
 sky130_fd_sc_hd__mux2_1 _40251_ (.A0(_02146_),
    .A1(\alu_add_sub[12] ),
    .S(_02133_),
    .X(\alu_out[12] ));
 sky130_fd_sc_hd__mux2_1 _40252_ (.A0(_02147_),
    .A1(\alu_add_sub[13] ),
    .S(_02133_),
    .X(\alu_out[13] ));
 sky130_fd_sc_hd__mux2_1 _40253_ (.A0(_02148_),
    .A1(\alu_add_sub[14] ),
    .S(_02133_),
    .X(\alu_out[14] ));
 sky130_fd_sc_hd__mux2_1 _40254_ (.A0(_02149_),
    .A1(\alu_add_sub[15] ),
    .S(_02133_),
    .X(\alu_out[15] ));
 sky130_fd_sc_hd__mux2_1 _40255_ (.A0(_02150_),
    .A1(\alu_add_sub[16] ),
    .S(_02133_),
    .X(\alu_out[16] ));
 sky130_fd_sc_hd__mux2_1 _40256_ (.A0(_02151_),
    .A1(\alu_add_sub[17] ),
    .S(_02133_),
    .X(\alu_out[17] ));
 sky130_fd_sc_hd__mux2_1 _40257_ (.A0(_02152_),
    .A1(\alu_add_sub[18] ),
    .S(_02133_),
    .X(\alu_out[18] ));
 sky130_fd_sc_hd__mux2_1 _40258_ (.A0(_02153_),
    .A1(\alu_add_sub[19] ),
    .S(_02133_),
    .X(\alu_out[19] ));
 sky130_fd_sc_hd__mux2_1 _40259_ (.A0(_02154_),
    .A1(\alu_add_sub[20] ),
    .S(_02133_),
    .X(\alu_out[20] ));
 sky130_fd_sc_hd__mux2_1 _40260_ (.A0(_02155_),
    .A1(\alu_add_sub[21] ),
    .S(_02133_),
    .X(\alu_out[21] ));
 sky130_fd_sc_hd__mux2_1 _40261_ (.A0(_02156_),
    .A1(\alu_add_sub[22] ),
    .S(_02133_),
    .X(\alu_out[22] ));
 sky130_fd_sc_hd__mux2_1 _40262_ (.A0(_02157_),
    .A1(\alu_add_sub[23] ),
    .S(_02133_),
    .X(\alu_out[23] ));
 sky130_fd_sc_hd__mux2_1 _40263_ (.A0(_02158_),
    .A1(\alu_add_sub[24] ),
    .S(_02133_),
    .X(\alu_out[24] ));
 sky130_fd_sc_hd__mux2_1 _40264_ (.A0(_02159_),
    .A1(\alu_add_sub[25] ),
    .S(_02133_),
    .X(\alu_out[25] ));
 sky130_fd_sc_hd__mux2_1 _40265_ (.A0(_02160_),
    .A1(\alu_add_sub[26] ),
    .S(_02133_),
    .X(\alu_out[26] ));
 sky130_fd_sc_hd__mux2_1 _40266_ (.A0(_02161_),
    .A1(\alu_add_sub[27] ),
    .S(_02133_),
    .X(\alu_out[27] ));
 sky130_fd_sc_hd__mux2_1 _40267_ (.A0(_02162_),
    .A1(\alu_add_sub[28] ),
    .S(_02133_),
    .X(\alu_out[28] ));
 sky130_fd_sc_hd__mux2_1 _40268_ (.A0(_02163_),
    .A1(\alu_add_sub[29] ),
    .S(_02133_),
    .X(\alu_out[29] ));
 sky130_fd_sc_hd__mux2_1 _40269_ (.A0(_02164_),
    .A1(\alu_add_sub[30] ),
    .S(_02133_),
    .X(\alu_out[30] ));
 sky130_fd_sc_hd__mux2_1 _40270_ (.A0(_02165_),
    .A1(\alu_add_sub[31] ),
    .S(_02133_),
    .X(\alu_out[31] ));
 sky130_fd_sc_hd__mux2_1 _40271_ (.A0(_02071_),
    .A1(\reg_next_pc[0] ),
    .S(_02069_),
    .X(\cpuregs_wrdata[0] ));
 sky130_fd_sc_hd__mux2_1 _40272_ (.A0(_02072_),
    .A1(\reg_pc[1] ),
    .S(_02069_),
    .X(\cpuregs_wrdata[1] ));
 sky130_fd_sc_hd__mux2_1 _40273_ (.A0(_02074_),
    .A1(_02073_),
    .S(_02069_),
    .X(\cpuregs_wrdata[2] ));
 sky130_fd_sc_hd__mux2_1 _40274_ (.A0(_02076_),
    .A1(_02075_),
    .S(_02069_),
    .X(\cpuregs_wrdata[3] ));
 sky130_fd_sc_hd__mux2_1 _40275_ (.A0(_02078_),
    .A1(_02077_),
    .S(_02069_),
    .X(\cpuregs_wrdata[4] ));
 sky130_fd_sc_hd__mux2_1 _40276_ (.A0(_02080_),
    .A1(_02079_),
    .S(_02069_),
    .X(\cpuregs_wrdata[5] ));
 sky130_fd_sc_hd__mux2_1 _40277_ (.A0(_02082_),
    .A1(_02081_),
    .S(_02069_),
    .X(\cpuregs_wrdata[6] ));
 sky130_fd_sc_hd__mux2_1 _40278_ (.A0(_02084_),
    .A1(_02083_),
    .S(_02069_),
    .X(\cpuregs_wrdata[7] ));
 sky130_fd_sc_hd__mux2_1 _40279_ (.A0(_02086_),
    .A1(_02085_),
    .S(_02069_),
    .X(\cpuregs_wrdata[8] ));
 sky130_fd_sc_hd__mux2_1 _40280_ (.A0(_02088_),
    .A1(_02087_),
    .S(_02069_),
    .X(\cpuregs_wrdata[9] ));
 sky130_fd_sc_hd__mux2_1 _40281_ (.A0(_02090_),
    .A1(_02089_),
    .S(_02069_),
    .X(\cpuregs_wrdata[10] ));
 sky130_fd_sc_hd__mux2_1 _40282_ (.A0(_02092_),
    .A1(_02091_),
    .S(_02069_),
    .X(\cpuregs_wrdata[11] ));
 sky130_fd_sc_hd__mux2_1 _40283_ (.A0(_02094_),
    .A1(_02093_),
    .S(_02069_),
    .X(\cpuregs_wrdata[12] ));
 sky130_fd_sc_hd__mux2_1 _40284_ (.A0(_02096_),
    .A1(_02095_),
    .S(_02069_),
    .X(\cpuregs_wrdata[13] ));
 sky130_fd_sc_hd__mux2_1 _40285_ (.A0(_02098_),
    .A1(_02097_),
    .S(_02069_),
    .X(\cpuregs_wrdata[14] ));
 sky130_fd_sc_hd__mux2_1 _40286_ (.A0(_02100_),
    .A1(_02099_),
    .S(_02069_),
    .X(\cpuregs_wrdata[15] ));
 sky130_fd_sc_hd__mux2_1 _40287_ (.A0(_02102_),
    .A1(_02101_),
    .S(_02069_),
    .X(\cpuregs_wrdata[16] ));
 sky130_fd_sc_hd__mux2_1 _40288_ (.A0(_02104_),
    .A1(_02103_),
    .S(_02069_),
    .X(\cpuregs_wrdata[17] ));
 sky130_fd_sc_hd__mux2_1 _40289_ (.A0(_02106_),
    .A1(_02105_),
    .S(_02069_),
    .X(\cpuregs_wrdata[18] ));
 sky130_fd_sc_hd__mux2_1 _40290_ (.A0(_02108_),
    .A1(_02107_),
    .S(_02069_),
    .X(\cpuregs_wrdata[19] ));
 sky130_fd_sc_hd__mux2_1 _40291_ (.A0(_02110_),
    .A1(_02109_),
    .S(_02069_),
    .X(\cpuregs_wrdata[20] ));
 sky130_fd_sc_hd__mux2_1 _40292_ (.A0(_02112_),
    .A1(_02111_),
    .S(_02069_),
    .X(\cpuregs_wrdata[21] ));
 sky130_fd_sc_hd__mux2_1 _40293_ (.A0(_02114_),
    .A1(_02113_),
    .S(_02069_),
    .X(\cpuregs_wrdata[22] ));
 sky130_fd_sc_hd__mux2_1 _40294_ (.A0(_02116_),
    .A1(_02115_),
    .S(_02069_),
    .X(\cpuregs_wrdata[23] ));
 sky130_fd_sc_hd__mux2_1 _40295_ (.A0(_02118_),
    .A1(_02117_),
    .S(_02069_),
    .X(\cpuregs_wrdata[24] ));
 sky130_fd_sc_hd__mux2_1 _40296_ (.A0(_02120_),
    .A1(_02119_),
    .S(_02069_),
    .X(\cpuregs_wrdata[25] ));
 sky130_fd_sc_hd__mux2_1 _40297_ (.A0(_02122_),
    .A1(_02121_),
    .S(_02069_),
    .X(\cpuregs_wrdata[26] ));
 sky130_fd_sc_hd__mux2_1 _40298_ (.A0(_02124_),
    .A1(_02123_),
    .S(_02069_),
    .X(\cpuregs_wrdata[27] ));
 sky130_fd_sc_hd__mux2_1 _40299_ (.A0(_02126_),
    .A1(_02125_),
    .S(_02069_),
    .X(\cpuregs_wrdata[28] ));
 sky130_fd_sc_hd__mux2_1 _40300_ (.A0(_02128_),
    .A1(_02127_),
    .S(_02069_),
    .X(\cpuregs_wrdata[29] ));
 sky130_fd_sc_hd__mux2_1 _40301_ (.A0(_02130_),
    .A1(_02129_),
    .S(_02069_),
    .X(\cpuregs_wrdata[30] ));
 sky130_fd_sc_hd__mux2_1 _40302_ (.A0(_02132_),
    .A1(_02131_),
    .S(_02069_),
    .X(\cpuregs_wrdata[31] ));
 sky130_fd_sc_hd__mux2_1 _40303_ (.A0(_02316_),
    .A1(_02317_),
    .S(_00307_),
    .X(_00004_));
 sky130_fd_sc_hd__mux2_1 _40304_ (.A0(_00347_),
    .A1(_20587_),
    .S(_00336_),
    .X(_00348_));
 sky130_fd_sc_hd__mux2_1 _40305_ (.A0(_20587_),
    .A1(_00348_),
    .S(resetn),
    .X(_00003_));
 sky130_fd_sc_hd__mux2_1 _40306_ (.A0(_02304_),
    .A1(_02305_),
    .S(\irq_state[1] ),
    .X(_02306_));
 sky130_fd_sc_hd__mux2_1 _40307_ (.A0(_02306_),
    .A1(_02304_),
    .S(_02217_),
    .X(_00008_));
 sky130_fd_sc_hd__mux2_1 _40308_ (.A0(_02214_),
    .A1(_02215_),
    .S(\irq_state[1] ),
    .X(_02216_));
 sky130_fd_sc_hd__mux2_1 _40309_ (.A0(_02216_),
    .A1(_02214_),
    .S(_02217_),
    .X(_00031_));
 sky130_fd_sc_hd__mux2_1 _40310_ (.A0(_02218_),
    .A1(_02219_),
    .S(\irq_state[1] ),
    .X(_02220_));
 sky130_fd_sc_hd__mux2_1 _40311_ (.A0(_02220_),
    .A1(_02218_),
    .S(_02217_),
    .X(_00032_));
 sky130_fd_sc_hd__mux2_1 _40312_ (.A0(_02221_),
    .A1(_02222_),
    .S(\irq_state[1] ),
    .X(_02223_));
 sky130_fd_sc_hd__mux2_1 _40313_ (.A0(_02223_),
    .A1(_02221_),
    .S(_02217_),
    .X(_00033_));
 sky130_fd_sc_hd__mux2_1 _40314_ (.A0(_02224_),
    .A1(_02225_),
    .S(\irq_state[1] ),
    .X(_02226_));
 sky130_fd_sc_hd__mux2_1 _40315_ (.A0(_02226_),
    .A1(_02224_),
    .S(_02217_),
    .X(_00034_));
 sky130_fd_sc_hd__mux2_1 _40316_ (.A0(_02227_),
    .A1(_02228_),
    .S(\irq_state[1] ),
    .X(_02229_));
 sky130_fd_sc_hd__mux2_1 _40317_ (.A0(_02229_),
    .A1(_02227_),
    .S(_02217_),
    .X(_00035_));
 sky130_fd_sc_hd__mux2_1 _40318_ (.A0(_02230_),
    .A1(_02231_),
    .S(\irq_state[1] ),
    .X(_02232_));
 sky130_fd_sc_hd__mux2_1 _40319_ (.A0(_02232_),
    .A1(_02230_),
    .S(_02217_),
    .X(_00036_));
 sky130_fd_sc_hd__mux2_1 _40320_ (.A0(_02233_),
    .A1(_02234_),
    .S(\irq_state[1] ),
    .X(_02235_));
 sky130_fd_sc_hd__mux2_1 _40321_ (.A0(_02235_),
    .A1(_02233_),
    .S(_02217_),
    .X(_00037_));
 sky130_fd_sc_hd__mux2_1 _40322_ (.A0(_02236_),
    .A1(_02237_),
    .S(\irq_state[1] ),
    .X(_02238_));
 sky130_fd_sc_hd__mux2_1 _40323_ (.A0(_02238_),
    .A1(_02236_),
    .S(_02217_),
    .X(_00009_));
 sky130_fd_sc_hd__mux2_1 _40324_ (.A0(_02239_),
    .A1(_02240_),
    .S(\irq_state[1] ),
    .X(_02241_));
 sky130_fd_sc_hd__mux2_1 _40325_ (.A0(_02241_),
    .A1(_02239_),
    .S(_02217_),
    .X(_00010_));
 sky130_fd_sc_hd__mux2_1 _40326_ (.A0(_02242_),
    .A1(_02243_),
    .S(\irq_state[1] ),
    .X(_02244_));
 sky130_fd_sc_hd__mux2_1 _40327_ (.A0(_02244_),
    .A1(_02242_),
    .S(_02217_),
    .X(_00011_));
 sky130_fd_sc_hd__mux2_1 _40328_ (.A0(_02245_),
    .A1(_02246_),
    .S(\irq_state[1] ),
    .X(_02247_));
 sky130_fd_sc_hd__mux2_1 _40329_ (.A0(_02247_),
    .A1(_02245_),
    .S(_02217_),
    .X(_00012_));
 sky130_fd_sc_hd__mux2_1 _40330_ (.A0(_02248_),
    .A1(_02249_),
    .S(\irq_state[1] ),
    .X(_02250_));
 sky130_fd_sc_hd__mux2_1 _40331_ (.A0(_02250_),
    .A1(_02248_),
    .S(_02217_),
    .X(_00013_));
 sky130_fd_sc_hd__mux2_1 _40332_ (.A0(_02251_),
    .A1(_02252_),
    .S(\irq_state[1] ),
    .X(_02253_));
 sky130_fd_sc_hd__mux2_1 _40333_ (.A0(_02253_),
    .A1(_02251_),
    .S(_02217_),
    .X(_00014_));
 sky130_fd_sc_hd__mux2_1 _40334_ (.A0(_02254_),
    .A1(_02255_),
    .S(\irq_state[1] ),
    .X(_02256_));
 sky130_fd_sc_hd__mux2_1 _40335_ (.A0(_02256_),
    .A1(_02254_),
    .S(_02217_),
    .X(_00015_));
 sky130_fd_sc_hd__mux2_1 _40336_ (.A0(_02257_),
    .A1(_02258_),
    .S(\irq_state[1] ),
    .X(_02259_));
 sky130_fd_sc_hd__mux2_1 _40337_ (.A0(_02259_),
    .A1(_02257_),
    .S(_02217_),
    .X(_00016_));
 sky130_fd_sc_hd__mux2_1 _40338_ (.A0(_02260_),
    .A1(_02261_),
    .S(\irq_state[1] ),
    .X(_02262_));
 sky130_fd_sc_hd__mux2_1 _40339_ (.A0(_02262_),
    .A1(_02260_),
    .S(_02217_),
    .X(_00017_));
 sky130_fd_sc_hd__mux2_1 _40340_ (.A0(_02263_),
    .A1(_02264_),
    .S(\irq_state[1] ),
    .X(_02265_));
 sky130_fd_sc_hd__mux2_1 _40341_ (.A0(_02265_),
    .A1(_02263_),
    .S(_02217_),
    .X(_00018_));
 sky130_fd_sc_hd__mux2_1 _40342_ (.A0(_02266_),
    .A1(_02267_),
    .S(\irq_state[1] ),
    .X(_02268_));
 sky130_fd_sc_hd__mux2_1 _40343_ (.A0(_02268_),
    .A1(_02266_),
    .S(_02217_),
    .X(_00019_));
 sky130_fd_sc_hd__mux2_1 _40344_ (.A0(_02269_),
    .A1(_02270_),
    .S(\irq_state[1] ),
    .X(_02271_));
 sky130_fd_sc_hd__mux2_1 _40345_ (.A0(_02271_),
    .A1(_02269_),
    .S(_02217_),
    .X(_00020_));
 sky130_fd_sc_hd__mux2_1 _40346_ (.A0(_02272_),
    .A1(_02273_),
    .S(\irq_state[1] ),
    .X(_02274_));
 sky130_fd_sc_hd__mux2_1 _40347_ (.A0(_02274_),
    .A1(_02272_),
    .S(_02217_),
    .X(_00021_));
 sky130_fd_sc_hd__mux2_1 _40348_ (.A0(_02275_),
    .A1(_02276_),
    .S(\irq_state[1] ),
    .X(_02277_));
 sky130_fd_sc_hd__mux2_1 _40349_ (.A0(_02277_),
    .A1(_02275_),
    .S(_02217_),
    .X(_00022_));
 sky130_fd_sc_hd__mux2_1 _40350_ (.A0(_02278_),
    .A1(_02279_),
    .S(\irq_state[1] ),
    .X(_02280_));
 sky130_fd_sc_hd__mux2_1 _40351_ (.A0(_02280_),
    .A1(_02278_),
    .S(_02217_),
    .X(_00023_));
 sky130_fd_sc_hd__mux2_1 _40352_ (.A0(_02281_),
    .A1(_02282_),
    .S(\irq_state[1] ),
    .X(_02283_));
 sky130_fd_sc_hd__mux2_1 _40353_ (.A0(_02283_),
    .A1(_02281_),
    .S(_02217_),
    .X(_00024_));
 sky130_fd_sc_hd__mux2_1 _40354_ (.A0(_02284_),
    .A1(_02285_),
    .S(\irq_state[1] ),
    .X(_02286_));
 sky130_fd_sc_hd__mux2_1 _40355_ (.A0(_02286_),
    .A1(_02284_),
    .S(_02217_),
    .X(_00025_));
 sky130_fd_sc_hd__mux2_1 _40356_ (.A0(_02287_),
    .A1(_02288_),
    .S(\irq_state[1] ),
    .X(_02289_));
 sky130_fd_sc_hd__mux2_1 _40357_ (.A0(_02289_),
    .A1(_02287_),
    .S(_02217_),
    .X(_00026_));
 sky130_fd_sc_hd__mux2_1 _40358_ (.A0(_02290_),
    .A1(_02291_),
    .S(\irq_state[1] ),
    .X(_02292_));
 sky130_fd_sc_hd__mux2_1 _40359_ (.A0(_02292_),
    .A1(_02290_),
    .S(_02217_),
    .X(_00027_));
 sky130_fd_sc_hd__mux2_1 _40360_ (.A0(_02293_),
    .A1(_02294_),
    .S(\irq_state[1] ),
    .X(_02295_));
 sky130_fd_sc_hd__mux2_1 _40361_ (.A0(_02295_),
    .A1(_02293_),
    .S(_02217_),
    .X(_00028_));
 sky130_fd_sc_hd__mux2_1 _40362_ (.A0(_02296_),
    .A1(_02297_),
    .S(\irq_state[1] ),
    .X(_02298_));
 sky130_fd_sc_hd__mux2_1 _40363_ (.A0(_02298_),
    .A1(_02296_),
    .S(_02217_),
    .X(_00029_));
 sky130_fd_sc_hd__mux2_1 _40364_ (.A0(_02299_),
    .A1(_02300_),
    .S(\irq_state[1] ),
    .X(_02301_));
 sky130_fd_sc_hd__mux2_1 _40365_ (.A0(_02301_),
    .A1(_02299_),
    .S(_02217_),
    .X(_00030_));
 sky130_fd_sc_hd__mux2_1 _40366_ (.A0(_01467_),
    .A1(\reg_next_pc[1] ),
    .S(_00292_),
    .X(_02590_));
 sky130_fd_sc_hd__mux2_1 _40367_ (.A0(_00295_),
    .A1(\reg_next_pc[2] ),
    .S(_00292_),
    .X(_02560_));
 sky130_fd_sc_hd__mux2_1 _40368_ (.A0(_01470_),
    .A1(\reg_next_pc[3] ),
    .S(_00292_),
    .X(_02571_));
 sky130_fd_sc_hd__mux2_1 _40369_ (.A0(_01478_),
    .A1(\reg_next_pc[5] ),
    .S(_00292_),
    .X(_02583_));
 sky130_fd_sc_hd__mux2_1 _40370_ (.A0(_01481_),
    .A1(\reg_next_pc[6] ),
    .S(_00292_),
    .X(_02584_));
 sky130_fd_sc_hd__mux2_1 _40371_ (.A0(_01484_),
    .A1(\reg_next_pc[7] ),
    .S(_00292_),
    .X(_02585_));
 sky130_fd_sc_hd__mux2_1 _40372_ (.A0(_01487_),
    .A1(\reg_next_pc[8] ),
    .S(_00292_),
    .X(_02586_));
 sky130_fd_sc_hd__mux2_1 _40373_ (.A0(_01490_),
    .A1(\reg_next_pc[9] ),
    .S(_00292_),
    .X(_02587_));
 sky130_fd_sc_hd__mux2_1 _40374_ (.A0(_01493_),
    .A1(\reg_next_pc[10] ),
    .S(_00292_),
    .X(_02588_));
 sky130_fd_sc_hd__mux2_1 _40375_ (.A0(_01496_),
    .A1(\reg_next_pc[11] ),
    .S(_00292_),
    .X(_02589_));
 sky130_fd_sc_hd__mux2_1 _40376_ (.A0(_01499_),
    .A1(\reg_next_pc[12] ),
    .S(_00292_),
    .X(_02561_));
 sky130_fd_sc_hd__mux2_1 _40377_ (.A0(_01502_),
    .A1(\reg_next_pc[13] ),
    .S(_00292_),
    .X(_02562_));
 sky130_fd_sc_hd__mux2_1 _40378_ (.A0(_01505_),
    .A1(\reg_next_pc[14] ),
    .S(_00292_),
    .X(_02563_));
 sky130_fd_sc_hd__mux2_1 _40379_ (.A0(_01508_),
    .A1(\reg_next_pc[15] ),
    .S(_00292_),
    .X(_02564_));
 sky130_fd_sc_hd__mux2_1 _40380_ (.A0(_01511_),
    .A1(\reg_next_pc[16] ),
    .S(_00292_),
    .X(_02565_));
 sky130_fd_sc_hd__mux2_1 _40381_ (.A0(_01514_),
    .A1(\reg_next_pc[17] ),
    .S(_00292_),
    .X(_02566_));
 sky130_fd_sc_hd__mux2_1 _40382_ (.A0(_01517_),
    .A1(\reg_next_pc[18] ),
    .S(_00292_),
    .X(_02567_));
 sky130_fd_sc_hd__mux2_1 _40383_ (.A0(_01520_),
    .A1(\reg_next_pc[19] ),
    .S(_00292_),
    .X(_02568_));
 sky130_fd_sc_hd__mux2_1 _40384_ (.A0(_01523_),
    .A1(\reg_next_pc[20] ),
    .S(_00292_),
    .X(_02569_));
 sky130_fd_sc_hd__mux2_1 _40385_ (.A0(_01526_),
    .A1(\reg_next_pc[21] ),
    .S(_00292_),
    .X(_02570_));
 sky130_fd_sc_hd__mux2_1 _40386_ (.A0(_01529_),
    .A1(\reg_next_pc[22] ),
    .S(_00292_),
    .X(_02572_));
 sky130_fd_sc_hd__mux2_1 _40387_ (.A0(_01532_),
    .A1(\reg_next_pc[23] ),
    .S(_00292_),
    .X(_02573_));
 sky130_fd_sc_hd__mux2_1 _40388_ (.A0(_01535_),
    .A1(\reg_next_pc[24] ),
    .S(_00292_),
    .X(_02574_));
 sky130_fd_sc_hd__mux2_1 _40389_ (.A0(_01538_),
    .A1(\reg_next_pc[25] ),
    .S(_00292_),
    .X(_02575_));
 sky130_fd_sc_hd__mux2_1 _40390_ (.A0(_01541_),
    .A1(\reg_next_pc[26] ),
    .S(_00292_),
    .X(_02576_));
 sky130_fd_sc_hd__mux2_1 _40391_ (.A0(_01544_),
    .A1(\reg_next_pc[27] ),
    .S(_00292_),
    .X(_02577_));
 sky130_fd_sc_hd__mux2_1 _40392_ (.A0(_01547_),
    .A1(\reg_next_pc[28] ),
    .S(_00292_),
    .X(_02578_));
 sky130_fd_sc_hd__mux2_1 _40393_ (.A0(_01550_),
    .A1(\reg_next_pc[29] ),
    .S(_00292_),
    .X(_02579_));
 sky130_fd_sc_hd__mux2_1 _40394_ (.A0(_01553_),
    .A1(\reg_next_pc[30] ),
    .S(_00292_),
    .X(_02580_));
 sky130_fd_sc_hd__mux2_1 _40395_ (.A0(_01556_),
    .A1(\reg_next_pc[31] ),
    .S(_00292_),
    .X(_02581_));
 sky130_fd_sc_hd__mux2_1 _40396_ (.A0(_00057_),
    .A1(_00064_),
    .S(mem_la_wdata[3]),
    .X(_00065_));
 sky130_fd_sc_hd__mux2_1 _40397_ (.A0(_00065_),
    .A1(_02543_),
    .S(mem_la_wdata[4]),
    .X(_20623_));
 sky130_fd_sc_hd__mux2_1 _40398_ (.A0(_00075_),
    .A1(_00082_),
    .S(mem_la_wdata[3]),
    .X(_00083_));
 sky130_fd_sc_hd__mux2_1 _40399_ (.A0(_00083_),
    .A1(_02544_),
    .S(mem_la_wdata[4]),
    .X(_20624_));
 sky130_fd_sc_hd__mux2_1 _40400_ (.A0(_00089_),
    .A1(_00092_),
    .S(mem_la_wdata[3]),
    .X(_00093_));
 sky130_fd_sc_hd__mux2_1 _40401_ (.A0(_00093_),
    .A1(_02545_),
    .S(mem_la_wdata[4]),
    .X(_20625_));
 sky130_fd_sc_hd__mux2_1 _40402_ (.A0(_00099_),
    .A1(_00102_),
    .S(mem_la_wdata[3]),
    .X(_00103_));
 sky130_fd_sc_hd__mux2_1 _40403_ (.A0(_00103_),
    .A1(_02546_),
    .S(mem_la_wdata[4]),
    .X(_20626_));
 sky130_fd_sc_hd__mux2_1 _40404_ (.A0(_00107_),
    .A1(_00108_),
    .S(mem_la_wdata[3]),
    .X(_00109_));
 sky130_fd_sc_hd__mux2_1 _40405_ (.A0(_00109_),
    .A1(_02547_),
    .S(mem_la_wdata[4]),
    .X(_20627_));
 sky130_fd_sc_hd__mux2_1 _40406_ (.A0(_00113_),
    .A1(_00114_),
    .S(mem_la_wdata[3]),
    .X(_00115_));
 sky130_fd_sc_hd__mux2_1 _40407_ (.A0(_00115_),
    .A1(_02548_),
    .S(mem_la_wdata[4]),
    .X(_20628_));
 sky130_fd_sc_hd__mux2_1 _40408_ (.A0(_00119_),
    .A1(_00120_),
    .S(mem_la_wdata[3]),
    .X(_00121_));
 sky130_fd_sc_hd__mux2_1 _40409_ (.A0(_00121_),
    .A1(_02549_),
    .S(mem_la_wdata[4]),
    .X(_20629_));
 sky130_fd_sc_hd__mux2_1 _40410_ (.A0(_00125_),
    .A1(_00126_),
    .S(mem_la_wdata[3]),
    .X(_00127_));
 sky130_fd_sc_hd__mux2_1 _40411_ (.A0(_00127_),
    .A1(_02550_),
    .S(mem_la_wdata[4]),
    .X(_20630_));
 sky130_fd_sc_hd__mux2_1 _40412_ (.A0(_00129_),
    .A1(_00106_),
    .S(mem_la_wdata[2]),
    .X(_00130_));
 sky130_fd_sc_hd__mux2_1 _40413_ (.A0(_00130_),
    .A1(_00057_),
    .S(mem_la_wdata[3]),
    .X(_00131_));
 sky130_fd_sc_hd__mux2_1 _40414_ (.A0(_00131_),
    .A1(_02551_),
    .S(mem_la_wdata[4]),
    .X(_20631_));
 sky130_fd_sc_hd__mux2_1 _40415_ (.A0(_00133_),
    .A1(_00112_),
    .S(mem_la_wdata[2]),
    .X(_00134_));
 sky130_fd_sc_hd__mux2_1 _40416_ (.A0(_00134_),
    .A1(_00075_),
    .S(mem_la_wdata[3]),
    .X(_00135_));
 sky130_fd_sc_hd__mux2_1 _40417_ (.A0(_00135_),
    .A1(_02552_),
    .S(mem_la_wdata[4]),
    .X(_20632_));
 sky130_fd_sc_hd__mux2_1 _40418_ (.A0(_00137_),
    .A1(_00118_),
    .S(mem_la_wdata[2]),
    .X(_00138_));
 sky130_fd_sc_hd__mux2_1 _40419_ (.A0(_00138_),
    .A1(_00089_),
    .S(mem_la_wdata[3]),
    .X(_00139_));
 sky130_fd_sc_hd__mux2_1 _40420_ (.A0(_00139_),
    .A1(_02553_),
    .S(mem_la_wdata[4]),
    .X(_20633_));
 sky130_fd_sc_hd__mux2_1 _40421_ (.A0(_00141_),
    .A1(_00124_),
    .S(mem_la_wdata[2]),
    .X(_00142_));
 sky130_fd_sc_hd__mux2_1 _40422_ (.A0(_00142_),
    .A1(_00099_),
    .S(mem_la_wdata[3]),
    .X(_00143_));
 sky130_fd_sc_hd__mux2_1 _40423_ (.A0(_00143_),
    .A1(_02554_),
    .S(mem_la_wdata[4]),
    .X(_20634_));
 sky130_fd_sc_hd__mux2_1 _40424_ (.A0(_00144_),
    .A1(_00136_),
    .S(mem_la_wdata[1]),
    .X(_00145_));
 sky130_fd_sc_hd__mux2_1 _40425_ (.A0(_00145_),
    .A1(_00129_),
    .S(mem_la_wdata[2]),
    .X(_00146_));
 sky130_fd_sc_hd__mux2_1 _40426_ (.A0(_00146_),
    .A1(_00107_),
    .S(mem_la_wdata[3]),
    .X(_00147_));
 sky130_fd_sc_hd__mux2_1 _40427_ (.A0(_00147_),
    .A1(_02555_),
    .S(mem_la_wdata[4]),
    .X(_20635_));
 sky130_fd_sc_hd__mux2_1 _40428_ (.A0(_00148_),
    .A1(_00140_),
    .S(mem_la_wdata[1]),
    .X(_00149_));
 sky130_fd_sc_hd__mux2_1 _40429_ (.A0(_00149_),
    .A1(_00133_),
    .S(mem_la_wdata[2]),
    .X(_00150_));
 sky130_fd_sc_hd__mux2_1 _40430_ (.A0(_00150_),
    .A1(_00113_),
    .S(mem_la_wdata[3]),
    .X(_00151_));
 sky130_fd_sc_hd__mux2_1 _40431_ (.A0(_00151_),
    .A1(_02556_),
    .S(mem_la_wdata[4]),
    .X(_20636_));
 sky130_fd_sc_hd__mux2_1 _40432_ (.A0(pcpi_rs1[30]),
    .A1(pcpi_rs1[29]),
    .S(mem_la_wdata[0]),
    .X(_00152_));
 sky130_fd_sc_hd__mux2_1 _40433_ (.A0(_00152_),
    .A1(_00144_),
    .S(mem_la_wdata[1]),
    .X(_00153_));
 sky130_fd_sc_hd__mux2_1 _40434_ (.A0(_00153_),
    .A1(_00137_),
    .S(mem_la_wdata[2]),
    .X(_00154_));
 sky130_fd_sc_hd__mux2_1 _40435_ (.A0(_00154_),
    .A1(_00119_),
    .S(mem_la_wdata[3]),
    .X(_00155_));
 sky130_fd_sc_hd__mux2_1 _40436_ (.A0(_00155_),
    .A1(_02557_),
    .S(mem_la_wdata[4]),
    .X(_20637_));
 sky130_fd_sc_hd__mux2_1 _40437_ (.A0(pcpi_rs1[31]),
    .A1(pcpi_rs1[30]),
    .S(mem_la_wdata[0]),
    .X(_00156_));
 sky130_fd_sc_hd__mux2_1 _40438_ (.A0(_00156_),
    .A1(_00148_),
    .S(mem_la_wdata[1]),
    .X(_00157_));
 sky130_fd_sc_hd__mux2_1 _40439_ (.A0(_00157_),
    .A1(_00141_),
    .S(mem_la_wdata[2]),
    .X(_00158_));
 sky130_fd_sc_hd__mux2_1 _40440_ (.A0(_00158_),
    .A1(_00125_),
    .S(mem_la_wdata[3]),
    .X(_00159_));
 sky130_fd_sc_hd__mux2_1 _40441_ (.A0(_00159_),
    .A1(_02558_),
    .S(mem_la_wdata[4]),
    .X(_20638_));
 sky130_fd_sc_hd__mux2_1 _40442_ (.A0(pcpi_rs1[0]),
    .A1(pcpi_rs1[1]),
    .S(mem_la_wdata[0]),
    .X(_00160_));
 sky130_fd_sc_hd__mux2_1 _40443_ (.A0(_00160_),
    .A1(_00161_),
    .S(mem_la_wdata[1]),
    .X(_00162_));
 sky130_fd_sc_hd__mux2_1 _40444_ (.A0(_00162_),
    .A1(_00165_),
    .S(mem_la_wdata[2]),
    .X(_00166_));
 sky130_fd_sc_hd__mux2_1 _40445_ (.A0(_00166_),
    .A1(_00173_),
    .S(mem_la_wdata[3]),
    .X(_00174_));
 sky130_fd_sc_hd__mux2_1 _40446_ (.A0(_00174_),
    .A1(_00189_),
    .S(mem_la_wdata[4]),
    .X(_20639_));
 sky130_fd_sc_hd__mux2_1 _40447_ (.A0(pcpi_rs1[1]),
    .A1(pcpi_rs1[2]),
    .S(mem_la_wdata[0]),
    .X(_00190_));
 sky130_fd_sc_hd__mux2_1 _40448_ (.A0(_00190_),
    .A1(_00191_),
    .S(mem_la_wdata[1]),
    .X(_00192_));
 sky130_fd_sc_hd__mux2_1 _40449_ (.A0(_00192_),
    .A1(_00195_),
    .S(mem_la_wdata[2]),
    .X(_00196_));
 sky130_fd_sc_hd__mux2_1 _40450_ (.A0(_00196_),
    .A1(_00203_),
    .S(mem_la_wdata[3]),
    .X(_00204_));
 sky130_fd_sc_hd__mux2_1 _40451_ (.A0(_00204_),
    .A1(_00220_),
    .S(mem_la_wdata[4]),
    .X(_20650_));
 sky130_fd_sc_hd__mux2_1 _40452_ (.A0(_00161_),
    .A1(_00163_),
    .S(mem_la_wdata[1]),
    .X(_00221_));
 sky130_fd_sc_hd__mux2_1 _40453_ (.A0(_00221_),
    .A1(_00222_),
    .S(mem_la_wdata[2]),
    .X(_00223_));
 sky130_fd_sc_hd__mux2_1 _40454_ (.A0(_00223_),
    .A1(_00226_),
    .S(mem_la_wdata[3]),
    .X(_00227_));
 sky130_fd_sc_hd__mux2_1 _40455_ (.A0(_00227_),
    .A1(_00234_),
    .S(mem_la_wdata[4]),
    .X(_20661_));
 sky130_fd_sc_hd__mux2_1 _40456_ (.A0(_00191_),
    .A1(_00193_),
    .S(mem_la_wdata[1]),
    .X(_00235_));
 sky130_fd_sc_hd__mux2_1 _40457_ (.A0(_00235_),
    .A1(_00236_),
    .S(mem_la_wdata[2]),
    .X(_00237_));
 sky130_fd_sc_hd__mux2_1 _40458_ (.A0(_00237_),
    .A1(_00240_),
    .S(mem_la_wdata[3]),
    .X(_00241_));
 sky130_fd_sc_hd__mux2_1 _40459_ (.A0(_00241_),
    .A1(_00248_),
    .S(mem_la_wdata[4]),
    .X(_20664_));
 sky130_fd_sc_hd__mux2_1 _40460_ (.A0(_00165_),
    .A1(_00169_),
    .S(mem_la_wdata[2]),
    .X(_00249_));
 sky130_fd_sc_hd__mux2_1 _40461_ (.A0(_00249_),
    .A1(_00250_),
    .S(mem_la_wdata[3]),
    .X(_00251_));
 sky130_fd_sc_hd__mux2_1 _40462_ (.A0(_00251_),
    .A1(_00254_),
    .S(mem_la_wdata[4]),
    .X(_20665_));
 sky130_fd_sc_hd__mux2_1 _40463_ (.A0(_00195_),
    .A1(_00199_),
    .S(mem_la_wdata[2]),
    .X(_00255_));
 sky130_fd_sc_hd__mux2_1 _40464_ (.A0(_00255_),
    .A1(_00256_),
    .S(mem_la_wdata[3]),
    .X(_00257_));
 sky130_fd_sc_hd__mux2_1 _40465_ (.A0(_00257_),
    .A1(_00260_),
    .S(mem_la_wdata[4]),
    .X(_20666_));
 sky130_fd_sc_hd__mux2_1 _40466_ (.A0(_00222_),
    .A1(_00224_),
    .S(mem_la_wdata[2]),
    .X(_00261_));
 sky130_fd_sc_hd__mux2_1 _40467_ (.A0(_00261_),
    .A1(_00262_),
    .S(mem_la_wdata[3]),
    .X(_00263_));
 sky130_fd_sc_hd__mux2_1 _40468_ (.A0(_00263_),
    .A1(_00266_),
    .S(mem_la_wdata[4]),
    .X(_20667_));
 sky130_fd_sc_hd__mux2_1 _40469_ (.A0(_00236_),
    .A1(_00238_),
    .S(mem_la_wdata[2]),
    .X(_00267_));
 sky130_fd_sc_hd__mux2_1 _40470_ (.A0(_00267_),
    .A1(_00268_),
    .S(mem_la_wdata[3]),
    .X(_00269_));
 sky130_fd_sc_hd__mux2_1 _40471_ (.A0(_00269_),
    .A1(_00272_),
    .S(mem_la_wdata[4]),
    .X(_20668_));
 sky130_fd_sc_hd__mux2_1 _40472_ (.A0(_00173_),
    .A1(_00181_),
    .S(mem_la_wdata[3]),
    .X(_00273_));
 sky130_fd_sc_hd__mux2_1 _40473_ (.A0(_00273_),
    .A1(_00274_),
    .S(mem_la_wdata[4]),
    .X(_20669_));
 sky130_fd_sc_hd__mux2_1 _40474_ (.A0(_00203_),
    .A1(_00211_),
    .S(mem_la_wdata[3]),
    .X(_00275_));
 sky130_fd_sc_hd__mux2_1 _40475_ (.A0(_00275_),
    .A1(_00276_),
    .S(mem_la_wdata[4]),
    .X(_20670_));
 sky130_fd_sc_hd__mux2_1 _40476_ (.A0(_00226_),
    .A1(_00230_),
    .S(mem_la_wdata[3]),
    .X(_00277_));
 sky130_fd_sc_hd__mux2_1 _40477_ (.A0(_00277_),
    .A1(_00278_),
    .S(mem_la_wdata[4]),
    .X(_20640_));
 sky130_fd_sc_hd__mux2_1 _40478_ (.A0(_00240_),
    .A1(_00244_),
    .S(mem_la_wdata[3]),
    .X(_00279_));
 sky130_fd_sc_hd__mux2_1 _40479_ (.A0(_00279_),
    .A1(_00280_),
    .S(mem_la_wdata[4]),
    .X(_20641_));
 sky130_fd_sc_hd__mux2_1 _40480_ (.A0(_00250_),
    .A1(_00252_),
    .S(mem_la_wdata[3]),
    .X(_00281_));
 sky130_fd_sc_hd__mux2_1 _40481_ (.A0(_00281_),
    .A1(_00282_),
    .S(mem_la_wdata[4]),
    .X(_20642_));
 sky130_fd_sc_hd__mux2_1 _40482_ (.A0(_00256_),
    .A1(_00258_),
    .S(mem_la_wdata[3]),
    .X(_00283_));
 sky130_fd_sc_hd__mux2_1 _40483_ (.A0(_00283_),
    .A1(_00284_),
    .S(mem_la_wdata[4]),
    .X(_20643_));
 sky130_fd_sc_hd__mux2_1 _40484_ (.A0(_00262_),
    .A1(_00264_),
    .S(mem_la_wdata[3]),
    .X(_00285_));
 sky130_fd_sc_hd__mux2_1 _40485_ (.A0(_00285_),
    .A1(_00286_),
    .S(mem_la_wdata[4]),
    .X(_20644_));
 sky130_fd_sc_hd__mux2_1 _40486_ (.A0(_00268_),
    .A1(_00270_),
    .S(mem_la_wdata[3]),
    .X(_00287_));
 sky130_fd_sc_hd__mux2_1 _40487_ (.A0(_00287_),
    .A1(_00288_),
    .S(mem_la_wdata[4]),
    .X(_20645_));
 sky130_fd_sc_hd__mux2_1 _40488_ (.A0(_00189_),
    .A1(_00216_),
    .S(mem_la_wdata[4]),
    .X(_20646_));
 sky130_fd_sc_hd__mux2_1 _40489_ (.A0(_00220_),
    .A1(_00216_),
    .S(mem_la_wdata[4]),
    .X(_20647_));
 sky130_fd_sc_hd__mux2_1 _40490_ (.A0(_00234_),
    .A1(_00216_),
    .S(mem_la_wdata[4]),
    .X(_20648_));
 sky130_fd_sc_hd__mux2_1 _40491_ (.A0(_00248_),
    .A1(_00216_),
    .S(mem_la_wdata[4]),
    .X(_20649_));
 sky130_fd_sc_hd__mux2_1 _40492_ (.A0(_00254_),
    .A1(_00216_),
    .S(mem_la_wdata[4]),
    .X(_20651_));
 sky130_fd_sc_hd__mux2_1 _40493_ (.A0(_00260_),
    .A1(_00216_),
    .S(mem_la_wdata[4]),
    .X(_20652_));
 sky130_fd_sc_hd__mux2_1 _40494_ (.A0(_00266_),
    .A1(_00216_),
    .S(mem_la_wdata[4]),
    .X(_20653_));
 sky130_fd_sc_hd__mux2_1 _40495_ (.A0(_00272_),
    .A1(_00216_),
    .S(mem_la_wdata[4]),
    .X(_20654_));
 sky130_fd_sc_hd__mux2_1 _40496_ (.A0(_00274_),
    .A1(_00216_),
    .S(mem_la_wdata[4]),
    .X(_20655_));
 sky130_fd_sc_hd__mux2_1 _40497_ (.A0(_00276_),
    .A1(_00216_),
    .S(mem_la_wdata[4]),
    .X(_20656_));
 sky130_fd_sc_hd__mux2_1 _40498_ (.A0(_00278_),
    .A1(_00216_),
    .S(mem_la_wdata[4]),
    .X(_20657_));
 sky130_fd_sc_hd__mux2_1 _40499_ (.A0(_00280_),
    .A1(_00216_),
    .S(mem_la_wdata[4]),
    .X(_20658_));
 sky130_fd_sc_hd__mux2_1 _40500_ (.A0(_00282_),
    .A1(_00216_),
    .S(mem_la_wdata[4]),
    .X(_20659_));
 sky130_fd_sc_hd__mux2_1 _40501_ (.A0(_00284_),
    .A1(_00216_),
    .S(mem_la_wdata[4]),
    .X(_20660_));
 sky130_fd_sc_hd__mux2_1 _40502_ (.A0(_00286_),
    .A1(_00216_),
    .S(mem_la_wdata[4]),
    .X(_20662_));
 sky130_fd_sc_hd__mux2_1 _40503_ (.A0(_00288_),
    .A1(_00216_),
    .S(mem_la_wdata[4]),
    .X(_20663_));
 sky130_fd_sc_hd__mux2_1 _40504_ (.A0(_01697_),
    .A1(_01698_),
    .S(\irq_state[1] ),
    .X(_01699_));
 sky130_fd_sc_hd__mux2_1 _40505_ (.A0(_01705_),
    .A1(_01699_),
    .S(_01700_),
    .X(_20622_));
 sky130_fd_sc_hd__mux2_1 _40506_ (.A0(_01720_),
    .A1(\irq_pending[0] ),
    .S(_01706_),
    .X(_20588_));
 sky130_fd_sc_hd__mux2_1 _40507_ (.A0(_01733_),
    .A1(\irq_pending[1] ),
    .S(_01706_),
    .X(_20599_));
 sky130_fd_sc_hd__mux2_1 _40508_ (.A0(_01746_),
    .A1(\irq_pending[2] ),
    .S(_01706_),
    .X(_20610_));
 sky130_fd_sc_hd__mux2_1 _40509_ (.A0(_01759_),
    .A1(\irq_pending[3] ),
    .S(_01706_),
    .X(_20613_));
 sky130_fd_sc_hd__mux2_1 _40510_ (.A0(_01772_),
    .A1(\irq_pending[4] ),
    .S(_01706_),
    .X(_20614_));
 sky130_fd_sc_hd__mux2_1 _40511_ (.A0(_01785_),
    .A1(\irq_pending[5] ),
    .S(_01706_),
    .X(_20615_));
 sky130_fd_sc_hd__mux2_1 _40512_ (.A0(_01798_),
    .A1(\irq_pending[6] ),
    .S(_01706_),
    .X(_20616_));
 sky130_fd_sc_hd__mux2_1 _40513_ (.A0(_01811_),
    .A1(\irq_pending[7] ),
    .S(_01706_),
    .X(_20617_));
 sky130_fd_sc_hd__mux2_1 _40514_ (.A0(_01825_),
    .A1(\irq_pending[8] ),
    .S(_01706_),
    .X(_20618_));
 sky130_fd_sc_hd__mux2_1 _40515_ (.A0(_01838_),
    .A1(\irq_pending[9] ),
    .S(_01706_),
    .X(_20619_));
 sky130_fd_sc_hd__mux2_1 _40516_ (.A0(_01851_),
    .A1(\irq_pending[10] ),
    .S(_01706_),
    .X(_20589_));
 sky130_fd_sc_hd__mux2_1 _40517_ (.A0(_01864_),
    .A1(\irq_pending[11] ),
    .S(_01706_),
    .X(_20590_));
 sky130_fd_sc_hd__mux2_1 _40518_ (.A0(_01877_),
    .A1(\irq_pending[12] ),
    .S(_01706_),
    .X(_20591_));
 sky130_fd_sc_hd__mux2_1 _40519_ (.A0(_01890_),
    .A1(\irq_pending[13] ),
    .S(_01706_),
    .X(_20592_));
 sky130_fd_sc_hd__mux2_1 _40520_ (.A0(_01903_),
    .A1(\irq_pending[14] ),
    .S(_01706_),
    .X(_20593_));
 sky130_fd_sc_hd__mux2_1 _40521_ (.A0(_01916_),
    .A1(\irq_pending[15] ),
    .S(_01706_),
    .X(_20594_));
 sky130_fd_sc_hd__mux2_1 _40522_ (.A0(_01925_),
    .A1(\irq_pending[16] ),
    .S(_01706_),
    .X(_20595_));
 sky130_fd_sc_hd__mux2_1 _40523_ (.A0(_01934_),
    .A1(\irq_pending[17] ),
    .S(_01706_),
    .X(_20596_));
 sky130_fd_sc_hd__mux2_1 _40524_ (.A0(_01943_),
    .A1(\irq_pending[18] ),
    .S(_01706_),
    .X(_20597_));
 sky130_fd_sc_hd__mux2_1 _40525_ (.A0(_01952_),
    .A1(\irq_pending[19] ),
    .S(_01706_),
    .X(_20598_));
 sky130_fd_sc_hd__mux2_1 _40526_ (.A0(_01961_),
    .A1(\irq_pending[20] ),
    .S(_01706_),
    .X(_20600_));
 sky130_fd_sc_hd__mux2_1 _40527_ (.A0(_01970_),
    .A1(\irq_pending[21] ),
    .S(_01706_),
    .X(_20601_));
 sky130_fd_sc_hd__mux2_1 _40528_ (.A0(_01979_),
    .A1(\irq_pending[22] ),
    .S(_01706_),
    .X(_20602_));
 sky130_fd_sc_hd__mux2_1 _40529_ (.A0(_01988_),
    .A1(\irq_pending[23] ),
    .S(_01706_),
    .X(_20603_));
 sky130_fd_sc_hd__mux2_1 _40530_ (.A0(_01997_),
    .A1(\irq_pending[24] ),
    .S(_01706_),
    .X(_20604_));
 sky130_fd_sc_hd__mux2_1 _40531_ (.A0(_02006_),
    .A1(\irq_pending[25] ),
    .S(_01706_),
    .X(_20605_));
 sky130_fd_sc_hd__mux2_1 _40532_ (.A0(_02015_),
    .A1(\irq_pending[26] ),
    .S(_01706_),
    .X(_20606_));
 sky130_fd_sc_hd__mux2_1 _40533_ (.A0(_02024_),
    .A1(\irq_pending[27] ),
    .S(_01706_),
    .X(_20607_));
 sky130_fd_sc_hd__mux2_1 _40534_ (.A0(_02033_),
    .A1(\irq_pending[28] ),
    .S(_01706_),
    .X(_20608_));
 sky130_fd_sc_hd__mux2_1 _40535_ (.A0(_02042_),
    .A1(\irq_pending[29] ),
    .S(_01706_),
    .X(_20609_));
 sky130_fd_sc_hd__mux2_1 _40536_ (.A0(_02051_),
    .A1(\irq_pending[30] ),
    .S(_01706_),
    .X(_20611_));
 sky130_fd_sc_hd__mux2_1 _40537_ (.A0(_02060_),
    .A1(\irq_pending[31] ),
    .S(_01706_),
    .X(_20612_));
 sky130_fd_sc_hd__mux2_1 _40538_ (.A0(_02061_),
    .A1(\cpu_state[2] ),
    .S(_02542_),
    .X(_20583_));
 sky130_fd_sc_hd__mux2_1 _40539_ (.A0(\decoded_rd[0] ),
    .A1(\irq_state[0] ),
    .S(_00308_),
    .X(_20582_));
 sky130_fd_sc_hd__mux2_1 _40540_ (.A0(_02062_),
    .A1(_02065_),
    .S(_02542_),
    .X(_20620_));
 sky130_fd_sc_hd__mux2_1 _40541_ (.A0(_02068_),
    .A1(_02066_),
    .S(_02067_),
    .X(_20621_));
 sky130_fd_sc_hd__mux2_1 _40542_ (.A0(_02166_),
    .A1(_00291_),
    .S(_00290_),
    .X(_20584_));
 sky130_fd_sc_hd__mux2_1 _40543_ (.A0(_02166_),
    .A1(mem_do_wdata),
    .S(_00290_),
    .X(_20585_));
 sky130_fd_sc_hd__mux2_1 _40544_ (.A0(_00271_),
    .A1(_00216_),
    .S(mem_la_wdata[3]),
    .X(_00288_));
 sky130_fd_sc_hd__mux2_1 _40545_ (.A0(_00265_),
    .A1(_00216_),
    .S(mem_la_wdata[3]),
    .X(_00286_));
 sky130_fd_sc_hd__mux2_1 _40546_ (.A0(_00259_),
    .A1(_00216_),
    .S(mem_la_wdata[3]),
    .X(_00284_));
 sky130_fd_sc_hd__mux2_1 _40547_ (.A0(_00253_),
    .A1(_00216_),
    .S(mem_la_wdata[3]),
    .X(_00282_));
 sky130_fd_sc_hd__mux2_1 _40548_ (.A0(_00247_),
    .A1(_00216_),
    .S(mem_la_wdata[3]),
    .X(_00280_));
 sky130_fd_sc_hd__mux2_1 _40549_ (.A0(_00233_),
    .A1(_00216_),
    .S(mem_la_wdata[3]),
    .X(_00278_));
 sky130_fd_sc_hd__mux2_1 _40550_ (.A0(_00219_),
    .A1(_00216_),
    .S(mem_la_wdata[3]),
    .X(_00276_));
 sky130_fd_sc_hd__mux2_1 _40551_ (.A0(_00188_),
    .A1(_00216_),
    .S(mem_la_wdata[3]),
    .X(_00274_));
 sky130_fd_sc_hd__mux2_1 _40552_ (.A0(_00270_),
    .A1(_00271_),
    .S(mem_la_wdata[3]),
    .X(_00272_));
 sky130_fd_sc_hd__mux2_1 _40553_ (.A0(_00246_),
    .A1(_00216_),
    .S(mem_la_wdata[2]),
    .X(_00271_));
 sky130_fd_sc_hd__mux2_1 _40554_ (.A0(_00243_),
    .A1(_00245_),
    .S(mem_la_wdata[2]),
    .X(_00270_));
 sky130_fd_sc_hd__mux2_1 _40555_ (.A0(_00239_),
    .A1(_00242_),
    .S(mem_la_wdata[2]),
    .X(_00268_));
 sky130_fd_sc_hd__mux2_1 _40556_ (.A0(_00264_),
    .A1(_00265_),
    .S(mem_la_wdata[3]),
    .X(_00266_));
 sky130_fd_sc_hd__mux2_1 _40557_ (.A0(_00232_),
    .A1(_00216_),
    .S(mem_la_wdata[2]),
    .X(_00265_));
 sky130_fd_sc_hd__mux2_1 _40558_ (.A0(_00229_),
    .A1(_00231_),
    .S(mem_la_wdata[2]),
    .X(_00264_));
 sky130_fd_sc_hd__mux2_1 _40559_ (.A0(_00225_),
    .A1(_00228_),
    .S(mem_la_wdata[2]),
    .X(_00262_));
 sky130_fd_sc_hd__mux2_1 _40560_ (.A0(_00258_),
    .A1(_00259_),
    .S(mem_la_wdata[3]),
    .X(_00260_));
 sky130_fd_sc_hd__mux2_1 _40561_ (.A0(_00218_),
    .A1(_00216_),
    .S(mem_la_wdata[2]),
    .X(_00259_));
 sky130_fd_sc_hd__mux2_1 _40562_ (.A0(_00210_),
    .A1(_00214_),
    .S(mem_la_wdata[2]),
    .X(_00258_));
 sky130_fd_sc_hd__mux2_1 _40563_ (.A0(_00202_),
    .A1(_00207_),
    .S(mem_la_wdata[2]),
    .X(_00256_));
 sky130_fd_sc_hd__mux2_1 _40564_ (.A0(_00252_),
    .A1(_00253_),
    .S(mem_la_wdata[3]),
    .X(_00254_));
 sky130_fd_sc_hd__mux2_1 _40565_ (.A0(_00187_),
    .A1(_00216_),
    .S(mem_la_wdata[2]),
    .X(_00253_));
 sky130_fd_sc_hd__mux2_1 _40566_ (.A0(_00180_),
    .A1(_00184_),
    .S(mem_la_wdata[2]),
    .X(_00252_));
 sky130_fd_sc_hd__mux2_1 _40567_ (.A0(_00172_),
    .A1(_00177_),
    .S(mem_la_wdata[2]),
    .X(_00250_));
 sky130_fd_sc_hd__mux2_1 _40568_ (.A0(_00244_),
    .A1(_00247_),
    .S(mem_la_wdata[3]),
    .X(_00248_));
 sky130_fd_sc_hd__mux2_1 _40569_ (.A0(_00245_),
    .A1(_00246_),
    .S(mem_la_wdata[2]),
    .X(_00247_));
 sky130_fd_sc_hd__mux2_1 _40570_ (.A0(_00217_),
    .A1(_00216_),
    .S(mem_la_wdata[1]),
    .X(_00246_));
 sky130_fd_sc_hd__mux2_1 _40571_ (.A0(_00213_),
    .A1(_00215_),
    .S(mem_la_wdata[1]),
    .X(_00245_));
 sky130_fd_sc_hd__mux2_1 _40572_ (.A0(_00242_),
    .A1(_00243_),
    .S(mem_la_wdata[2]),
    .X(_00244_));
 sky130_fd_sc_hd__mux2_1 _40573_ (.A0(_00209_),
    .A1(_00212_),
    .S(mem_la_wdata[1]),
    .X(_00243_));
 sky130_fd_sc_hd__mux2_1 _40574_ (.A0(_00206_),
    .A1(_00208_),
    .S(mem_la_wdata[1]),
    .X(_00242_));
 sky130_fd_sc_hd__mux2_1 _40575_ (.A0(_00238_),
    .A1(_00239_),
    .S(mem_la_wdata[2]),
    .X(_00240_));
 sky130_fd_sc_hd__mux2_1 _40576_ (.A0(_00201_),
    .A1(_00205_),
    .S(mem_la_wdata[1]),
    .X(_00239_));
 sky130_fd_sc_hd__mux2_1 _40577_ (.A0(_00198_),
    .A1(_00200_),
    .S(mem_la_wdata[1]),
    .X(_00238_));
 sky130_fd_sc_hd__mux2_1 _40578_ (.A0(_00194_),
    .A1(_00197_),
    .S(mem_la_wdata[1]),
    .X(_00236_));
 sky130_fd_sc_hd__mux2_1 _40579_ (.A0(_00230_),
    .A1(_00233_),
    .S(mem_la_wdata[3]),
    .X(_00234_));
 sky130_fd_sc_hd__mux2_1 _40580_ (.A0(_00231_),
    .A1(_00232_),
    .S(mem_la_wdata[2]),
    .X(_00233_));
 sky130_fd_sc_hd__mux2_1 _40581_ (.A0(_00186_),
    .A1(_00216_),
    .S(mem_la_wdata[1]),
    .X(_00232_));
 sky130_fd_sc_hd__mux2_1 _40582_ (.A0(_00183_),
    .A1(_00185_),
    .S(mem_la_wdata[1]),
    .X(_00231_));
 sky130_fd_sc_hd__mux2_1 _40583_ (.A0(_00228_),
    .A1(_00229_),
    .S(mem_la_wdata[2]),
    .X(_00230_));
 sky130_fd_sc_hd__mux2_1 _40584_ (.A0(_00179_),
    .A1(_00182_),
    .S(mem_la_wdata[1]),
    .X(_00229_));
 sky130_fd_sc_hd__mux2_1 _40585_ (.A0(_00176_),
    .A1(_00178_),
    .S(mem_la_wdata[1]),
    .X(_00228_));
 sky130_fd_sc_hd__mux2_1 _40586_ (.A0(_00224_),
    .A1(_00225_),
    .S(mem_la_wdata[2]),
    .X(_00226_));
 sky130_fd_sc_hd__mux2_1 _40587_ (.A0(_00171_),
    .A1(_00175_),
    .S(mem_la_wdata[1]),
    .X(_00225_));
 sky130_fd_sc_hd__mux2_1 _40588_ (.A0(_00168_),
    .A1(_00170_),
    .S(mem_la_wdata[1]),
    .X(_00224_));
 sky130_fd_sc_hd__mux2_1 _40589_ (.A0(_00164_),
    .A1(_00167_),
    .S(mem_la_wdata[1]),
    .X(_00222_));
 sky130_fd_sc_hd__mux2_1 _40590_ (.A0(_00211_),
    .A1(_00219_),
    .S(mem_la_wdata[3]),
    .X(_00220_));
 sky130_fd_sc_hd__mux2_1 _40591_ (.A0(_00214_),
    .A1(_00218_),
    .S(mem_la_wdata[2]),
    .X(_00219_));
 sky130_fd_sc_hd__mux2_1 _40592_ (.A0(_00215_),
    .A1(_00217_),
    .S(mem_la_wdata[1]),
    .X(_00218_));
 sky130_fd_sc_hd__mux2_1 _40593_ (.A0(pcpi_rs1[31]),
    .A1(_00216_),
    .S(mem_la_wdata[0]),
    .X(_00217_));
 sky130_fd_sc_hd__mux2_1 _40594_ (.A0(pcpi_rs1[29]),
    .A1(pcpi_rs1[30]),
    .S(mem_la_wdata[0]),
    .X(_00215_));
 sky130_fd_sc_hd__mux2_1 _40595_ (.A0(_00212_),
    .A1(_00213_),
    .S(mem_la_wdata[1]),
    .X(_00214_));
 sky130_fd_sc_hd__mux2_1 _40596_ (.A0(pcpi_rs1[27]),
    .A1(pcpi_rs1[28]),
    .S(mem_la_wdata[0]),
    .X(_00213_));
 sky130_fd_sc_hd__mux2_1 _40597_ (.A0(pcpi_rs1[25]),
    .A1(pcpi_rs1[26]),
    .S(mem_la_wdata[0]),
    .X(_00212_));
 sky130_fd_sc_hd__mux2_1 _40598_ (.A0(_00207_),
    .A1(_00210_),
    .S(mem_la_wdata[2]),
    .X(_00211_));
 sky130_fd_sc_hd__mux2_1 _40599_ (.A0(_00208_),
    .A1(_00209_),
    .S(mem_la_wdata[1]),
    .X(_00210_));
 sky130_fd_sc_hd__mux2_1 _40600_ (.A0(pcpi_rs1[23]),
    .A1(pcpi_rs1[24]),
    .S(mem_la_wdata[0]),
    .X(_00209_));
 sky130_fd_sc_hd__mux2_1 _40601_ (.A0(pcpi_rs1[21]),
    .A1(pcpi_rs1[22]),
    .S(mem_la_wdata[0]),
    .X(_00208_));
 sky130_fd_sc_hd__mux2_1 _40602_ (.A0(_00205_),
    .A1(_00206_),
    .S(mem_la_wdata[1]),
    .X(_00207_));
 sky130_fd_sc_hd__mux2_1 _40603_ (.A0(pcpi_rs1[19]),
    .A1(pcpi_rs1[20]),
    .S(mem_la_wdata[0]),
    .X(_00206_));
 sky130_fd_sc_hd__mux2_1 _40604_ (.A0(pcpi_rs1[17]),
    .A1(pcpi_rs1[18]),
    .S(mem_la_wdata[0]),
    .X(_00205_));
 sky130_fd_sc_hd__mux2_1 _40605_ (.A0(_00199_),
    .A1(_00202_),
    .S(mem_la_wdata[2]),
    .X(_00203_));
 sky130_fd_sc_hd__mux2_1 _40606_ (.A0(_00200_),
    .A1(_00201_),
    .S(mem_la_wdata[1]),
    .X(_00202_));
 sky130_fd_sc_hd__mux2_1 _40607_ (.A0(pcpi_rs1[15]),
    .A1(pcpi_rs1[16]),
    .S(mem_la_wdata[0]),
    .X(_00201_));
 sky130_fd_sc_hd__mux2_1 _40608_ (.A0(pcpi_rs1[13]),
    .A1(pcpi_rs1[14]),
    .S(mem_la_wdata[0]),
    .X(_00200_));
 sky130_fd_sc_hd__mux2_1 _40609_ (.A0(_00197_),
    .A1(_00198_),
    .S(mem_la_wdata[1]),
    .X(_00199_));
 sky130_fd_sc_hd__mux2_1 _40610_ (.A0(pcpi_rs1[11]),
    .A1(pcpi_rs1[12]),
    .S(mem_la_wdata[0]),
    .X(_00198_));
 sky130_fd_sc_hd__mux2_1 _40611_ (.A0(pcpi_rs1[9]),
    .A1(pcpi_rs1[10]),
    .S(mem_la_wdata[0]),
    .X(_00197_));
 sky130_fd_sc_hd__mux2_1 _40612_ (.A0(_00193_),
    .A1(_00194_),
    .S(mem_la_wdata[1]),
    .X(_00195_));
 sky130_fd_sc_hd__mux2_1 _40613_ (.A0(pcpi_rs1[7]),
    .A1(pcpi_rs1[8]),
    .S(mem_la_wdata[0]),
    .X(_00194_));
 sky130_fd_sc_hd__mux2_1 _40614_ (.A0(pcpi_rs1[5]),
    .A1(pcpi_rs1[6]),
    .S(mem_la_wdata[0]),
    .X(_00193_));
 sky130_fd_sc_hd__mux2_1 _40615_ (.A0(pcpi_rs1[3]),
    .A1(pcpi_rs1[4]),
    .S(mem_la_wdata[0]),
    .X(_00191_));
 sky130_fd_sc_hd__mux2_1 _40616_ (.A0(_00181_),
    .A1(_00188_),
    .S(mem_la_wdata[3]),
    .X(_00189_));
 sky130_fd_sc_hd__mux2_1 _40617_ (.A0(_00184_),
    .A1(_00187_),
    .S(mem_la_wdata[2]),
    .X(_00188_));
 sky130_fd_sc_hd__mux2_1 _40618_ (.A0(_00185_),
    .A1(_00186_),
    .S(mem_la_wdata[1]),
    .X(_00187_));
 sky130_fd_sc_hd__mux2_1 _40619_ (.A0(pcpi_rs1[30]),
    .A1(pcpi_rs1[31]),
    .S(mem_la_wdata[0]),
    .X(_00186_));
 sky130_fd_sc_hd__mux2_1 _40620_ (.A0(pcpi_rs1[28]),
    .A1(pcpi_rs1[29]),
    .S(mem_la_wdata[0]),
    .X(_00185_));
 sky130_fd_sc_hd__mux2_1 _40621_ (.A0(_00182_),
    .A1(_00183_),
    .S(mem_la_wdata[1]),
    .X(_00184_));
 sky130_fd_sc_hd__mux2_1 _40622_ (.A0(pcpi_rs1[26]),
    .A1(pcpi_rs1[27]),
    .S(mem_la_wdata[0]),
    .X(_00183_));
 sky130_fd_sc_hd__mux2_1 _40623_ (.A0(pcpi_rs1[24]),
    .A1(pcpi_rs1[25]),
    .S(mem_la_wdata[0]),
    .X(_00182_));
 sky130_fd_sc_hd__mux2_1 _40624_ (.A0(_00177_),
    .A1(_00180_),
    .S(mem_la_wdata[2]),
    .X(_00181_));
 sky130_fd_sc_hd__mux2_1 _40625_ (.A0(_00178_),
    .A1(_00179_),
    .S(mem_la_wdata[1]),
    .X(_00180_));
 sky130_fd_sc_hd__mux2_1 _40626_ (.A0(pcpi_rs1[22]),
    .A1(pcpi_rs1[23]),
    .S(mem_la_wdata[0]),
    .X(_00179_));
 sky130_fd_sc_hd__mux2_1 _40627_ (.A0(pcpi_rs1[20]),
    .A1(pcpi_rs1[21]),
    .S(mem_la_wdata[0]),
    .X(_00178_));
 sky130_fd_sc_hd__mux2_1 _40628_ (.A0(_00175_),
    .A1(_00176_),
    .S(mem_la_wdata[1]),
    .X(_00177_));
 sky130_fd_sc_hd__mux2_1 _40629_ (.A0(pcpi_rs1[18]),
    .A1(pcpi_rs1[19]),
    .S(mem_la_wdata[0]),
    .X(_00176_));
 sky130_fd_sc_hd__mux2_1 _40630_ (.A0(pcpi_rs1[16]),
    .A1(pcpi_rs1[17]),
    .S(mem_la_wdata[0]),
    .X(_00175_));
 sky130_fd_sc_hd__mux2_1 _40631_ (.A0(_00169_),
    .A1(_00172_),
    .S(mem_la_wdata[2]),
    .X(_00173_));
 sky130_fd_sc_hd__mux2_1 _40632_ (.A0(_00170_),
    .A1(_00171_),
    .S(mem_la_wdata[1]),
    .X(_00172_));
 sky130_fd_sc_hd__mux2_1 _40633_ (.A0(pcpi_rs1[14]),
    .A1(pcpi_rs1[15]),
    .S(mem_la_wdata[0]),
    .X(_00171_));
 sky130_fd_sc_hd__mux2_1 _40634_ (.A0(pcpi_rs1[12]),
    .A1(pcpi_rs1[13]),
    .S(mem_la_wdata[0]),
    .X(_00170_));
 sky130_fd_sc_hd__mux2_1 _40635_ (.A0(_00167_),
    .A1(_00168_),
    .S(mem_la_wdata[1]),
    .X(_00169_));
 sky130_fd_sc_hd__mux2_1 _40636_ (.A0(pcpi_rs1[10]),
    .A1(pcpi_rs1[11]),
    .S(mem_la_wdata[0]),
    .X(_00168_));
 sky130_fd_sc_hd__mux2_1 _40637_ (.A0(pcpi_rs1[8]),
    .A1(pcpi_rs1[9]),
    .S(mem_la_wdata[0]),
    .X(_00167_));
 sky130_fd_sc_hd__mux2_1 _40638_ (.A0(_00163_),
    .A1(_00164_),
    .S(mem_la_wdata[1]),
    .X(_00165_));
 sky130_fd_sc_hd__mux2_1 _40639_ (.A0(pcpi_rs1[6]),
    .A1(pcpi_rs1[7]),
    .S(mem_la_wdata[0]),
    .X(_00164_));
 sky130_fd_sc_hd__mux2_1 _40640_ (.A0(pcpi_rs1[4]),
    .A1(pcpi_rs1[5]),
    .S(mem_la_wdata[0]),
    .X(_00163_));
 sky130_fd_sc_hd__mux2_1 _40641_ (.A0(pcpi_rs1[2]),
    .A1(pcpi_rs1[3]),
    .S(mem_la_wdata[0]),
    .X(_00161_));
 sky130_fd_sc_hd__mux2_1 _40642_ (.A0(pcpi_rs1[29]),
    .A1(pcpi_rs1[28]),
    .S(mem_la_wdata[0]),
    .X(_00148_));
 sky130_fd_sc_hd__mux2_1 _40643_ (.A0(pcpi_rs1[28]),
    .A1(pcpi_rs1[27]),
    .S(mem_la_wdata[0]),
    .X(_00144_));
 sky130_fd_sc_hd__mux2_1 _40644_ (.A0(_00140_),
    .A1(_00132_),
    .S(mem_la_wdata[1]),
    .X(_00141_));
 sky130_fd_sc_hd__mux2_1 _40645_ (.A0(pcpi_rs1[27]),
    .A1(pcpi_rs1[26]),
    .S(mem_la_wdata[0]),
    .X(_00140_));
 sky130_fd_sc_hd__mux2_1 _40646_ (.A0(_00136_),
    .A1(_00128_),
    .S(mem_la_wdata[1]),
    .X(_00137_));
 sky130_fd_sc_hd__mux2_1 _40647_ (.A0(pcpi_rs1[26]),
    .A1(pcpi_rs1[25]),
    .S(mem_la_wdata[0]),
    .X(_00136_));
 sky130_fd_sc_hd__mux2_1 _40648_ (.A0(_00132_),
    .A1(_00123_),
    .S(mem_la_wdata[1]),
    .X(_00133_));
 sky130_fd_sc_hd__mux2_1 _40649_ (.A0(pcpi_rs1[25]),
    .A1(pcpi_rs1[24]),
    .S(mem_la_wdata[0]),
    .X(_00132_));
 sky130_fd_sc_hd__mux2_1 _40650_ (.A0(_00128_),
    .A1(_00117_),
    .S(mem_la_wdata[1]),
    .X(_00129_));
 sky130_fd_sc_hd__mux2_1 _40651_ (.A0(pcpi_rs1[24]),
    .A1(pcpi_rs1[23]),
    .S(mem_la_wdata[0]),
    .X(_00128_));
 sky130_fd_sc_hd__mux2_1 _40652_ (.A0(_00098_),
    .A1(_00100_),
    .S(mem_la_wdata[2]),
    .X(_00126_));
 sky130_fd_sc_hd__mux2_1 _40653_ (.A0(_00124_),
    .A1(_00097_),
    .S(mem_la_wdata[2]),
    .X(_00125_));
 sky130_fd_sc_hd__mux2_1 _40654_ (.A0(_00123_),
    .A1(_00111_),
    .S(mem_la_wdata[1]),
    .X(_00124_));
 sky130_fd_sc_hd__mux2_1 _40655_ (.A0(pcpi_rs1[23]),
    .A1(pcpi_rs1[22]),
    .S(mem_la_wdata[0]),
    .X(_00123_));
 sky130_fd_sc_hd__mux2_1 _40656_ (.A0(_00101_),
    .A1(_00094_),
    .S(mem_la_wdata[2]),
    .X(_00122_));
 sky130_fd_sc_hd__mux2_1 _40657_ (.A0(_00088_),
    .A1(_00090_),
    .S(mem_la_wdata[2]),
    .X(_00120_));
 sky130_fd_sc_hd__mux2_1 _40658_ (.A0(_00118_),
    .A1(_00087_),
    .S(mem_la_wdata[2]),
    .X(_00119_));
 sky130_fd_sc_hd__mux2_1 _40659_ (.A0(_00117_),
    .A1(_00105_),
    .S(mem_la_wdata[1]),
    .X(_00118_));
 sky130_fd_sc_hd__mux2_1 _40660_ (.A0(pcpi_rs1[22]),
    .A1(pcpi_rs1[21]),
    .S(mem_la_wdata[0]),
    .X(_00117_));
 sky130_fd_sc_hd__mux2_1 _40661_ (.A0(_00091_),
    .A1(_00084_),
    .S(mem_la_wdata[2]),
    .X(_00116_));
 sky130_fd_sc_hd__mux2_1 _40662_ (.A0(_00074_),
    .A1(_00078_),
    .S(mem_la_wdata[2]),
    .X(_00114_));
 sky130_fd_sc_hd__mux2_1 _40663_ (.A0(_00112_),
    .A1(_00071_),
    .S(mem_la_wdata[2]),
    .X(_00113_));
 sky130_fd_sc_hd__mux2_1 _40664_ (.A0(_00111_),
    .A1(_00096_),
    .S(mem_la_wdata[1]),
    .X(_00112_));
 sky130_fd_sc_hd__mux2_1 _40665_ (.A0(pcpi_rs1[21]),
    .A1(pcpi_rs1[20]),
    .S(mem_la_wdata[0]),
    .X(_00111_));
 sky130_fd_sc_hd__mux2_1 _40666_ (.A0(_00081_),
    .A1(_00067_),
    .S(mem_la_wdata[2]),
    .X(_00110_));
 sky130_fd_sc_hd__mux2_1 _40667_ (.A0(_00056_),
    .A1(_00060_),
    .S(mem_la_wdata[2]),
    .X(_00108_));
 sky130_fd_sc_hd__mux2_1 _40668_ (.A0(_00106_),
    .A1(_00053_),
    .S(mem_la_wdata[2]),
    .X(_00107_));
 sky130_fd_sc_hd__mux2_1 _40669_ (.A0(_00105_),
    .A1(_00086_),
    .S(mem_la_wdata[1]),
    .X(_00106_));
 sky130_fd_sc_hd__mux2_1 _40670_ (.A0(pcpi_rs1[20]),
    .A1(pcpi_rs1[19]),
    .S(mem_la_wdata[0]),
    .X(_00105_));
 sky130_fd_sc_hd__mux2_1 _40671_ (.A0(_00063_),
    .A1(_00049_),
    .S(mem_la_wdata[2]),
    .X(_00104_));
 sky130_fd_sc_hd__mux2_1 _40672_ (.A0(_00100_),
    .A1(_00101_),
    .S(mem_la_wdata[2]),
    .X(_00102_));
 sky130_fd_sc_hd__mux2_1 _40673_ (.A0(_00077_),
    .A1(_00079_),
    .S(mem_la_wdata[1]),
    .X(_00101_));
 sky130_fd_sc_hd__mux2_1 _40674_ (.A0(_00073_),
    .A1(_00076_),
    .S(mem_la_wdata[1]),
    .X(_00100_));
 sky130_fd_sc_hd__mux2_1 _40675_ (.A0(_00097_),
    .A1(_00098_),
    .S(mem_la_wdata[2]),
    .X(_00099_));
 sky130_fd_sc_hd__mux2_1 _40676_ (.A0(_00070_),
    .A1(_00072_),
    .S(mem_la_wdata[1]),
    .X(_00098_));
 sky130_fd_sc_hd__mux2_1 _40677_ (.A0(_00096_),
    .A1(_00069_),
    .S(mem_la_wdata[1]),
    .X(_00097_));
 sky130_fd_sc_hd__mux2_1 _40678_ (.A0(pcpi_rs1[19]),
    .A1(pcpi_rs1[18]),
    .S(mem_la_wdata[0]),
    .X(_00096_));
 sky130_fd_sc_hd__mux2_1 _40679_ (.A0(_00080_),
    .A1(_00066_),
    .S(mem_la_wdata[1]),
    .X(_00094_));
 sky130_fd_sc_hd__mux2_1 _40680_ (.A0(_00090_),
    .A1(_00091_),
    .S(mem_la_wdata[2]),
    .X(_00092_));
 sky130_fd_sc_hd__mux2_1 _40681_ (.A0(_00059_),
    .A1(_00061_),
    .S(mem_la_wdata[1]),
    .X(_00091_));
 sky130_fd_sc_hd__mux2_1 _40682_ (.A0(_00055_),
    .A1(_00058_),
    .S(mem_la_wdata[1]),
    .X(_00090_));
 sky130_fd_sc_hd__mux2_1 _40683_ (.A0(_00087_),
    .A1(_00088_),
    .S(mem_la_wdata[2]),
    .X(_00089_));
 sky130_fd_sc_hd__mux2_1 _40684_ (.A0(_00052_),
    .A1(_00054_),
    .S(mem_la_wdata[1]),
    .X(_00088_));
 sky130_fd_sc_hd__mux2_1 _40685_ (.A0(_00086_),
    .A1(_00051_),
    .S(mem_la_wdata[1]),
    .X(_00087_));
 sky130_fd_sc_hd__mux2_1 _40686_ (.A0(pcpi_rs1[18]),
    .A1(pcpi_rs1[17]),
    .S(mem_la_wdata[0]),
    .X(_00086_));
 sky130_fd_sc_hd__mux2_1 _40687_ (.A0(_00062_),
    .A1(_00048_),
    .S(mem_la_wdata[1]),
    .X(_00084_));
 sky130_fd_sc_hd__mux2_1 _40688_ (.A0(_00078_),
    .A1(_00081_),
    .S(mem_la_wdata[2]),
    .X(_00082_));
 sky130_fd_sc_hd__mux2_1 _40689_ (.A0(_00079_),
    .A1(_00080_),
    .S(mem_la_wdata[1]),
    .X(_00081_));
 sky130_fd_sc_hd__mux2_1 _40690_ (.A0(pcpi_rs1[3]),
    .A1(pcpi_rs1[2]),
    .S(mem_la_wdata[0]),
    .X(_00080_));
 sky130_fd_sc_hd__mux2_1 _40691_ (.A0(pcpi_rs1[5]),
    .A1(pcpi_rs1[4]),
    .S(mem_la_wdata[0]),
    .X(_00079_));
 sky130_fd_sc_hd__mux2_1 _40692_ (.A0(_00076_),
    .A1(_00077_),
    .S(mem_la_wdata[1]),
    .X(_00078_));
 sky130_fd_sc_hd__mux2_1 _40693_ (.A0(pcpi_rs1[7]),
    .A1(pcpi_rs1[6]),
    .S(mem_la_wdata[0]),
    .X(_00077_));
 sky130_fd_sc_hd__mux2_1 _40694_ (.A0(pcpi_rs1[9]),
    .A1(pcpi_rs1[8]),
    .S(mem_la_wdata[0]),
    .X(_00076_));
 sky130_fd_sc_hd__mux2_1 _40695_ (.A0(_00071_),
    .A1(_00074_),
    .S(mem_la_wdata[2]),
    .X(_00075_));
 sky130_fd_sc_hd__mux2_1 _40696_ (.A0(_00072_),
    .A1(_00073_),
    .S(mem_la_wdata[1]),
    .X(_00074_));
 sky130_fd_sc_hd__mux2_1 _40697_ (.A0(pcpi_rs1[11]),
    .A1(pcpi_rs1[10]),
    .S(mem_la_wdata[0]),
    .X(_00073_));
 sky130_fd_sc_hd__mux2_1 _40698_ (.A0(pcpi_rs1[13]),
    .A1(pcpi_rs1[12]),
    .S(mem_la_wdata[0]),
    .X(_00072_));
 sky130_fd_sc_hd__mux2_1 _40699_ (.A0(_00069_),
    .A1(_00070_),
    .S(mem_la_wdata[1]),
    .X(_00071_));
 sky130_fd_sc_hd__mux2_1 _40700_ (.A0(pcpi_rs1[15]),
    .A1(pcpi_rs1[14]),
    .S(mem_la_wdata[0]),
    .X(_00070_));
 sky130_fd_sc_hd__mux2_1 _40701_ (.A0(pcpi_rs1[17]),
    .A1(pcpi_rs1[16]),
    .S(mem_la_wdata[0]),
    .X(_00069_));
 sky130_fd_sc_hd__mux2_1 _40702_ (.A0(pcpi_rs1[1]),
    .A1(pcpi_rs1[0]),
    .S(mem_la_wdata[0]),
    .X(_00066_));
 sky130_fd_sc_hd__mux2_1 _40703_ (.A0(_00060_),
    .A1(_00063_),
    .S(mem_la_wdata[2]),
    .X(_00064_));
 sky130_fd_sc_hd__mux2_1 _40704_ (.A0(_00061_),
    .A1(_00062_),
    .S(mem_la_wdata[1]),
    .X(_00063_));
 sky130_fd_sc_hd__mux2_1 _40705_ (.A0(pcpi_rs1[2]),
    .A1(pcpi_rs1[1]),
    .S(mem_la_wdata[0]),
    .X(_00062_));
 sky130_fd_sc_hd__mux2_1 _40706_ (.A0(pcpi_rs1[4]),
    .A1(pcpi_rs1[3]),
    .S(mem_la_wdata[0]),
    .X(_00061_));
 sky130_fd_sc_hd__mux2_1 _40707_ (.A0(_00058_),
    .A1(_00059_),
    .S(mem_la_wdata[1]),
    .X(_00060_));
 sky130_fd_sc_hd__mux2_1 _40708_ (.A0(pcpi_rs1[6]),
    .A1(pcpi_rs1[5]),
    .S(mem_la_wdata[0]),
    .X(_00059_));
 sky130_fd_sc_hd__mux2_1 _40709_ (.A0(pcpi_rs1[8]),
    .A1(pcpi_rs1[7]),
    .S(mem_la_wdata[0]),
    .X(_00058_));
 sky130_fd_sc_hd__mux2_1 _40710_ (.A0(_00053_),
    .A1(_00056_),
    .S(mem_la_wdata[2]),
    .X(_00057_));
 sky130_fd_sc_hd__mux2_1 _40711_ (.A0(_00054_),
    .A1(_00055_),
    .S(mem_la_wdata[1]),
    .X(_00056_));
 sky130_fd_sc_hd__mux2_1 _40712_ (.A0(pcpi_rs1[10]),
    .A1(pcpi_rs1[9]),
    .S(mem_la_wdata[0]),
    .X(_00055_));
 sky130_fd_sc_hd__mux2_1 _40713_ (.A0(pcpi_rs1[12]),
    .A1(pcpi_rs1[11]),
    .S(mem_la_wdata[0]),
    .X(_00054_));
 sky130_fd_sc_hd__mux2_1 _40714_ (.A0(_00051_),
    .A1(_00052_),
    .S(mem_la_wdata[1]),
    .X(_00053_));
 sky130_fd_sc_hd__mux2_1 _40715_ (.A0(pcpi_rs1[14]),
    .A1(pcpi_rs1[13]),
    .S(mem_la_wdata[0]),
    .X(_00052_));
 sky130_fd_sc_hd__mux2_1 _40716_ (.A0(pcpi_rs1[16]),
    .A1(pcpi_rs1[15]),
    .S(mem_la_wdata[0]),
    .X(_00051_));
 sky130_fd_sc_hd__mux2_1 _40717_ (.A0(_02408_),
    .A1(pcpi_rs2[31]),
    .S(instr_sub),
    .X(_02409_));
 sky130_fd_sc_hd__mux2_1 _40718_ (.A0(_02406_),
    .A1(_02405_),
    .S(instr_sub),
    .X(_02407_));
 sky130_fd_sc_hd__mux2_1 _40719_ (.A0(_02403_),
    .A1(_02402_),
    .S(instr_sub),
    .X(_02404_));
 sky130_fd_sc_hd__mux2_1 _40720_ (.A0(_02400_),
    .A1(_02399_),
    .S(instr_sub),
    .X(_02401_));
 sky130_fd_sc_hd__mux2_1 _40721_ (.A0(_02397_),
    .A1(_02396_),
    .S(instr_sub),
    .X(_02398_));
 sky130_fd_sc_hd__mux2_1 _40722_ (.A0(_02394_),
    .A1(_02393_),
    .S(instr_sub),
    .X(_02395_));
 sky130_fd_sc_hd__mux2_1 _40723_ (.A0(_02391_),
    .A1(_02390_),
    .S(instr_sub),
    .X(_02392_));
 sky130_fd_sc_hd__mux2_1 _40724_ (.A0(_02388_),
    .A1(_02387_),
    .S(instr_sub),
    .X(_02389_));
 sky130_fd_sc_hd__mux2_1 _40725_ (.A0(_02385_),
    .A1(_02384_),
    .S(instr_sub),
    .X(_02386_));
 sky130_fd_sc_hd__mux2_1 _40726_ (.A0(_02382_),
    .A1(_02381_),
    .S(instr_sub),
    .X(_02383_));
 sky130_fd_sc_hd__mux2_1 _40727_ (.A0(_02379_),
    .A1(_02378_),
    .S(instr_sub),
    .X(_02380_));
 sky130_fd_sc_hd__mux2_1 _40728_ (.A0(_02376_),
    .A1(_02375_),
    .S(instr_sub),
    .X(_02377_));
 sky130_fd_sc_hd__mux2_1 _40729_ (.A0(_02373_),
    .A1(_02372_),
    .S(instr_sub),
    .X(_02374_));
 sky130_fd_sc_hd__mux2_1 _40730_ (.A0(_02370_),
    .A1(_02369_),
    .S(instr_sub),
    .X(_02371_));
 sky130_fd_sc_hd__mux2_1 _40731_ (.A0(_02367_),
    .A1(_02366_),
    .S(instr_sub),
    .X(_02368_));
 sky130_fd_sc_hd__mux2_1 _40732_ (.A0(_02364_),
    .A1(_02363_),
    .S(instr_sub),
    .X(_02365_));
 sky130_fd_sc_hd__mux2_1 _40733_ (.A0(_02361_),
    .A1(_02360_),
    .S(instr_sub),
    .X(_02362_));
 sky130_fd_sc_hd__mux2_1 _40734_ (.A0(_02358_),
    .A1(_02357_),
    .S(instr_sub),
    .X(_02359_));
 sky130_fd_sc_hd__mux2_1 _40735_ (.A0(_02355_),
    .A1(_02354_),
    .S(instr_sub),
    .X(_02356_));
 sky130_fd_sc_hd__mux2_1 _40736_ (.A0(_02352_),
    .A1(_02351_),
    .S(instr_sub),
    .X(_02353_));
 sky130_fd_sc_hd__mux2_1 _40737_ (.A0(_02349_),
    .A1(_02348_),
    .S(instr_sub),
    .X(_02350_));
 sky130_fd_sc_hd__mux2_1 _40738_ (.A0(_02346_),
    .A1(_02345_),
    .S(instr_sub),
    .X(_02347_));
 sky130_fd_sc_hd__mux2_1 _40739_ (.A0(_02343_),
    .A1(_02342_),
    .S(instr_sub),
    .X(_02344_));
 sky130_fd_sc_hd__mux2_1 _40740_ (.A0(_02340_),
    .A1(_02339_),
    .S(instr_sub),
    .X(_02341_));
 sky130_fd_sc_hd__mux2_1 _40741_ (.A0(_02337_),
    .A1(_02336_),
    .S(instr_sub),
    .X(_02338_));
 sky130_fd_sc_hd__mux2_1 _40742_ (.A0(_02334_),
    .A1(_02333_),
    .S(instr_sub),
    .X(_02335_));
 sky130_fd_sc_hd__mux2_1 _40743_ (.A0(_02331_),
    .A1(_02330_),
    .S(instr_sub),
    .X(_02332_));
 sky130_fd_sc_hd__mux2_1 _40744_ (.A0(_02328_),
    .A1(_02327_),
    .S(instr_sub),
    .X(_02329_));
 sky130_fd_sc_hd__mux2_1 _40745_ (.A0(_02325_),
    .A1(_02324_),
    .S(instr_sub),
    .X(_02326_));
 sky130_fd_sc_hd__mux2_1 _40746_ (.A0(_02322_),
    .A1(_02321_),
    .S(instr_sub),
    .X(_02323_));
 sky130_fd_sc_hd__mux2_1 _40747_ (.A0(_02319_),
    .A1(_02318_),
    .S(instr_sub),
    .X(_02320_));
 sky130_fd_sc_hd__mux2_1 _40748_ (.A0(_02313_),
    .A1(_02314_),
    .S(_00306_),
    .X(_02315_));
 sky130_fd_sc_hd__mux2_1 _40749_ (.A0(_02311_),
    .A1(_02315_),
    .S(_00303_),
    .X(_02316_));
 sky130_fd_sc_hd__mux2_1 _40750_ (.A0(_02311_),
    .A1(_02312_),
    .S(_00305_),
    .X(_02313_));
 sky130_fd_sc_hd__mux2_1 _40751_ (.A0(_02307_),
    .A1(_02308_),
    .S(\irq_state[1] ),
    .X(_02309_));
 sky130_fd_sc_hd__mux2_1 _40752_ (.A0(_02309_),
    .A1(_02307_),
    .S(_02217_),
    .X(_02310_));
 sky130_fd_sc_hd__mux2_1 _40753_ (.A0(_02302_),
    .A1(\irq_pending[0] ),
    .S(_01208_),
    .X(_02303_));
 sky130_fd_sc_hd__mux2_1 _40754_ (.A0(\reg_out[0] ),
    .A1(\alu_out_q[0] ),
    .S(latched_stalu),
    .X(_02070_));
 sky130_fd_sc_hd__mux2_1 _40755_ (.A0(_02063_),
    .A1(_00343_),
    .S(is_beq_bne_blt_bge_bltu_bgeu),
    .X(_02064_));
 sky130_fd_sc_hd__mux2_1 _40756_ (.A0(_02056_),
    .A1(_02055_),
    .S(_01714_),
    .X(_02057_));
 sky130_fd_sc_hd__mux2_1 _40757_ (.A0(_02058_),
    .A1(_02057_),
    .S(_01717_),
    .X(_02059_));
 sky130_fd_sc_hd__mux2_1 _40758_ (.A0(\pcpi_mul.rd[31] ),
    .A1(\pcpi_mul.rd[63] ),
    .S(\pcpi_mul.shift_out ),
    .X(_02054_));
 sky130_fd_sc_hd__mux2_1 _40759_ (.A0(_01908_),
    .A1(_02052_),
    .S(_01816_),
    .X(_02053_));
 sky130_fd_sc_hd__mux2_1 _40760_ (.A0(_02047_),
    .A1(_02046_),
    .S(_01714_),
    .X(_02048_));
 sky130_fd_sc_hd__mux2_1 _40761_ (.A0(_02049_),
    .A1(_02048_),
    .S(_01717_),
    .X(_02050_));
 sky130_fd_sc_hd__mux2_1 _40762_ (.A0(\pcpi_mul.rd[30] ),
    .A1(\pcpi_mul.rd[62] ),
    .S(\pcpi_mul.shift_out ),
    .X(_02045_));
 sky130_fd_sc_hd__mux2_1 _40763_ (.A0(_01908_),
    .A1(_02043_),
    .S(_01816_),
    .X(_02044_));
 sky130_fd_sc_hd__mux2_1 _40764_ (.A0(_02038_),
    .A1(_02037_),
    .S(_01714_),
    .X(_02039_));
 sky130_fd_sc_hd__mux2_1 _40765_ (.A0(_02040_),
    .A1(_02039_),
    .S(_01717_),
    .X(_02041_));
 sky130_fd_sc_hd__mux2_1 _40766_ (.A0(\pcpi_mul.rd[29] ),
    .A1(\pcpi_mul.rd[61] ),
    .S(\pcpi_mul.shift_out ),
    .X(_02036_));
 sky130_fd_sc_hd__mux2_1 _40767_ (.A0(_01908_),
    .A1(_02034_),
    .S(_01816_),
    .X(_02035_));
 sky130_fd_sc_hd__mux2_1 _40768_ (.A0(_02029_),
    .A1(_02028_),
    .S(_01714_),
    .X(_02030_));
 sky130_fd_sc_hd__mux2_1 _40769_ (.A0(_02031_),
    .A1(_02030_),
    .S(_01717_),
    .X(_02032_));
 sky130_fd_sc_hd__mux2_1 _40770_ (.A0(\pcpi_mul.rd[28] ),
    .A1(\pcpi_mul.rd[60] ),
    .S(\pcpi_mul.shift_out ),
    .X(_02027_));
 sky130_fd_sc_hd__mux2_1 _40771_ (.A0(_01908_),
    .A1(_02025_),
    .S(_01816_),
    .X(_02026_));
 sky130_fd_sc_hd__mux2_1 _40772_ (.A0(_02020_),
    .A1(_02019_),
    .S(_01714_),
    .X(_02021_));
 sky130_fd_sc_hd__mux2_1 _40773_ (.A0(_02022_),
    .A1(_02021_),
    .S(_01717_),
    .X(_02023_));
 sky130_fd_sc_hd__mux2_1 _40774_ (.A0(\pcpi_mul.rd[27] ),
    .A1(\pcpi_mul.rd[59] ),
    .S(\pcpi_mul.shift_out ),
    .X(_02018_));
 sky130_fd_sc_hd__mux2_1 _40775_ (.A0(_01908_),
    .A1(_02016_),
    .S(_01816_),
    .X(_02017_));
 sky130_fd_sc_hd__mux2_1 _40776_ (.A0(_02011_),
    .A1(_02010_),
    .S(_01714_),
    .X(_02012_));
 sky130_fd_sc_hd__mux2_1 _40777_ (.A0(_02013_),
    .A1(_02012_),
    .S(_01717_),
    .X(_02014_));
 sky130_fd_sc_hd__mux2_1 _40778_ (.A0(\pcpi_mul.rd[26] ),
    .A1(\pcpi_mul.rd[58] ),
    .S(\pcpi_mul.shift_out ),
    .X(_02009_));
 sky130_fd_sc_hd__mux2_1 _40779_ (.A0(_01908_),
    .A1(_02007_),
    .S(_01816_),
    .X(_02008_));
 sky130_fd_sc_hd__mux2_1 _40780_ (.A0(_02002_),
    .A1(_02001_),
    .S(_01714_),
    .X(_02003_));
 sky130_fd_sc_hd__mux2_1 _40781_ (.A0(_02004_),
    .A1(_02003_),
    .S(_01717_),
    .X(_02005_));
 sky130_fd_sc_hd__mux2_1 _40782_ (.A0(\pcpi_mul.rd[25] ),
    .A1(\pcpi_mul.rd[57] ),
    .S(\pcpi_mul.shift_out ),
    .X(_02000_));
 sky130_fd_sc_hd__mux2_1 _40783_ (.A0(_01908_),
    .A1(_01998_),
    .S(_01816_),
    .X(_01999_));
 sky130_fd_sc_hd__mux2_1 _40784_ (.A0(_01993_),
    .A1(_01992_),
    .S(_01714_),
    .X(_01994_));
 sky130_fd_sc_hd__mux2_1 _40785_ (.A0(_01995_),
    .A1(_01994_),
    .S(_01717_),
    .X(_01996_));
 sky130_fd_sc_hd__mux2_1 _40786_ (.A0(\pcpi_mul.rd[24] ),
    .A1(\pcpi_mul.rd[56] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01991_));
 sky130_fd_sc_hd__mux2_1 _40787_ (.A0(_01908_),
    .A1(_01989_),
    .S(_01816_),
    .X(_01990_));
 sky130_fd_sc_hd__mux2_1 _40788_ (.A0(_01984_),
    .A1(_01983_),
    .S(_01714_),
    .X(_01985_));
 sky130_fd_sc_hd__mux2_1 _40789_ (.A0(_01986_),
    .A1(_01985_),
    .S(_01717_),
    .X(_01987_));
 sky130_fd_sc_hd__mux2_1 _40790_ (.A0(\pcpi_mul.rd[23] ),
    .A1(\pcpi_mul.rd[55] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01982_));
 sky130_fd_sc_hd__mux2_1 _40791_ (.A0(_01908_),
    .A1(_01980_),
    .S(_01816_),
    .X(_01981_));
 sky130_fd_sc_hd__mux2_1 _40792_ (.A0(_01975_),
    .A1(_01974_),
    .S(_01714_),
    .X(_01976_));
 sky130_fd_sc_hd__mux2_1 _40793_ (.A0(_01977_),
    .A1(_01976_),
    .S(_01717_),
    .X(_01978_));
 sky130_fd_sc_hd__mux2_1 _40794_ (.A0(\pcpi_mul.rd[22] ),
    .A1(\pcpi_mul.rd[54] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01973_));
 sky130_fd_sc_hd__mux2_1 _40795_ (.A0(_01908_),
    .A1(_01971_),
    .S(_01816_),
    .X(_01972_));
 sky130_fd_sc_hd__mux2_1 _40796_ (.A0(_01966_),
    .A1(_01965_),
    .S(_01714_),
    .X(_01967_));
 sky130_fd_sc_hd__mux2_1 _40797_ (.A0(_01968_),
    .A1(_01967_),
    .S(_01717_),
    .X(_01969_));
 sky130_fd_sc_hd__mux2_1 _40798_ (.A0(\pcpi_mul.rd[21] ),
    .A1(\pcpi_mul.rd[53] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01964_));
 sky130_fd_sc_hd__mux2_1 _40799_ (.A0(_01908_),
    .A1(_01962_),
    .S(_01816_),
    .X(_01963_));
 sky130_fd_sc_hd__mux2_1 _40800_ (.A0(_01957_),
    .A1(_01956_),
    .S(_01714_),
    .X(_01958_));
 sky130_fd_sc_hd__mux2_1 _40801_ (.A0(_01959_),
    .A1(_01958_),
    .S(_01717_),
    .X(_01960_));
 sky130_fd_sc_hd__mux2_1 _40802_ (.A0(\pcpi_mul.rd[20] ),
    .A1(\pcpi_mul.rd[52] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01955_));
 sky130_fd_sc_hd__mux2_1 _40803_ (.A0(_01908_),
    .A1(_01953_),
    .S(_01816_),
    .X(_01954_));
 sky130_fd_sc_hd__mux2_1 _40804_ (.A0(_01948_),
    .A1(_01947_),
    .S(_01714_),
    .X(_01949_));
 sky130_fd_sc_hd__mux2_1 _40805_ (.A0(_01950_),
    .A1(_01949_),
    .S(_01717_),
    .X(_01951_));
 sky130_fd_sc_hd__mux2_1 _40806_ (.A0(\pcpi_mul.rd[19] ),
    .A1(\pcpi_mul.rd[51] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01946_));
 sky130_fd_sc_hd__mux2_1 _40807_ (.A0(_01908_),
    .A1(_01944_),
    .S(_01816_),
    .X(_01945_));
 sky130_fd_sc_hd__mux2_1 _40808_ (.A0(_01939_),
    .A1(_01938_),
    .S(_01714_),
    .X(_01940_));
 sky130_fd_sc_hd__mux2_1 _40809_ (.A0(_01941_),
    .A1(_01940_),
    .S(_01717_),
    .X(_01942_));
 sky130_fd_sc_hd__mux2_1 _40810_ (.A0(\pcpi_mul.rd[18] ),
    .A1(\pcpi_mul.rd[50] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01937_));
 sky130_fd_sc_hd__mux2_1 _40811_ (.A0(_01908_),
    .A1(_01935_),
    .S(_01816_),
    .X(_01936_));
 sky130_fd_sc_hd__mux2_1 _40812_ (.A0(_01930_),
    .A1(_01929_),
    .S(_01714_),
    .X(_01931_));
 sky130_fd_sc_hd__mux2_1 _40813_ (.A0(_01932_),
    .A1(_01931_),
    .S(_01717_),
    .X(_01933_));
 sky130_fd_sc_hd__mux2_1 _40814_ (.A0(\pcpi_mul.rd[17] ),
    .A1(\pcpi_mul.rd[49] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01928_));
 sky130_fd_sc_hd__mux2_1 _40815_ (.A0(_01908_),
    .A1(_01926_),
    .S(_01816_),
    .X(_01927_));
 sky130_fd_sc_hd__mux2_1 _40816_ (.A0(_01921_),
    .A1(_01920_),
    .S(_01714_),
    .X(_01922_));
 sky130_fd_sc_hd__mux2_1 _40817_ (.A0(_01923_),
    .A1(_01922_),
    .S(_01717_),
    .X(_01924_));
 sky130_fd_sc_hd__mux2_1 _40818_ (.A0(\pcpi_mul.rd[16] ),
    .A1(\pcpi_mul.rd[48] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01919_));
 sky130_fd_sc_hd__mux2_1 _40819_ (.A0(_01908_),
    .A1(_01917_),
    .S(_01816_),
    .X(_01918_));
 sky130_fd_sc_hd__mux2_1 _40820_ (.A0(_01912_),
    .A1(_01911_),
    .S(_01714_),
    .X(_01913_));
 sky130_fd_sc_hd__mux2_1 _40821_ (.A0(_01914_),
    .A1(_01913_),
    .S(_01717_),
    .X(_01915_));
 sky130_fd_sc_hd__mux2_1 _40822_ (.A0(\pcpi_mul.rd[15] ),
    .A1(\pcpi_mul.rd[47] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01910_));
 sky130_fd_sc_hd__mux2_1 _40823_ (.A0(_01908_),
    .A1(_01907_),
    .S(_01816_),
    .X(_01909_));
 sky130_fd_sc_hd__mux2_1 _40824_ (.A0(_01906_),
    .A1(_01904_),
    .S(_01683_),
    .X(_01907_));
 sky130_fd_sc_hd__mux2_1 _40825_ (.A0(mem_rdata[15]),
    .A1(mem_rdata[31]),
    .S(pcpi_rs1[1]),
    .X(_01905_));
 sky130_fd_sc_hd__mux2_1 _40826_ (.A0(_01899_),
    .A1(_01898_),
    .S(_01714_),
    .X(_01900_));
 sky130_fd_sc_hd__mux2_1 _40827_ (.A0(_01901_),
    .A1(_01900_),
    .S(_01717_),
    .X(_01902_));
 sky130_fd_sc_hd__mux2_1 _40828_ (.A0(\pcpi_mul.rd[14] ),
    .A1(\pcpi_mul.rd[46] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01897_));
 sky130_fd_sc_hd__mux2_1 _40829_ (.A0(_01895_),
    .A1(_01894_),
    .S(_01816_),
    .X(_01896_));
 sky130_fd_sc_hd__mux2_1 _40830_ (.A0(_01893_),
    .A1(_01891_),
    .S(_01683_),
    .X(_01894_));
 sky130_fd_sc_hd__mux2_1 _40831_ (.A0(mem_rdata[14]),
    .A1(mem_rdata[30]),
    .S(pcpi_rs1[1]),
    .X(_01892_));
 sky130_fd_sc_hd__mux2_1 _40832_ (.A0(_01886_),
    .A1(_01885_),
    .S(_01714_),
    .X(_01887_));
 sky130_fd_sc_hd__mux2_1 _40833_ (.A0(_01888_),
    .A1(_01887_),
    .S(_01717_),
    .X(_01889_));
 sky130_fd_sc_hd__mux2_1 _40834_ (.A0(\pcpi_mul.rd[13] ),
    .A1(\pcpi_mul.rd[45] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01884_));
 sky130_fd_sc_hd__mux2_1 _40835_ (.A0(_01882_),
    .A1(_01881_),
    .S(_01816_),
    .X(_01883_));
 sky130_fd_sc_hd__mux2_1 _40836_ (.A0(_01880_),
    .A1(_01878_),
    .S(_01683_),
    .X(_01881_));
 sky130_fd_sc_hd__mux2_1 _40837_ (.A0(mem_rdata[13]),
    .A1(mem_rdata[29]),
    .S(pcpi_rs1[1]),
    .X(_01879_));
 sky130_fd_sc_hd__mux2_1 _40838_ (.A0(_01873_),
    .A1(_01872_),
    .S(_01714_),
    .X(_01874_));
 sky130_fd_sc_hd__mux2_1 _40839_ (.A0(_01875_),
    .A1(_01874_),
    .S(_01717_),
    .X(_01876_));
 sky130_fd_sc_hd__mux2_1 _40840_ (.A0(\pcpi_mul.rd[12] ),
    .A1(\pcpi_mul.rd[44] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01871_));
 sky130_fd_sc_hd__mux2_1 _40841_ (.A0(_01869_),
    .A1(_01868_),
    .S(_01816_),
    .X(_01870_));
 sky130_fd_sc_hd__mux2_1 _40842_ (.A0(_01867_),
    .A1(_01865_),
    .S(_01683_),
    .X(_01868_));
 sky130_fd_sc_hd__mux2_1 _40843_ (.A0(mem_rdata[12]),
    .A1(mem_rdata[28]),
    .S(pcpi_rs1[1]),
    .X(_01866_));
 sky130_fd_sc_hd__mux2_1 _40844_ (.A0(_01860_),
    .A1(_01859_),
    .S(_01714_),
    .X(_01861_));
 sky130_fd_sc_hd__mux2_1 _40845_ (.A0(_01862_),
    .A1(_01861_),
    .S(_01717_),
    .X(_01863_));
 sky130_fd_sc_hd__mux2_1 _40846_ (.A0(\pcpi_mul.rd[11] ),
    .A1(\pcpi_mul.rd[43] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01858_));
 sky130_fd_sc_hd__mux2_1 _40847_ (.A0(_01856_),
    .A1(_01855_),
    .S(_01816_),
    .X(_01857_));
 sky130_fd_sc_hd__mux2_1 _40848_ (.A0(_01854_),
    .A1(_01852_),
    .S(_01683_),
    .X(_01855_));
 sky130_fd_sc_hd__mux2_1 _40849_ (.A0(mem_rdata[11]),
    .A1(mem_rdata[27]),
    .S(pcpi_rs1[1]),
    .X(_01853_));
 sky130_fd_sc_hd__mux2_1 _40850_ (.A0(_01847_),
    .A1(_01846_),
    .S(_01714_),
    .X(_01848_));
 sky130_fd_sc_hd__mux2_1 _40851_ (.A0(_01849_),
    .A1(_01848_),
    .S(_01717_),
    .X(_01850_));
 sky130_fd_sc_hd__mux2_1 _40852_ (.A0(\pcpi_mul.rd[10] ),
    .A1(\pcpi_mul.rd[42] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01845_));
 sky130_fd_sc_hd__mux2_1 _40853_ (.A0(_01843_),
    .A1(_01842_),
    .S(_01816_),
    .X(_01844_));
 sky130_fd_sc_hd__mux2_1 _40854_ (.A0(_01841_),
    .A1(_01839_),
    .S(_01683_),
    .X(_01842_));
 sky130_fd_sc_hd__mux2_1 _40855_ (.A0(mem_rdata[10]),
    .A1(mem_rdata[26]),
    .S(pcpi_rs1[1]),
    .X(_01840_));
 sky130_fd_sc_hd__mux2_1 _40856_ (.A0(_01834_),
    .A1(_01833_),
    .S(_01714_),
    .X(_01835_));
 sky130_fd_sc_hd__mux2_1 _40857_ (.A0(_01836_),
    .A1(_01835_),
    .S(_01717_),
    .X(_01837_));
 sky130_fd_sc_hd__mux2_1 _40858_ (.A0(\pcpi_mul.rd[9] ),
    .A1(\pcpi_mul.rd[41] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01832_));
 sky130_fd_sc_hd__mux2_1 _40859_ (.A0(_01830_),
    .A1(_01829_),
    .S(_01816_),
    .X(_01831_));
 sky130_fd_sc_hd__mux2_1 _40860_ (.A0(_01828_),
    .A1(_01826_),
    .S(_01683_),
    .X(_01829_));
 sky130_fd_sc_hd__mux2_1 _40861_ (.A0(mem_rdata[9]),
    .A1(mem_rdata[25]),
    .S(pcpi_rs1[1]),
    .X(_01827_));
 sky130_fd_sc_hd__mux2_1 _40862_ (.A0(_01821_),
    .A1(_01820_),
    .S(_01714_),
    .X(_01822_));
 sky130_fd_sc_hd__mux2_1 _40863_ (.A0(_01823_),
    .A1(_01822_),
    .S(_01717_),
    .X(_01824_));
 sky130_fd_sc_hd__mux2_1 _40864_ (.A0(\pcpi_mul.rd[8] ),
    .A1(\pcpi_mul.rd[40] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01819_));
 sky130_fd_sc_hd__mux2_1 _40865_ (.A0(_01817_),
    .A1(_01815_),
    .S(_01816_),
    .X(_01818_));
 sky130_fd_sc_hd__mux2_1 _40866_ (.A0(_01814_),
    .A1(_01812_),
    .S(_01683_),
    .X(_01815_));
 sky130_fd_sc_hd__mux2_1 _40867_ (.A0(mem_rdata[8]),
    .A1(mem_rdata[24]),
    .S(pcpi_rs1[1]),
    .X(_01813_));
 sky130_fd_sc_hd__mux2_1 _40868_ (.A0(_01807_),
    .A1(_01806_),
    .S(_01714_),
    .X(_01808_));
 sky130_fd_sc_hd__mux2_1 _40869_ (.A0(_01809_),
    .A1(_01808_),
    .S(_01717_),
    .X(_01810_));
 sky130_fd_sc_hd__mux2_1 _40870_ (.A0(\pcpi_mul.rd[7] ),
    .A1(\pcpi_mul.rd[39] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01805_));
 sky130_fd_sc_hd__mux2_1 _40871_ (.A0(_01803_),
    .A1(_01799_),
    .S(_01683_),
    .X(_01804_));
 sky130_fd_sc_hd__mux2_1 _40872_ (.A0(mem_rdata[7]),
    .A1(mem_rdata[23]),
    .S(pcpi_rs1[1]),
    .X(_01802_));
 sky130_fd_sc_hd__mux2_1 _40873_ (.A0(_01800_),
    .A1(_01799_),
    .S(_00304_),
    .X(_01801_));
 sky130_fd_sc_hd__mux2_1 _40874_ (.A0(_01794_),
    .A1(_01793_),
    .S(_01714_),
    .X(_01795_));
 sky130_fd_sc_hd__mux2_1 _40875_ (.A0(_01796_),
    .A1(_01795_),
    .S(_01717_),
    .X(_01797_));
 sky130_fd_sc_hd__mux2_1 _40876_ (.A0(\pcpi_mul.rd[6] ),
    .A1(\pcpi_mul.rd[38] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01792_));
 sky130_fd_sc_hd__mux2_1 _40877_ (.A0(_01790_),
    .A1(_01786_),
    .S(_01683_),
    .X(_01791_));
 sky130_fd_sc_hd__mux2_1 _40878_ (.A0(mem_rdata[6]),
    .A1(mem_rdata[22]),
    .S(pcpi_rs1[1]),
    .X(_01789_));
 sky130_fd_sc_hd__mux2_1 _40879_ (.A0(_01787_),
    .A1(_01786_),
    .S(_00304_),
    .X(_01788_));
 sky130_fd_sc_hd__mux2_1 _40880_ (.A0(_01781_),
    .A1(_01780_),
    .S(_01714_),
    .X(_01782_));
 sky130_fd_sc_hd__mux2_1 _40881_ (.A0(_01783_),
    .A1(_01782_),
    .S(_01717_),
    .X(_01784_));
 sky130_fd_sc_hd__mux2_1 _40882_ (.A0(\pcpi_mul.rd[5] ),
    .A1(\pcpi_mul.rd[37] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01779_));
 sky130_fd_sc_hd__mux2_1 _40883_ (.A0(_01777_),
    .A1(_01773_),
    .S(_01683_),
    .X(_01778_));
 sky130_fd_sc_hd__mux2_1 _40884_ (.A0(mem_rdata[5]),
    .A1(mem_rdata[21]),
    .S(pcpi_rs1[1]),
    .X(_01776_));
 sky130_fd_sc_hd__mux2_1 _40885_ (.A0(_01774_),
    .A1(_01773_),
    .S(_00304_),
    .X(_01775_));
 sky130_fd_sc_hd__mux2_1 _40886_ (.A0(_01768_),
    .A1(_01767_),
    .S(_01714_),
    .X(_01769_));
 sky130_fd_sc_hd__mux2_1 _40887_ (.A0(_01770_),
    .A1(_01769_),
    .S(_01717_),
    .X(_01771_));
 sky130_fd_sc_hd__mux2_1 _40888_ (.A0(\pcpi_mul.rd[4] ),
    .A1(\pcpi_mul.rd[36] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01766_));
 sky130_fd_sc_hd__mux2_1 _40889_ (.A0(_01764_),
    .A1(_01760_),
    .S(_01683_),
    .X(_01765_));
 sky130_fd_sc_hd__mux2_1 _40890_ (.A0(mem_rdata[4]),
    .A1(mem_rdata[20]),
    .S(pcpi_rs1[1]),
    .X(_01763_));
 sky130_fd_sc_hd__mux2_1 _40891_ (.A0(_01761_),
    .A1(_01760_),
    .S(_00304_),
    .X(_01762_));
 sky130_fd_sc_hd__mux2_1 _40892_ (.A0(_01755_),
    .A1(_01754_),
    .S(_01714_),
    .X(_01756_));
 sky130_fd_sc_hd__mux2_1 _40893_ (.A0(_01757_),
    .A1(_01756_),
    .S(_01717_),
    .X(_01758_));
 sky130_fd_sc_hd__mux2_1 _40894_ (.A0(\pcpi_mul.rd[3] ),
    .A1(\pcpi_mul.rd[35] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01753_));
 sky130_fd_sc_hd__mux2_1 _40895_ (.A0(_01751_),
    .A1(_01747_),
    .S(_01683_),
    .X(_01752_));
 sky130_fd_sc_hd__mux2_1 _40896_ (.A0(mem_rdata[3]),
    .A1(mem_rdata[19]),
    .S(pcpi_rs1[1]),
    .X(_01750_));
 sky130_fd_sc_hd__mux2_1 _40897_ (.A0(_01748_),
    .A1(_01747_),
    .S(_00304_),
    .X(_01749_));
 sky130_fd_sc_hd__mux2_1 _40898_ (.A0(_01742_),
    .A1(_01741_),
    .S(_01714_),
    .X(_01743_));
 sky130_fd_sc_hd__mux2_1 _40899_ (.A0(_01744_),
    .A1(_01743_),
    .S(_01717_),
    .X(_01745_));
 sky130_fd_sc_hd__mux2_1 _40900_ (.A0(\pcpi_mul.rd[2] ),
    .A1(\pcpi_mul.rd[34] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01740_));
 sky130_fd_sc_hd__mux2_1 _40901_ (.A0(_01738_),
    .A1(_01734_),
    .S(_01683_),
    .X(_01739_));
 sky130_fd_sc_hd__mux2_1 _40902_ (.A0(mem_rdata[2]),
    .A1(mem_rdata[18]),
    .S(pcpi_rs1[1]),
    .X(_01737_));
 sky130_fd_sc_hd__mux2_1 _40903_ (.A0(_01735_),
    .A1(_01734_),
    .S(_00304_),
    .X(_01736_));
 sky130_fd_sc_hd__mux2_1 _40904_ (.A0(_01729_),
    .A1(_01728_),
    .S(_01714_),
    .X(_01730_));
 sky130_fd_sc_hd__mux2_1 _40905_ (.A0(_01731_),
    .A1(_01730_),
    .S(_01717_),
    .X(_01732_));
 sky130_fd_sc_hd__mux2_1 _40906_ (.A0(\pcpi_mul.rd[1] ),
    .A1(\pcpi_mul.rd[33] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01727_));
 sky130_fd_sc_hd__mux2_1 _40907_ (.A0(_01725_),
    .A1(_01721_),
    .S(_01683_),
    .X(_01726_));
 sky130_fd_sc_hd__mux2_1 _40908_ (.A0(mem_rdata[1]),
    .A1(mem_rdata[17]),
    .S(pcpi_rs1[1]),
    .X(_01724_));
 sky130_fd_sc_hd__mux2_1 _40909_ (.A0(_01722_),
    .A1(_01721_),
    .S(_00304_),
    .X(_01723_));
 sky130_fd_sc_hd__mux2_1 _40910_ (.A0(_01715_),
    .A1(_02559_),
    .S(_01714_),
    .X(_01716_));
 sky130_fd_sc_hd__mux2_1 _40911_ (.A0(_01718_),
    .A1(_01716_),
    .S(_01717_),
    .X(_01719_));
 sky130_fd_sc_hd__mux2_1 _40912_ (.A0(\pcpi_mul.rd[0] ),
    .A1(\pcpi_mul.rd[32] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01713_));
 sky130_fd_sc_hd__mux2_1 _40913_ (.A0(_01711_),
    .A1(_01707_),
    .S(_01683_),
    .X(_01712_));
 sky130_fd_sc_hd__mux2_1 _40914_ (.A0(mem_rdata[0]),
    .A1(mem_rdata[16]),
    .S(pcpi_rs1[1]),
    .X(_01710_));
 sky130_fd_sc_hd__mux2_1 _40915_ (.A0(_01708_),
    .A1(_01707_),
    .S(_00304_),
    .X(_01709_));
 sky130_fd_sc_hd__mux2_1 _40916_ (.A0(_01701_),
    .A1(_01696_),
    .S(_00311_),
    .X(_01702_));
 sky130_fd_sc_hd__mux2_1 _40917_ (.A0(_01702_),
    .A1(_01696_),
    .S(\pcpi_mul.active[1] ),
    .X(_01703_));
 sky130_fd_sc_hd__mux2_1 _40918_ (.A0(_01696_),
    .A1(_01703_),
    .S(_00310_),
    .X(_01704_));
 sky130_fd_sc_hd__mux2_1 _40919_ (.A0(_01693_),
    .A1(mem_wstrb[3]),
    .S(_00316_),
    .X(_01694_));
 sky130_fd_sc_hd__mux2_1 _40920_ (.A0(_01690_),
    .A1(mem_wstrb[2]),
    .S(_00316_),
    .X(_01691_));
 sky130_fd_sc_hd__mux2_1 _40921_ (.A0(_01687_),
    .A1(mem_wstrb[1]),
    .S(_00316_),
    .X(_01688_));
 sky130_fd_sc_hd__mux2_1 _40922_ (.A0(_01684_),
    .A1(mem_wstrb[0]),
    .S(_00316_),
    .X(_01685_));
 sky130_fd_sc_hd__mux2_1 _40923_ (.A0(\reg_next_pc[31] ),
    .A1(_01554_),
    .S(latched_store),
    .X(_01555_));
 sky130_fd_sc_hd__mux2_1 _40924_ (.A0(\reg_out[31] ),
    .A1(\alu_out_q[31] ),
    .S(latched_stalu),
    .X(_01554_));
 sky130_fd_sc_hd__mux2_1 _40925_ (.A0(\reg_next_pc[30] ),
    .A1(_01551_),
    .S(latched_store),
    .X(_01552_));
 sky130_fd_sc_hd__mux2_1 _40926_ (.A0(\reg_out[30] ),
    .A1(\alu_out_q[30] ),
    .S(latched_stalu),
    .X(_01551_));
 sky130_fd_sc_hd__mux2_1 _40927_ (.A0(\reg_next_pc[29] ),
    .A1(_01548_),
    .S(latched_store),
    .X(_01549_));
 sky130_fd_sc_hd__mux2_1 _40928_ (.A0(\reg_out[29] ),
    .A1(\alu_out_q[29] ),
    .S(latched_stalu),
    .X(_01548_));
 sky130_fd_sc_hd__mux2_1 _40929_ (.A0(\reg_next_pc[28] ),
    .A1(_01545_),
    .S(latched_store),
    .X(_01546_));
 sky130_fd_sc_hd__mux2_1 _40930_ (.A0(\reg_out[28] ),
    .A1(\alu_out_q[28] ),
    .S(latched_stalu),
    .X(_01545_));
 sky130_fd_sc_hd__mux2_1 _40931_ (.A0(\reg_next_pc[27] ),
    .A1(_01542_),
    .S(latched_store),
    .X(_01543_));
 sky130_fd_sc_hd__mux2_1 _40932_ (.A0(\reg_out[27] ),
    .A1(\alu_out_q[27] ),
    .S(latched_stalu),
    .X(_01542_));
 sky130_fd_sc_hd__mux2_1 _40933_ (.A0(\reg_next_pc[26] ),
    .A1(_01539_),
    .S(latched_store),
    .X(_01540_));
 sky130_fd_sc_hd__mux2_1 _40934_ (.A0(\reg_out[26] ),
    .A1(\alu_out_q[26] ),
    .S(latched_stalu),
    .X(_01539_));
 sky130_fd_sc_hd__mux2_1 _40935_ (.A0(\reg_next_pc[25] ),
    .A1(_01536_),
    .S(latched_store),
    .X(_01537_));
 sky130_fd_sc_hd__mux2_1 _40936_ (.A0(\reg_out[25] ),
    .A1(\alu_out_q[25] ),
    .S(latched_stalu),
    .X(_01536_));
 sky130_fd_sc_hd__mux2_1 _40937_ (.A0(\reg_next_pc[24] ),
    .A1(_01533_),
    .S(latched_store),
    .X(_01534_));
 sky130_fd_sc_hd__mux2_1 _40938_ (.A0(\reg_out[24] ),
    .A1(\alu_out_q[24] ),
    .S(latched_stalu),
    .X(_01533_));
 sky130_fd_sc_hd__mux2_1 _40939_ (.A0(\reg_next_pc[23] ),
    .A1(_01530_),
    .S(latched_store),
    .X(_01531_));
 sky130_fd_sc_hd__mux2_1 _40940_ (.A0(\reg_out[23] ),
    .A1(\alu_out_q[23] ),
    .S(latched_stalu),
    .X(_01530_));
 sky130_fd_sc_hd__mux2_1 _40941_ (.A0(\reg_next_pc[22] ),
    .A1(_01527_),
    .S(latched_store),
    .X(_01528_));
 sky130_fd_sc_hd__mux2_1 _40942_ (.A0(\reg_out[22] ),
    .A1(\alu_out_q[22] ),
    .S(latched_stalu),
    .X(_01527_));
 sky130_fd_sc_hd__mux2_1 _40943_ (.A0(\reg_next_pc[21] ),
    .A1(_01524_),
    .S(latched_store),
    .X(_01525_));
 sky130_fd_sc_hd__mux2_1 _40944_ (.A0(\reg_out[21] ),
    .A1(\alu_out_q[21] ),
    .S(latched_stalu),
    .X(_01524_));
 sky130_fd_sc_hd__mux2_1 _40945_ (.A0(\reg_next_pc[20] ),
    .A1(_01521_),
    .S(latched_store),
    .X(_01522_));
 sky130_fd_sc_hd__mux2_1 _40946_ (.A0(\reg_out[20] ),
    .A1(\alu_out_q[20] ),
    .S(latched_stalu),
    .X(_01521_));
 sky130_fd_sc_hd__mux2_1 _40947_ (.A0(\reg_next_pc[19] ),
    .A1(_01518_),
    .S(latched_store),
    .X(_01519_));
 sky130_fd_sc_hd__mux2_1 _40948_ (.A0(\reg_out[19] ),
    .A1(\alu_out_q[19] ),
    .S(latched_stalu),
    .X(_01518_));
 sky130_fd_sc_hd__mux2_1 _40949_ (.A0(\reg_next_pc[18] ),
    .A1(_01515_),
    .S(latched_store),
    .X(_01516_));
 sky130_fd_sc_hd__mux2_1 _40950_ (.A0(\reg_out[18] ),
    .A1(\alu_out_q[18] ),
    .S(latched_stalu),
    .X(_01515_));
 sky130_fd_sc_hd__mux2_1 _40951_ (.A0(\reg_next_pc[17] ),
    .A1(_01512_),
    .S(latched_store),
    .X(_01513_));
 sky130_fd_sc_hd__mux2_1 _40952_ (.A0(\reg_out[17] ),
    .A1(\alu_out_q[17] ),
    .S(latched_stalu),
    .X(_01512_));
 sky130_fd_sc_hd__mux2_1 _40953_ (.A0(\reg_next_pc[16] ),
    .A1(_01509_),
    .S(latched_store),
    .X(_01510_));
 sky130_fd_sc_hd__mux2_1 _40954_ (.A0(\reg_out[16] ),
    .A1(\alu_out_q[16] ),
    .S(latched_stalu),
    .X(_01509_));
 sky130_fd_sc_hd__mux2_1 _40955_ (.A0(\reg_next_pc[15] ),
    .A1(_01506_),
    .S(latched_store),
    .X(_01507_));
 sky130_fd_sc_hd__mux2_1 _40956_ (.A0(\reg_out[15] ),
    .A1(\alu_out_q[15] ),
    .S(latched_stalu),
    .X(_01506_));
 sky130_fd_sc_hd__mux2_1 _40957_ (.A0(\reg_next_pc[14] ),
    .A1(_01503_),
    .S(latched_store),
    .X(_01504_));
 sky130_fd_sc_hd__mux2_1 _40958_ (.A0(\reg_out[14] ),
    .A1(\alu_out_q[14] ),
    .S(latched_stalu),
    .X(_01503_));
 sky130_fd_sc_hd__mux2_1 _40959_ (.A0(\reg_next_pc[13] ),
    .A1(_01500_),
    .S(latched_store),
    .X(_01501_));
 sky130_fd_sc_hd__mux2_1 _40960_ (.A0(\reg_out[13] ),
    .A1(\alu_out_q[13] ),
    .S(latched_stalu),
    .X(_01500_));
 sky130_fd_sc_hd__mux2_1 _40961_ (.A0(\reg_next_pc[12] ),
    .A1(_01497_),
    .S(latched_store),
    .X(_01498_));
 sky130_fd_sc_hd__mux2_1 _40962_ (.A0(\reg_out[12] ),
    .A1(\alu_out_q[12] ),
    .S(latched_stalu),
    .X(_01497_));
 sky130_fd_sc_hd__mux2_1 _40963_ (.A0(\reg_next_pc[11] ),
    .A1(_01494_),
    .S(latched_store),
    .X(_01495_));
 sky130_fd_sc_hd__mux2_1 _40964_ (.A0(\reg_out[11] ),
    .A1(\alu_out_q[11] ),
    .S(latched_stalu),
    .X(_01494_));
 sky130_fd_sc_hd__mux2_1 _40965_ (.A0(\reg_next_pc[10] ),
    .A1(_01491_),
    .S(latched_store),
    .X(_01492_));
 sky130_fd_sc_hd__mux2_1 _40966_ (.A0(\reg_out[10] ),
    .A1(\alu_out_q[10] ),
    .S(latched_stalu),
    .X(_01491_));
 sky130_fd_sc_hd__mux2_1 _40967_ (.A0(\reg_next_pc[9] ),
    .A1(_01488_),
    .S(latched_store),
    .X(_01489_));
 sky130_fd_sc_hd__mux2_1 _40968_ (.A0(\reg_out[9] ),
    .A1(\alu_out_q[9] ),
    .S(latched_stalu),
    .X(_01488_));
 sky130_fd_sc_hd__mux2_1 _40969_ (.A0(\reg_next_pc[8] ),
    .A1(_01485_),
    .S(latched_store),
    .X(_01486_));
 sky130_fd_sc_hd__mux2_1 _40970_ (.A0(\reg_out[8] ),
    .A1(\alu_out_q[8] ),
    .S(latched_stalu),
    .X(_01485_));
 sky130_fd_sc_hd__mux2_1 _40971_ (.A0(\reg_next_pc[7] ),
    .A1(_01482_),
    .S(latched_store),
    .X(_01483_));
 sky130_fd_sc_hd__mux2_1 _40972_ (.A0(\reg_out[7] ),
    .A1(\alu_out_q[7] ),
    .S(latched_stalu),
    .X(_01482_));
 sky130_fd_sc_hd__mux2_1 _40973_ (.A0(\reg_next_pc[6] ),
    .A1(_01479_),
    .S(latched_store),
    .X(_01480_));
 sky130_fd_sc_hd__mux2_1 _40974_ (.A0(\reg_out[6] ),
    .A1(\alu_out_q[6] ),
    .S(latched_stalu),
    .X(_01479_));
 sky130_fd_sc_hd__mux2_1 _40975_ (.A0(\reg_next_pc[5] ),
    .A1(_01476_),
    .S(latched_store),
    .X(_01477_));
 sky130_fd_sc_hd__mux2_1 _40976_ (.A0(\reg_out[5] ),
    .A1(\alu_out_q[5] ),
    .S(latched_stalu),
    .X(_01476_));
 sky130_fd_sc_hd__mux2_1 _40977_ (.A0(_01474_),
    .A1(_01471_),
    .S(_00292_),
    .X(_01475_));
 sky130_fd_sc_hd__mux2_1 _40978_ (.A0(\reg_next_pc[4] ),
    .A1(_01472_),
    .S(latched_store),
    .X(_01473_));
 sky130_fd_sc_hd__mux2_1 _40979_ (.A0(\reg_out[4] ),
    .A1(\alu_out_q[4] ),
    .S(latched_stalu),
    .X(_01472_));
 sky130_fd_sc_hd__mux2_1 _40980_ (.A0(\reg_next_pc[3] ),
    .A1(_01468_),
    .S(latched_store),
    .X(_01469_));
 sky130_fd_sc_hd__mux2_1 _40981_ (.A0(\reg_out[3] ),
    .A1(\alu_out_q[3] ),
    .S(latched_stalu),
    .X(_01468_));
 sky130_fd_sc_hd__mux2_1 _40982_ (.A0(\reg_next_pc[1] ),
    .A1(_01465_),
    .S(latched_store),
    .X(_01466_));
 sky130_fd_sc_hd__mux2_1 _40983_ (.A0(\reg_out[1] ),
    .A1(\alu_out_q[1] ),
    .S(latched_stalu),
    .X(_01465_));
 sky130_fd_sc_hd__mux2_1 _40984_ (.A0(_01301_),
    .A1(\timer[31] ),
    .S(_01208_),
    .X(_01302_));
 sky130_fd_sc_hd__mux2_1 _40985_ (.A0(_01298_),
    .A1(\timer[30] ),
    .S(_01208_),
    .X(_01299_));
 sky130_fd_sc_hd__mux2_1 _40986_ (.A0(_01295_),
    .A1(\timer[29] ),
    .S(_01208_),
    .X(_01296_));
 sky130_fd_sc_hd__mux2_1 _40987_ (.A0(_01292_),
    .A1(\timer[28] ),
    .S(_01208_),
    .X(_01293_));
 sky130_fd_sc_hd__mux2_1 _40988_ (.A0(_01289_),
    .A1(\timer[27] ),
    .S(_01208_),
    .X(_01290_));
 sky130_fd_sc_hd__mux2_1 _40989_ (.A0(_01286_),
    .A1(\timer[26] ),
    .S(_01208_),
    .X(_01287_));
 sky130_fd_sc_hd__mux2_1 _40990_ (.A0(_01283_),
    .A1(\timer[25] ),
    .S(_01208_),
    .X(_01284_));
 sky130_fd_sc_hd__mux2_1 _40991_ (.A0(_01280_),
    .A1(\timer[24] ),
    .S(_01208_),
    .X(_01281_));
 sky130_fd_sc_hd__mux2_1 _40992_ (.A0(_01277_),
    .A1(\timer[23] ),
    .S(_01208_),
    .X(_01278_));
 sky130_fd_sc_hd__mux2_1 _40993_ (.A0(_01274_),
    .A1(\timer[22] ),
    .S(_01208_),
    .X(_01275_));
 sky130_fd_sc_hd__mux2_1 _40994_ (.A0(_01271_),
    .A1(\timer[21] ),
    .S(_01208_),
    .X(_01272_));
 sky130_fd_sc_hd__mux2_1 _40995_ (.A0(_01268_),
    .A1(\timer[20] ),
    .S(_01208_),
    .X(_01269_));
 sky130_fd_sc_hd__mux2_1 _40996_ (.A0(_01265_),
    .A1(\timer[19] ),
    .S(_01208_),
    .X(_01266_));
 sky130_fd_sc_hd__mux2_1 _40997_ (.A0(_01262_),
    .A1(\timer[18] ),
    .S(_01208_),
    .X(_01263_));
 sky130_fd_sc_hd__mux2_1 _40998_ (.A0(_01259_),
    .A1(\timer[17] ),
    .S(_01208_),
    .X(_01260_));
 sky130_fd_sc_hd__mux2_1 _40999_ (.A0(_01256_),
    .A1(\timer[16] ),
    .S(_01208_),
    .X(_01257_));
 sky130_fd_sc_hd__mux2_1 _41000_ (.A0(_01253_),
    .A1(\timer[15] ),
    .S(_01208_),
    .X(_01254_));
 sky130_fd_sc_hd__mux2_1 _41001_ (.A0(_01250_),
    .A1(\timer[14] ),
    .S(_01208_),
    .X(_01251_));
 sky130_fd_sc_hd__mux2_1 _41002_ (.A0(_01247_),
    .A1(\timer[13] ),
    .S(_01208_),
    .X(_01248_));
 sky130_fd_sc_hd__mux2_1 _41003_ (.A0(_01244_),
    .A1(\timer[12] ),
    .S(_01208_),
    .X(_01245_));
 sky130_fd_sc_hd__mux2_1 _41004_ (.A0(_01241_),
    .A1(\timer[11] ),
    .S(_01208_),
    .X(_01242_));
 sky130_fd_sc_hd__mux2_1 _41005_ (.A0(_01238_),
    .A1(\timer[10] ),
    .S(_01208_),
    .X(_01239_));
 sky130_fd_sc_hd__mux2_1 _41006_ (.A0(_01235_),
    .A1(\timer[9] ),
    .S(_01208_),
    .X(_01236_));
 sky130_fd_sc_hd__mux2_1 _41007_ (.A0(_01232_),
    .A1(\timer[8] ),
    .S(_01208_),
    .X(_01233_));
 sky130_fd_sc_hd__mux2_1 _41008_ (.A0(_01229_),
    .A1(\timer[7] ),
    .S(_01208_),
    .X(_01230_));
 sky130_fd_sc_hd__mux2_1 _41009_ (.A0(_01226_),
    .A1(\timer[6] ),
    .S(_01208_),
    .X(_01227_));
 sky130_fd_sc_hd__mux2_1 _41010_ (.A0(_01223_),
    .A1(\timer[5] ),
    .S(_01208_),
    .X(_01224_));
 sky130_fd_sc_hd__mux2_1 _41011_ (.A0(_01220_),
    .A1(\timer[4] ),
    .S(_01208_),
    .X(_01221_));
 sky130_fd_sc_hd__mux2_1 _41012_ (.A0(_01217_),
    .A1(\timer[3] ),
    .S(_01208_),
    .X(_01218_));
 sky130_fd_sc_hd__mux2_1 _41013_ (.A0(_01214_),
    .A1(\timer[2] ),
    .S(_01208_),
    .X(_01215_));
 sky130_fd_sc_hd__mux2_1 _41014_ (.A0(_01211_),
    .A1(\timer[1] ),
    .S(_01208_),
    .X(_01212_));
 sky130_fd_sc_hd__mux2_1 _41015_ (.A0(_01206_),
    .A1(_01201_),
    .S(_00368_),
    .X(_01207_));
 sky130_fd_sc_hd__mux2_1 _41016_ (.A0(_01179_),
    .A1(_01174_),
    .S(_00368_),
    .X(_01180_));
 sky130_fd_sc_hd__mux2_1 _41017_ (.A0(_01152_),
    .A1(_01147_),
    .S(_00368_),
    .X(_01153_));
 sky130_fd_sc_hd__mux2_1 _41018_ (.A0(_01125_),
    .A1(_01120_),
    .S(_00368_),
    .X(_01126_));
 sky130_fd_sc_hd__mux2_1 _41019_ (.A0(_01098_),
    .A1(_01093_),
    .S(_00368_),
    .X(_01099_));
 sky130_fd_sc_hd__mux2_1 _41020_ (.A0(_01071_),
    .A1(_01066_),
    .S(_00368_),
    .X(_01072_));
 sky130_fd_sc_hd__mux2_1 _41021_ (.A0(_01044_),
    .A1(_01039_),
    .S(_00368_),
    .X(_01045_));
 sky130_fd_sc_hd__mux2_1 _41022_ (.A0(_01017_),
    .A1(_01012_),
    .S(_00368_),
    .X(_01018_));
 sky130_fd_sc_hd__mux2_1 _41023_ (.A0(_00990_),
    .A1(_00985_),
    .S(_00368_),
    .X(_00991_));
 sky130_fd_sc_hd__mux2_1 _41024_ (.A0(_00963_),
    .A1(_00958_),
    .S(_00368_),
    .X(_00964_));
 sky130_fd_sc_hd__mux2_1 _41025_ (.A0(_00936_),
    .A1(_00931_),
    .S(_00368_),
    .X(_00937_));
 sky130_fd_sc_hd__mux2_1 _41026_ (.A0(_00909_),
    .A1(_00904_),
    .S(_00368_),
    .X(_00910_));
 sky130_fd_sc_hd__mux2_1 _41027_ (.A0(_00882_),
    .A1(_00877_),
    .S(_00368_),
    .X(_00883_));
 sky130_fd_sc_hd__mux2_1 _41028_ (.A0(_00855_),
    .A1(_00850_),
    .S(_00368_),
    .X(_00856_));
 sky130_fd_sc_hd__mux2_1 _41029_ (.A0(_00828_),
    .A1(_00823_),
    .S(_00368_),
    .X(_00829_));
 sky130_fd_sc_hd__mux2_1 _41030_ (.A0(_00801_),
    .A1(_00796_),
    .S(_00368_),
    .X(_00802_));
 sky130_fd_sc_hd__mux2_1 _41031_ (.A0(_00774_),
    .A1(_00769_),
    .S(_00368_),
    .X(_00775_));
 sky130_fd_sc_hd__mux2_1 _41032_ (.A0(_00747_),
    .A1(_00742_),
    .S(_00368_),
    .X(_00748_));
 sky130_fd_sc_hd__mux2_1 _41033_ (.A0(_00720_),
    .A1(_00715_),
    .S(_00368_),
    .X(_00721_));
 sky130_fd_sc_hd__mux2_1 _41034_ (.A0(_00693_),
    .A1(_00688_),
    .S(_00368_),
    .X(_00694_));
 sky130_fd_sc_hd__mux2_1 _41035_ (.A0(_00666_),
    .A1(_00661_),
    .S(_00368_),
    .X(_00667_));
 sky130_fd_sc_hd__mux2_1 _41036_ (.A0(_00639_),
    .A1(_00634_),
    .S(_00368_),
    .X(_00640_));
 sky130_fd_sc_hd__mux2_1 _41037_ (.A0(_00612_),
    .A1(_00607_),
    .S(_00368_),
    .X(_00613_));
 sky130_fd_sc_hd__mux2_1 _41038_ (.A0(_00585_),
    .A1(_00580_),
    .S(_00368_),
    .X(_00586_));
 sky130_fd_sc_hd__mux2_1 _41039_ (.A0(_00558_),
    .A1(_00553_),
    .S(_00368_),
    .X(_00559_));
 sky130_fd_sc_hd__mux2_1 _41040_ (.A0(_00531_),
    .A1(_00526_),
    .S(_00368_),
    .X(_00532_));
 sky130_fd_sc_hd__mux2_1 _41041_ (.A0(_00504_),
    .A1(_00499_),
    .S(_00368_),
    .X(_00505_));
 sky130_fd_sc_hd__mux2_1 _41042_ (.A0(_00477_),
    .A1(_00472_),
    .S(_00368_),
    .X(_00478_));
 sky130_fd_sc_hd__mux2_1 _41043_ (.A0(_00450_),
    .A1(_00445_),
    .S(_00368_),
    .X(_00451_));
 sky130_fd_sc_hd__mux2_1 _41044_ (.A0(_00423_),
    .A1(_00418_),
    .S(_00368_),
    .X(_00424_));
 sky130_fd_sc_hd__mux2_1 _41045_ (.A0(_00396_),
    .A1(_00391_),
    .S(_00368_),
    .X(_00397_));
 sky130_fd_sc_hd__mux2_1 _41046_ (.A0(_00369_),
    .A1(_00365_),
    .S(_00368_),
    .X(_00370_));
 sky130_fd_sc_hd__mux2_1 _41047_ (.A0(_00366_),
    .A1(_00367_),
    .S(\cpu_state[3] ),
    .X(_00368_));
 sky130_fd_sc_hd__mux2_1 _41048_ (.A0(\decoded_rs1[3] ),
    .A1(\decoded_imm_uj[3] ),
    .S(\cpu_state[3] ),
    .X(_00362_));
 sky130_fd_sc_hd__mux2_1 _41049_ (.A0(\decoded_rs1[2] ),
    .A1(\decoded_imm_uj[2] ),
    .S(\cpu_state[3] ),
    .X(_00360_));
 sky130_fd_sc_hd__mux2_1 _41050_ (.A0(\decoded_rs1[1] ),
    .A1(\decoded_imm_uj[1] ),
    .S(\cpu_state[3] ),
    .X(_00358_));
 sky130_fd_sc_hd__mux2_1 _41051_ (.A0(\decoded_rs1[0] ),
    .A1(\decoded_imm_uj[11] ),
    .S(\cpu_state[3] ),
    .X(_00357_));
 sky130_fd_sc_hd__mux2_1 _41052_ (.A0(_00349_),
    .A1(_00323_),
    .S(decoder_trigger),
    .X(_00350_));
 sky130_fd_sc_hd__mux2_1 _41053_ (.A0(_00350_),
    .A1(_00351_),
    .S(_00309_),
    .X(_00352_));
 sky130_fd_sc_hd__mux2_1 _41054_ (.A0(_00352_),
    .A1(_00349_),
    .S(_00308_),
    .X(_00353_));
 sky130_fd_sc_hd__mux2_1 _41055_ (.A0(_00355_),
    .A1(_00353_),
    .S(_00354_),
    .X(_00356_));
 sky130_fd_sc_hd__mux2_1 _41056_ (.A0(_00337_),
    .A1(_00344_),
    .S(is_beq_bne_blt_bge_bltu_bgeu),
    .X(_00345_));
 sky130_fd_sc_hd__mux2_1 _41057_ (.A0(_00345_),
    .A1(_00337_),
    .S(alu_wait),
    .X(_00346_));
 sky130_fd_sc_hd__mux2_1 _41058_ (.A0(_00342_),
    .A1(_00340_),
    .S(_00341_),
    .X(_00343_));
 sky130_fd_sc_hd__mux2_1 _41059_ (.A0(_00338_),
    .A1(_00337_),
    .S(_00296_),
    .X(_00339_));
 sky130_fd_sc_hd__mux2_1 _41060_ (.A0(\mem_rdata_q[12] ),
    .A1(_00334_),
    .S(\mem_rdata_q[13] ),
    .X(_00335_));
 sky130_fd_sc_hd__mux2_1 _41061_ (.A0(\cpu_state[1] ),
    .A1(_00302_),
    .S(\cpu_state[4] ),
    .X(_00333_));
 sky130_fd_sc_hd__mux2_1 _41062_ (.A0(_00322_),
    .A1(_00296_),
    .S(\cpu_state[6] ),
    .X(_00332_));
 sky130_fd_sc_hd__mux2_1 _41063_ (.A0(_00315_),
    .A1(alu_wait),
    .S(\cpu_state[4] ),
    .X(_00331_));
 sky130_fd_sc_hd__mux2_1 _41064_ (.A0(\mem_rdata_q[6] ),
    .A1(mem_rdata[6]),
    .S(mem_xfer),
    .X(_00330_));
 sky130_fd_sc_hd__mux2_1 _41065_ (.A0(\mem_rdata_q[5] ),
    .A1(mem_rdata[5]),
    .S(mem_xfer),
    .X(_00329_));
 sky130_fd_sc_hd__mux2_1 _41066_ (.A0(\mem_rdata_q[4] ),
    .A1(mem_rdata[4]),
    .S(mem_xfer),
    .X(_00328_));
 sky130_fd_sc_hd__mux2_1 _41067_ (.A0(\mem_rdata_q[3] ),
    .A1(mem_rdata[3]),
    .S(mem_xfer),
    .X(_00327_));
 sky130_fd_sc_hd__mux2_1 _41068_ (.A0(\mem_rdata_q[2] ),
    .A1(mem_rdata[2]),
    .S(mem_xfer),
    .X(_00326_));
 sky130_fd_sc_hd__mux2_1 _41069_ (.A0(\mem_rdata_q[1] ),
    .A1(mem_rdata[1]),
    .S(mem_xfer),
    .X(_00325_));
 sky130_fd_sc_hd__mux2_1 _41070_ (.A0(\mem_rdata_q[0] ),
    .A1(mem_rdata[0]),
    .S(mem_xfer),
    .X(_00324_));
 sky130_fd_sc_hd__mux2_1 _41071_ (.A0(\cpu_state[1] ),
    .A1(instr_retirq),
    .S(\cpu_state[2] ),
    .X(_00321_));
 sky130_fd_sc_hd__mux2_1 _41072_ (.A0(_00319_),
    .A1(\cpu_state[5] ),
    .S(_00296_),
    .X(_00320_));
 sky130_fd_sc_hd__mux2_1 _41073_ (.A0(_00317_),
    .A1(\cpu_state[6] ),
    .S(_00296_),
    .X(_00318_));
 sky130_fd_sc_hd__mux2_1 _41074_ (.A0(_00313_),
    .A1(_00312_),
    .S(_00307_),
    .X(_00314_));
 sky130_fd_sc_hd__mux2_1 _41075_ (.A0(_00298_),
    .A1(_00299_),
    .S(_00289_),
    .X(_00300_));
 sky130_fd_sc_hd__mux2_1 _41076_ (.A0(\reg_next_pc[2] ),
    .A1(_00293_),
    .S(latched_store),
    .X(_00294_));
 sky130_fd_sc_hd__mux2_1 _41077_ (.A0(\reg_out[2] ),
    .A1(\alu_out_q[2] ),
    .S(latched_stalu),
    .X(_00293_));
 sky130_fd_sc_hd__mux2_1 _41078_ (.A0(_00126_),
    .A1(_00122_),
    .S(mem_la_wdata[3]),
    .X(_02558_));
 sky130_fd_sc_hd__mux2_1 _41079_ (.A0(_00120_),
    .A1(_00116_),
    .S(mem_la_wdata[3]),
    .X(_02557_));
 sky130_fd_sc_hd__mux2_1 _41080_ (.A0(_00114_),
    .A1(_00110_),
    .S(mem_la_wdata[3]),
    .X(_02556_));
 sky130_fd_sc_hd__mux2_1 _41081_ (.A0(_00108_),
    .A1(_00104_),
    .S(mem_la_wdata[3]),
    .X(_02555_));
 sky130_fd_sc_hd__mux2_1 _41082_ (.A0(_00102_),
    .A1(_00095_),
    .S(mem_la_wdata[3]),
    .X(_02554_));
 sky130_fd_sc_hd__mux2_1 _41083_ (.A0(_00092_),
    .A1(_00085_),
    .S(mem_la_wdata[3]),
    .X(_02553_));
 sky130_fd_sc_hd__mux2_1 _41084_ (.A0(_00082_),
    .A1(_00068_),
    .S(mem_la_wdata[3]),
    .X(_02552_));
 sky130_fd_sc_hd__mux2_1 _41085_ (.A0(_00064_),
    .A1(_00050_),
    .S(mem_la_wdata[3]),
    .X(_02551_));
 sky130_fd_sc_hd__mux2_1 _41086_ (.A0(_01694_),
    .A1(_01695_),
    .S(_00290_),
    .X(_02541_));
 sky130_fd_sc_hd__mux2_1 _41087_ (.A0(_01691_),
    .A1(_01692_),
    .S(_00290_),
    .X(_02540_));
 sky130_fd_sc_hd__mux2_1 _41088_ (.A0(_01688_),
    .A1(_01689_),
    .S(_00290_),
    .X(_02539_));
 sky130_fd_sc_hd__mux2_1 _41089_ (.A0(_01685_),
    .A1(_01686_),
    .S(_00290_),
    .X(_02538_));
 sky130_fd_sc_hd__mux2_1 _41090_ (.A0(_01679_),
    .A1(_01680_),
    .S(instr_jal),
    .X(_01681_));
 sky130_fd_sc_hd__mux2_1 _41091_ (.A0(_01682_),
    .A1(_02581_),
    .S(_00308_),
    .X(_02530_));
 sky130_fd_sc_hd__mux2_1 _41092_ (.A0(_01675_),
    .A1(_01676_),
    .S(instr_jal),
    .X(_01677_));
 sky130_fd_sc_hd__mux2_1 _41093_ (.A0(_01678_),
    .A1(_02580_),
    .S(_00308_),
    .X(_02529_));
 sky130_fd_sc_hd__mux2_1 _41094_ (.A0(_01671_),
    .A1(_01672_),
    .S(instr_jal),
    .X(_01673_));
 sky130_fd_sc_hd__mux2_1 _41095_ (.A0(_01674_),
    .A1(_02579_),
    .S(_00308_),
    .X(_02527_));
 sky130_fd_sc_hd__mux2_1 _41096_ (.A0(_01667_),
    .A1(_01668_),
    .S(instr_jal),
    .X(_01669_));
 sky130_fd_sc_hd__mux2_1 _41097_ (.A0(_01670_),
    .A1(_02578_),
    .S(_00308_),
    .X(_02526_));
 sky130_fd_sc_hd__mux2_1 _41098_ (.A0(_01663_),
    .A1(_01664_),
    .S(instr_jal),
    .X(_01665_));
 sky130_fd_sc_hd__mux2_1 _41099_ (.A0(_01666_),
    .A1(_02577_),
    .S(_00308_),
    .X(_02525_));
 sky130_fd_sc_hd__mux2_1 _41100_ (.A0(_01659_),
    .A1(_01660_),
    .S(instr_jal),
    .X(_01661_));
 sky130_fd_sc_hd__mux2_1 _41101_ (.A0(_01662_),
    .A1(_02576_),
    .S(_00308_),
    .X(_02524_));
 sky130_fd_sc_hd__mux2_1 _41102_ (.A0(_01655_),
    .A1(_01656_),
    .S(instr_jal),
    .X(_01657_));
 sky130_fd_sc_hd__mux2_1 _41103_ (.A0(_01658_),
    .A1(_02575_),
    .S(_00308_),
    .X(_02523_));
 sky130_fd_sc_hd__mux2_1 _41104_ (.A0(_01651_),
    .A1(_01652_),
    .S(instr_jal),
    .X(_01653_));
 sky130_fd_sc_hd__mux2_1 _41105_ (.A0(_01654_),
    .A1(_02574_),
    .S(_00308_),
    .X(_02522_));
 sky130_fd_sc_hd__mux2_1 _41106_ (.A0(_01647_),
    .A1(_01648_),
    .S(instr_jal),
    .X(_01649_));
 sky130_fd_sc_hd__mux2_1 _41107_ (.A0(_01650_),
    .A1(_02573_),
    .S(_00308_),
    .X(_02521_));
 sky130_fd_sc_hd__mux2_1 _41108_ (.A0(_01643_),
    .A1(_01644_),
    .S(instr_jal),
    .X(_01645_));
 sky130_fd_sc_hd__mux2_1 _41109_ (.A0(_01646_),
    .A1(_02572_),
    .S(_00308_),
    .X(_02520_));
 sky130_fd_sc_hd__mux2_1 _41110_ (.A0(_01639_),
    .A1(_01640_),
    .S(instr_jal),
    .X(_01641_));
 sky130_fd_sc_hd__mux2_1 _41111_ (.A0(_01642_),
    .A1(_02570_),
    .S(_00308_),
    .X(_02519_));
 sky130_fd_sc_hd__mux2_1 _41112_ (.A0(_01635_),
    .A1(_01636_),
    .S(instr_jal),
    .X(_01637_));
 sky130_fd_sc_hd__mux2_1 _41113_ (.A0(_01638_),
    .A1(_02569_),
    .S(_00308_),
    .X(_02518_));
 sky130_fd_sc_hd__mux2_1 _41114_ (.A0(_01631_),
    .A1(_01632_),
    .S(instr_jal),
    .X(_01633_));
 sky130_fd_sc_hd__mux2_1 _41115_ (.A0(_01634_),
    .A1(_02568_),
    .S(_00308_),
    .X(_02516_));
 sky130_fd_sc_hd__mux2_1 _41116_ (.A0(_01627_),
    .A1(_01628_),
    .S(instr_jal),
    .X(_01629_));
 sky130_fd_sc_hd__mux2_1 _41117_ (.A0(_01630_),
    .A1(_02567_),
    .S(_00308_),
    .X(_02515_));
 sky130_fd_sc_hd__mux2_1 _41118_ (.A0(_01623_),
    .A1(_01624_),
    .S(instr_jal),
    .X(_01625_));
 sky130_fd_sc_hd__mux2_1 _41119_ (.A0(_01626_),
    .A1(_02566_),
    .S(_00308_),
    .X(_02514_));
 sky130_fd_sc_hd__mux2_1 _41120_ (.A0(_01619_),
    .A1(_01620_),
    .S(instr_jal),
    .X(_01621_));
 sky130_fd_sc_hd__mux2_1 _41121_ (.A0(_01622_),
    .A1(_02565_),
    .S(_00308_),
    .X(_02513_));
 sky130_fd_sc_hd__mux2_1 _41122_ (.A0(_01615_),
    .A1(_01616_),
    .S(instr_jal),
    .X(_01617_));
 sky130_fd_sc_hd__mux2_1 _41123_ (.A0(_01618_),
    .A1(_02564_),
    .S(_00308_),
    .X(_02512_));
 sky130_fd_sc_hd__mux2_1 _41124_ (.A0(_01611_),
    .A1(_01612_),
    .S(instr_jal),
    .X(_01613_));
 sky130_fd_sc_hd__mux2_1 _41125_ (.A0(_01614_),
    .A1(_02563_),
    .S(_00308_),
    .X(_02511_));
 sky130_fd_sc_hd__mux2_1 _41126_ (.A0(_01607_),
    .A1(_01608_),
    .S(instr_jal),
    .X(_01609_));
 sky130_fd_sc_hd__mux2_1 _41127_ (.A0(_01610_),
    .A1(_02562_),
    .S(_00308_),
    .X(_02510_));
 sky130_fd_sc_hd__mux2_1 _41128_ (.A0(_01603_),
    .A1(_01604_),
    .S(instr_jal),
    .X(_01605_));
 sky130_fd_sc_hd__mux2_1 _41129_ (.A0(_01606_),
    .A1(_02561_),
    .S(_00308_),
    .X(_02509_));
 sky130_fd_sc_hd__mux2_1 _41130_ (.A0(_01599_),
    .A1(_01600_),
    .S(instr_jal),
    .X(_01601_));
 sky130_fd_sc_hd__mux2_1 _41131_ (.A0(_01602_),
    .A1(_02589_),
    .S(_00308_),
    .X(_02508_));
 sky130_fd_sc_hd__mux2_1 _41132_ (.A0(_01595_),
    .A1(_01596_),
    .S(instr_jal),
    .X(_01597_));
 sky130_fd_sc_hd__mux2_1 _41133_ (.A0(_01598_),
    .A1(_02588_),
    .S(_00308_),
    .X(_02507_));
 sky130_fd_sc_hd__mux2_1 _41134_ (.A0(_01591_),
    .A1(_01592_),
    .S(instr_jal),
    .X(_01593_));
 sky130_fd_sc_hd__mux2_1 _41135_ (.A0(_01594_),
    .A1(_02587_),
    .S(_00308_),
    .X(_02537_));
 sky130_fd_sc_hd__mux2_1 _41136_ (.A0(_01587_),
    .A1(_01588_),
    .S(instr_jal),
    .X(_01589_));
 sky130_fd_sc_hd__mux2_1 _41137_ (.A0(_01590_),
    .A1(_02586_),
    .S(_00308_),
    .X(_02536_));
 sky130_fd_sc_hd__mux2_1 _41138_ (.A0(_01583_),
    .A1(_01584_),
    .S(instr_jal),
    .X(_01585_));
 sky130_fd_sc_hd__mux2_1 _41139_ (.A0(_01586_),
    .A1(_02585_),
    .S(_00308_),
    .X(_02535_));
 sky130_fd_sc_hd__mux2_1 _41140_ (.A0(_01579_),
    .A1(_01580_),
    .S(instr_jal),
    .X(_01581_));
 sky130_fd_sc_hd__mux2_1 _41141_ (.A0(_01582_),
    .A1(_02584_),
    .S(_00308_),
    .X(_02534_));
 sky130_fd_sc_hd__mux2_1 _41142_ (.A0(_01575_),
    .A1(_01576_),
    .S(instr_jal),
    .X(_01577_));
 sky130_fd_sc_hd__mux2_1 _41143_ (.A0(_01578_),
    .A1(_02583_),
    .S(_00308_),
    .X(_02533_));
 sky130_fd_sc_hd__mux2_1 _41144_ (.A0(_01571_),
    .A1(_01572_),
    .S(instr_jal),
    .X(_01573_));
 sky130_fd_sc_hd__mux2_1 _41145_ (.A0(_01574_),
    .A1(_02582_),
    .S(_00308_),
    .X(_02532_));
 sky130_fd_sc_hd__mux2_1 _41146_ (.A0(_01567_),
    .A1(_01568_),
    .S(instr_jal),
    .X(_01569_));
 sky130_fd_sc_hd__mux2_1 _41147_ (.A0(_01570_),
    .A1(_02571_),
    .S(_00308_),
    .X(_02531_));
 sky130_fd_sc_hd__mux2_1 _41148_ (.A0(_01561_),
    .A1(_01562_),
    .S(instr_jal),
    .X(_01563_));
 sky130_fd_sc_hd__mux2_1 _41149_ (.A0(_02560_),
    .A1(_01563_),
    .S(decoder_trigger),
    .X(_01564_));
 sky130_fd_sc_hd__mux2_1 _41150_ (.A0(_01564_),
    .A1(_01565_),
    .S(_00309_),
    .X(_01566_));
 sky130_fd_sc_hd__mux2_1 _41151_ (.A0(_01566_),
    .A1(_02560_),
    .S(_00308_),
    .X(_02528_));
 sky130_fd_sc_hd__mux2_1 _41152_ (.A0(_02590_),
    .A1(_01557_),
    .S(instr_jal),
    .X(_01558_));
 sky130_fd_sc_hd__mux2_1 _41153_ (.A0(_02590_),
    .A1(_01558_),
    .S(decoder_trigger),
    .X(_01559_));
 sky130_fd_sc_hd__mux2_1 _41154_ (.A0(_01559_),
    .A1(_02590_),
    .S(_00309_),
    .X(_01560_));
 sky130_fd_sc_hd__mux2_1 _41155_ (.A0(_01560_),
    .A1(_02590_),
    .S(_00308_),
    .X(_02517_));
 sky130_fd_sc_hd__mux2_1 _41156_ (.A0(\cpuregs_rs1[31] ),
    .A1(_01462_),
    .S(is_lui_auipc_jal),
    .X(_01463_));
 sky130_fd_sc_hd__mux2_1 _41157_ (.A0(_01464_),
    .A1(_01463_),
    .S(_00297_),
    .X(_02499_));
 sky130_fd_sc_hd__mux2_1 _41158_ (.A0(\cpuregs_rs1[30] ),
    .A1(_01459_),
    .S(is_lui_auipc_jal),
    .X(_01460_));
 sky130_fd_sc_hd__mux2_1 _41159_ (.A0(_01461_),
    .A1(_01460_),
    .S(_00297_),
    .X(_02498_));
 sky130_fd_sc_hd__mux2_1 _41160_ (.A0(\cpuregs_rs1[29] ),
    .A1(_01456_),
    .S(is_lui_auipc_jal),
    .X(_01457_));
 sky130_fd_sc_hd__mux2_1 _41161_ (.A0(_01458_),
    .A1(_01457_),
    .S(_00297_),
    .X(_02496_));
 sky130_fd_sc_hd__mux2_1 _41162_ (.A0(\cpuregs_rs1[28] ),
    .A1(_01453_),
    .S(is_lui_auipc_jal),
    .X(_01454_));
 sky130_fd_sc_hd__mux2_1 _41163_ (.A0(_01455_),
    .A1(_01454_),
    .S(_00297_),
    .X(_02495_));
 sky130_fd_sc_hd__mux2_1 _41164_ (.A0(\cpuregs_rs1[27] ),
    .A1(_01450_),
    .S(is_lui_auipc_jal),
    .X(_01451_));
 sky130_fd_sc_hd__mux2_1 _41165_ (.A0(_01452_),
    .A1(_01451_),
    .S(_00297_),
    .X(_02494_));
 sky130_fd_sc_hd__mux2_1 _41166_ (.A0(\cpuregs_rs1[26] ),
    .A1(_01447_),
    .S(is_lui_auipc_jal),
    .X(_01448_));
 sky130_fd_sc_hd__mux2_1 _41167_ (.A0(_01449_),
    .A1(_01448_),
    .S(_00297_),
    .X(_02493_));
 sky130_fd_sc_hd__mux2_1 _41168_ (.A0(\cpuregs_rs1[25] ),
    .A1(_01444_),
    .S(is_lui_auipc_jal),
    .X(_01445_));
 sky130_fd_sc_hd__mux2_1 _41169_ (.A0(_01446_),
    .A1(_01445_),
    .S(_00297_),
    .X(_02492_));
 sky130_fd_sc_hd__mux2_1 _41170_ (.A0(\cpuregs_rs1[24] ),
    .A1(_01441_),
    .S(is_lui_auipc_jal),
    .X(_01442_));
 sky130_fd_sc_hd__mux2_1 _41171_ (.A0(_01443_),
    .A1(_01442_),
    .S(_00297_),
    .X(_02491_));
 sky130_fd_sc_hd__mux2_1 _41172_ (.A0(\cpuregs_rs1[23] ),
    .A1(_01438_),
    .S(is_lui_auipc_jal),
    .X(_01439_));
 sky130_fd_sc_hd__mux2_1 _41173_ (.A0(_01440_),
    .A1(_01439_),
    .S(_00297_),
    .X(_02490_));
 sky130_fd_sc_hd__mux2_1 _41174_ (.A0(\cpuregs_rs1[22] ),
    .A1(_01435_),
    .S(is_lui_auipc_jal),
    .X(_01436_));
 sky130_fd_sc_hd__mux2_1 _41175_ (.A0(_01437_),
    .A1(_01436_),
    .S(_00297_),
    .X(_02489_));
 sky130_fd_sc_hd__mux2_1 _41176_ (.A0(\cpuregs_rs1[21] ),
    .A1(_01432_),
    .S(is_lui_auipc_jal),
    .X(_01433_));
 sky130_fd_sc_hd__mux2_1 _41177_ (.A0(_01434_),
    .A1(_01433_),
    .S(_00297_),
    .X(_02488_));
 sky130_fd_sc_hd__mux2_1 _41178_ (.A0(\cpuregs_rs1[20] ),
    .A1(_01429_),
    .S(is_lui_auipc_jal),
    .X(_01430_));
 sky130_fd_sc_hd__mux2_1 _41179_ (.A0(_01431_),
    .A1(_01430_),
    .S(_00297_),
    .X(_02487_));
 sky130_fd_sc_hd__mux2_1 _41180_ (.A0(\cpuregs_rs1[19] ),
    .A1(_01426_),
    .S(is_lui_auipc_jal),
    .X(_01427_));
 sky130_fd_sc_hd__mux2_1 _41181_ (.A0(_01428_),
    .A1(_01427_),
    .S(_00297_),
    .X(_02485_));
 sky130_fd_sc_hd__mux2_1 _41182_ (.A0(\cpuregs_rs1[18] ),
    .A1(_01423_),
    .S(is_lui_auipc_jal),
    .X(_01424_));
 sky130_fd_sc_hd__mux2_1 _41183_ (.A0(_01425_),
    .A1(_01424_),
    .S(_00297_),
    .X(_02484_));
 sky130_fd_sc_hd__mux2_1 _41184_ (.A0(\cpuregs_rs1[17] ),
    .A1(_01420_),
    .S(is_lui_auipc_jal),
    .X(_01421_));
 sky130_fd_sc_hd__mux2_1 _41185_ (.A0(_01422_),
    .A1(_01421_),
    .S(_00297_),
    .X(_02483_));
 sky130_fd_sc_hd__mux2_1 _41186_ (.A0(\cpuregs_rs1[16] ),
    .A1(_01417_),
    .S(is_lui_auipc_jal),
    .X(_01418_));
 sky130_fd_sc_hd__mux2_1 _41187_ (.A0(_01419_),
    .A1(_01418_),
    .S(_00297_),
    .X(_02482_));
 sky130_fd_sc_hd__mux2_1 _41188_ (.A0(\cpuregs_rs1[15] ),
    .A1(_01414_),
    .S(is_lui_auipc_jal),
    .X(_01415_));
 sky130_fd_sc_hd__mux2_1 _41189_ (.A0(_01416_),
    .A1(_01415_),
    .S(_00297_),
    .X(_02481_));
 sky130_fd_sc_hd__mux2_1 _41190_ (.A0(\cpuregs_rs1[14] ),
    .A1(_01411_),
    .S(is_lui_auipc_jal),
    .X(_01412_));
 sky130_fd_sc_hd__mux2_1 _41191_ (.A0(_01413_),
    .A1(_01412_),
    .S(_00297_),
    .X(_02480_));
 sky130_fd_sc_hd__mux2_1 _41192_ (.A0(\cpuregs_rs1[13] ),
    .A1(_01408_),
    .S(is_lui_auipc_jal),
    .X(_01409_));
 sky130_fd_sc_hd__mux2_1 _41193_ (.A0(_01410_),
    .A1(_01409_),
    .S(_00297_),
    .X(_02479_));
 sky130_fd_sc_hd__mux2_1 _41194_ (.A0(\cpuregs_rs1[12] ),
    .A1(_01405_),
    .S(is_lui_auipc_jal),
    .X(_01406_));
 sky130_fd_sc_hd__mux2_1 _41195_ (.A0(_01407_),
    .A1(_01406_),
    .S(_00297_),
    .X(_02478_));
 sky130_fd_sc_hd__mux2_1 _41196_ (.A0(\cpuregs_rs1[11] ),
    .A1(_01402_),
    .S(is_lui_auipc_jal),
    .X(_01403_));
 sky130_fd_sc_hd__mux2_1 _41197_ (.A0(_01404_),
    .A1(_01403_),
    .S(_00297_),
    .X(_02477_));
 sky130_fd_sc_hd__mux2_1 _41198_ (.A0(\cpuregs_rs1[10] ),
    .A1(_01399_),
    .S(is_lui_auipc_jal),
    .X(_01400_));
 sky130_fd_sc_hd__mux2_1 _41199_ (.A0(_01401_),
    .A1(_01400_),
    .S(_00297_),
    .X(_02476_));
 sky130_fd_sc_hd__mux2_1 _41200_ (.A0(\cpuregs_rs1[9] ),
    .A1(_01396_),
    .S(is_lui_auipc_jal),
    .X(_01397_));
 sky130_fd_sc_hd__mux2_1 _41201_ (.A0(_01398_),
    .A1(_01397_),
    .S(_00297_),
    .X(_02506_));
 sky130_fd_sc_hd__mux2_1 _41202_ (.A0(\cpuregs_rs1[8] ),
    .A1(_01393_),
    .S(is_lui_auipc_jal),
    .X(_01394_));
 sky130_fd_sc_hd__mux2_1 _41203_ (.A0(_01395_),
    .A1(_01394_),
    .S(_00297_),
    .X(_02505_));
 sky130_fd_sc_hd__mux2_1 _41204_ (.A0(\cpuregs_rs1[7] ),
    .A1(_01390_),
    .S(is_lui_auipc_jal),
    .X(_01391_));
 sky130_fd_sc_hd__mux2_1 _41205_ (.A0(_01392_),
    .A1(_01391_),
    .S(_00297_),
    .X(_02504_));
 sky130_fd_sc_hd__mux2_1 _41206_ (.A0(\cpuregs_rs1[6] ),
    .A1(_01387_),
    .S(is_lui_auipc_jal),
    .X(_01388_));
 sky130_fd_sc_hd__mux2_1 _41207_ (.A0(_01389_),
    .A1(_01388_),
    .S(_00297_),
    .X(_02503_));
 sky130_fd_sc_hd__mux2_1 _41208_ (.A0(\cpuregs_rs1[5] ),
    .A1(_01384_),
    .S(is_lui_auipc_jal),
    .X(_01385_));
 sky130_fd_sc_hd__mux2_1 _41209_ (.A0(_01386_),
    .A1(_01385_),
    .S(_00297_),
    .X(_02502_));
 sky130_fd_sc_hd__mux2_1 _41210_ (.A0(\cpuregs_rs1[4] ),
    .A1(_01381_),
    .S(is_lui_auipc_jal),
    .X(_01382_));
 sky130_fd_sc_hd__mux2_1 _41211_ (.A0(_01383_),
    .A1(_01382_),
    .S(_00297_),
    .X(_02501_));
 sky130_fd_sc_hd__mux2_1 _41212_ (.A0(\cpuregs_rs1[3] ),
    .A1(_01378_),
    .S(is_lui_auipc_jal),
    .X(_01379_));
 sky130_fd_sc_hd__mux2_1 _41213_ (.A0(_01380_),
    .A1(_01379_),
    .S(_00297_),
    .X(_02500_));
 sky130_fd_sc_hd__mux2_1 _41214_ (.A0(\cpuregs_rs1[2] ),
    .A1(_01375_),
    .S(is_lui_auipc_jal),
    .X(_01376_));
 sky130_fd_sc_hd__mux2_1 _41215_ (.A0(_01377_),
    .A1(_01376_),
    .S(_00297_),
    .X(_02497_));
 sky130_fd_sc_hd__mux2_1 _41216_ (.A0(\cpuregs_rs1[1] ),
    .A1(_01372_),
    .S(is_lui_auipc_jal),
    .X(_01373_));
 sky130_fd_sc_hd__mux2_1 _41217_ (.A0(_01374_),
    .A1(_01373_),
    .S(_00297_),
    .X(_02486_));
 sky130_fd_sc_hd__mux2_1 _41218_ (.A0(\cpuregs_rs1[0] ),
    .A1(_01369_),
    .S(is_lui_auipc_jal),
    .X(_01370_));
 sky130_fd_sc_hd__mux2_1 _41219_ (.A0(_01371_),
    .A1(_01370_),
    .S(_00297_),
    .X(_02475_));
 sky130_fd_sc_hd__mux2_1 _41220_ (.A0(_01367_),
    .A1(\decoded_imm[31] ),
    .S(_01304_),
    .X(_01368_));
 sky130_fd_sc_hd__mux2_1 _41221_ (.A0(_01368_),
    .A1(\cpuregs_rs1[31] ),
    .S(\cpu_state[3] ),
    .X(_02467_));
 sky130_fd_sc_hd__mux2_1 _41222_ (.A0(_01365_),
    .A1(\decoded_imm[30] ),
    .S(_01304_),
    .X(_01366_));
 sky130_fd_sc_hd__mux2_1 _41223_ (.A0(_01366_),
    .A1(\cpuregs_rs1[30] ),
    .S(\cpu_state[3] ),
    .X(_02466_));
 sky130_fd_sc_hd__mux2_1 _41224_ (.A0(_01363_),
    .A1(\decoded_imm[29] ),
    .S(_01304_),
    .X(_01364_));
 sky130_fd_sc_hd__mux2_1 _41225_ (.A0(_01364_),
    .A1(\cpuregs_rs1[29] ),
    .S(\cpu_state[3] ),
    .X(_02464_));
 sky130_fd_sc_hd__mux2_1 _41226_ (.A0(_01361_),
    .A1(\decoded_imm[28] ),
    .S(_01304_),
    .X(_01362_));
 sky130_fd_sc_hd__mux2_1 _41227_ (.A0(_01362_),
    .A1(\cpuregs_rs1[28] ),
    .S(\cpu_state[3] ),
    .X(_02463_));
 sky130_fd_sc_hd__mux2_1 _41228_ (.A0(_01359_),
    .A1(\decoded_imm[27] ),
    .S(_01304_),
    .X(_01360_));
 sky130_fd_sc_hd__mux2_1 _41229_ (.A0(_01360_),
    .A1(\cpuregs_rs1[27] ),
    .S(\cpu_state[3] ),
    .X(_02462_));
 sky130_fd_sc_hd__mux2_1 _41230_ (.A0(_01357_),
    .A1(\decoded_imm[26] ),
    .S(_01304_),
    .X(_01358_));
 sky130_fd_sc_hd__mux2_1 _41231_ (.A0(_01358_),
    .A1(\cpuregs_rs1[26] ),
    .S(\cpu_state[3] ),
    .X(_02461_));
 sky130_fd_sc_hd__mux2_1 _41232_ (.A0(_01355_),
    .A1(\decoded_imm[25] ),
    .S(_01304_),
    .X(_01356_));
 sky130_fd_sc_hd__mux2_1 _41233_ (.A0(_01356_),
    .A1(\cpuregs_rs1[25] ),
    .S(\cpu_state[3] ),
    .X(_02460_));
 sky130_fd_sc_hd__mux2_1 _41234_ (.A0(_01353_),
    .A1(\decoded_imm[24] ),
    .S(_01304_),
    .X(_01354_));
 sky130_fd_sc_hd__mux2_1 _41235_ (.A0(_01354_),
    .A1(\cpuregs_rs1[24] ),
    .S(\cpu_state[3] ),
    .X(_02459_));
 sky130_fd_sc_hd__mux2_1 _41236_ (.A0(_01351_),
    .A1(\decoded_imm[23] ),
    .S(_01304_),
    .X(_01352_));
 sky130_fd_sc_hd__mux2_1 _41237_ (.A0(_01352_),
    .A1(\cpuregs_rs1[23] ),
    .S(\cpu_state[3] ),
    .X(_02458_));
 sky130_fd_sc_hd__mux2_1 _41238_ (.A0(_01349_),
    .A1(\decoded_imm[22] ),
    .S(_01304_),
    .X(_01350_));
 sky130_fd_sc_hd__mux2_1 _41239_ (.A0(_01350_),
    .A1(\cpuregs_rs1[22] ),
    .S(\cpu_state[3] ),
    .X(_02457_));
 sky130_fd_sc_hd__mux2_1 _41240_ (.A0(_01347_),
    .A1(\decoded_imm[21] ),
    .S(_01304_),
    .X(_01348_));
 sky130_fd_sc_hd__mux2_1 _41241_ (.A0(_01348_),
    .A1(\cpuregs_rs1[21] ),
    .S(\cpu_state[3] ),
    .X(_02456_));
 sky130_fd_sc_hd__mux2_1 _41242_ (.A0(_01345_),
    .A1(\decoded_imm[20] ),
    .S(_01304_),
    .X(_01346_));
 sky130_fd_sc_hd__mux2_1 _41243_ (.A0(_01346_),
    .A1(\cpuregs_rs1[20] ),
    .S(\cpu_state[3] ),
    .X(_02455_));
 sky130_fd_sc_hd__mux2_1 _41244_ (.A0(_01343_),
    .A1(\decoded_imm[19] ),
    .S(_01304_),
    .X(_01344_));
 sky130_fd_sc_hd__mux2_1 _41245_ (.A0(_01344_),
    .A1(\cpuregs_rs1[19] ),
    .S(\cpu_state[3] ),
    .X(_02453_));
 sky130_fd_sc_hd__mux2_1 _41246_ (.A0(_01341_),
    .A1(\decoded_imm[18] ),
    .S(_01304_),
    .X(_01342_));
 sky130_fd_sc_hd__mux2_1 _41247_ (.A0(_01342_),
    .A1(\cpuregs_rs1[18] ),
    .S(\cpu_state[3] ),
    .X(_02452_));
 sky130_fd_sc_hd__mux2_1 _41248_ (.A0(_01339_),
    .A1(\decoded_imm[17] ),
    .S(_01304_),
    .X(_01340_));
 sky130_fd_sc_hd__mux2_1 _41249_ (.A0(_01340_),
    .A1(\cpuregs_rs1[17] ),
    .S(\cpu_state[3] ),
    .X(_02451_));
 sky130_fd_sc_hd__mux2_1 _41250_ (.A0(_01337_),
    .A1(\decoded_imm[16] ),
    .S(_01304_),
    .X(_01338_));
 sky130_fd_sc_hd__mux2_1 _41251_ (.A0(_01338_),
    .A1(\cpuregs_rs1[16] ),
    .S(\cpu_state[3] ),
    .X(_02450_));
 sky130_fd_sc_hd__mux2_1 _41252_ (.A0(_01335_),
    .A1(\decoded_imm[15] ),
    .S(_01304_),
    .X(_01336_));
 sky130_fd_sc_hd__mux2_1 _41253_ (.A0(_01336_),
    .A1(\cpuregs_rs1[15] ),
    .S(\cpu_state[3] ),
    .X(_02449_));
 sky130_fd_sc_hd__mux2_1 _41254_ (.A0(_01333_),
    .A1(\decoded_imm[14] ),
    .S(_01304_),
    .X(_01334_));
 sky130_fd_sc_hd__mux2_1 _41255_ (.A0(_01334_),
    .A1(\cpuregs_rs1[14] ),
    .S(\cpu_state[3] ),
    .X(_02448_));
 sky130_fd_sc_hd__mux2_1 _41256_ (.A0(_01331_),
    .A1(\decoded_imm[13] ),
    .S(_01304_),
    .X(_01332_));
 sky130_fd_sc_hd__mux2_1 _41257_ (.A0(_01332_),
    .A1(\cpuregs_rs1[13] ),
    .S(\cpu_state[3] ),
    .X(_02447_));
 sky130_fd_sc_hd__mux2_1 _41258_ (.A0(_01329_),
    .A1(\decoded_imm[12] ),
    .S(_01304_),
    .X(_01330_));
 sky130_fd_sc_hd__mux2_1 _41259_ (.A0(_01330_),
    .A1(\cpuregs_rs1[12] ),
    .S(\cpu_state[3] ),
    .X(_02446_));
 sky130_fd_sc_hd__mux2_1 _41260_ (.A0(_01327_),
    .A1(\decoded_imm[11] ),
    .S(_01304_),
    .X(_01328_));
 sky130_fd_sc_hd__mux2_1 _41261_ (.A0(_01328_),
    .A1(\cpuregs_rs1[11] ),
    .S(\cpu_state[3] ),
    .X(_02445_));
 sky130_fd_sc_hd__mux2_1 _41262_ (.A0(_01325_),
    .A1(\decoded_imm[10] ),
    .S(_01304_),
    .X(_01326_));
 sky130_fd_sc_hd__mux2_1 _41263_ (.A0(_01326_),
    .A1(\cpuregs_rs1[10] ),
    .S(\cpu_state[3] ),
    .X(_02444_));
 sky130_fd_sc_hd__mux2_1 _41264_ (.A0(_01323_),
    .A1(\decoded_imm[9] ),
    .S(_01304_),
    .X(_01324_));
 sky130_fd_sc_hd__mux2_1 _41265_ (.A0(_01324_),
    .A1(\cpuregs_rs1[9] ),
    .S(\cpu_state[3] ),
    .X(_02474_));
 sky130_fd_sc_hd__mux2_1 _41266_ (.A0(_01321_),
    .A1(\decoded_imm[8] ),
    .S(_01304_),
    .X(_01322_));
 sky130_fd_sc_hd__mux2_1 _41267_ (.A0(_01322_),
    .A1(\cpuregs_rs1[8] ),
    .S(\cpu_state[3] ),
    .X(_02473_));
 sky130_fd_sc_hd__mux2_1 _41268_ (.A0(_01319_),
    .A1(\decoded_imm[7] ),
    .S(_01304_),
    .X(_01320_));
 sky130_fd_sc_hd__mux2_1 _41269_ (.A0(_01320_),
    .A1(\cpuregs_rs1[7] ),
    .S(\cpu_state[3] ),
    .X(_02472_));
 sky130_fd_sc_hd__mux2_1 _41270_ (.A0(_01317_),
    .A1(\decoded_imm[6] ),
    .S(_01304_),
    .X(_01318_));
 sky130_fd_sc_hd__mux2_1 _41271_ (.A0(_01318_),
    .A1(\cpuregs_rs1[6] ),
    .S(\cpu_state[3] ),
    .X(_02471_));
 sky130_fd_sc_hd__mux2_1 _41272_ (.A0(_01315_),
    .A1(\decoded_imm[5] ),
    .S(_01304_),
    .X(_01316_));
 sky130_fd_sc_hd__mux2_1 _41273_ (.A0(_01316_),
    .A1(\cpuregs_rs1[5] ),
    .S(\cpu_state[3] ),
    .X(_02470_));
 sky130_fd_sc_hd__mux2_1 _41274_ (.A0(\decoded_imm[4] ),
    .A1(\decoded_imm_uj[4] ),
    .S(is_slli_srli_srai),
    .X(_01313_));
 sky130_fd_sc_hd__mux2_1 _41275_ (.A0(_01313_),
    .A1(\decoded_imm[4] ),
    .S(_01304_),
    .X(_01314_));
 sky130_fd_sc_hd__mux2_1 _41276_ (.A0(_01314_),
    .A1(\cpuregs_rs1[4] ),
    .S(\cpu_state[3] ),
    .X(_02469_));
 sky130_fd_sc_hd__mux2_1 _41277_ (.A0(\decoded_imm[3] ),
    .A1(\decoded_imm_uj[3] ),
    .S(is_slli_srli_srai),
    .X(_01311_));
 sky130_fd_sc_hd__mux2_1 _41278_ (.A0(_01311_),
    .A1(\decoded_imm[3] ),
    .S(_01304_),
    .X(_01312_));
 sky130_fd_sc_hd__mux2_1 _41279_ (.A0(_01312_),
    .A1(\cpuregs_rs1[3] ),
    .S(\cpu_state[3] ),
    .X(_02468_));
 sky130_fd_sc_hd__mux2_1 _41280_ (.A0(\decoded_imm[2] ),
    .A1(\decoded_imm_uj[2] ),
    .S(is_slli_srli_srai),
    .X(_01309_));
 sky130_fd_sc_hd__mux2_1 _41281_ (.A0(_01309_),
    .A1(\decoded_imm[2] ),
    .S(_01304_),
    .X(_01310_));
 sky130_fd_sc_hd__mux2_1 _41282_ (.A0(_01310_),
    .A1(\cpuregs_rs1[2] ),
    .S(\cpu_state[3] ),
    .X(_02465_));
 sky130_fd_sc_hd__mux2_1 _41283_ (.A0(\decoded_imm[1] ),
    .A1(\decoded_imm_uj[1] ),
    .S(is_slli_srli_srai),
    .X(_01307_));
 sky130_fd_sc_hd__mux2_1 _41284_ (.A0(_01307_),
    .A1(\decoded_imm[1] ),
    .S(_01304_),
    .X(_01308_));
 sky130_fd_sc_hd__mux2_1 _41285_ (.A0(_01308_),
    .A1(\cpuregs_rs1[1] ),
    .S(\cpu_state[3] ),
    .X(_02454_));
 sky130_fd_sc_hd__mux2_1 _41286_ (.A0(\decoded_imm[0] ),
    .A1(\decoded_imm_uj[11] ),
    .S(is_slli_srli_srai),
    .X(_01305_));
 sky130_fd_sc_hd__mux2_1 _41287_ (.A0(_01305_),
    .A1(\decoded_imm[0] ),
    .S(_01304_),
    .X(_01306_));
 sky130_fd_sc_hd__mux2_1 _41288_ (.A0(_01306_),
    .A1(\cpuregs_rs1[0] ),
    .S(\cpu_state[3] ),
    .X(_02443_));
 sky130_fd_sc_hd__mux2_1 _41289_ (.A0(_01302_),
    .A1(\cpuregs_rs1[31] ),
    .S(instr_timer),
    .X(_01303_));
 sky130_fd_sc_hd__mux2_1 _41290_ (.A0(_01302_),
    .A1(_01303_),
    .S(\cpu_state[2] ),
    .X(_02435_));
 sky130_fd_sc_hd__mux2_1 _41291_ (.A0(_01299_),
    .A1(\cpuregs_rs1[30] ),
    .S(instr_timer),
    .X(_01300_));
 sky130_fd_sc_hd__mux2_1 _41292_ (.A0(_01299_),
    .A1(_01300_),
    .S(\cpu_state[2] ),
    .X(_02434_));
 sky130_fd_sc_hd__mux2_1 _41293_ (.A0(_01296_),
    .A1(\cpuregs_rs1[29] ),
    .S(instr_timer),
    .X(_01297_));
 sky130_fd_sc_hd__mux2_1 _41294_ (.A0(_01296_),
    .A1(_01297_),
    .S(\cpu_state[2] ),
    .X(_02432_));
 sky130_fd_sc_hd__mux2_1 _41295_ (.A0(_01293_),
    .A1(\cpuregs_rs1[28] ),
    .S(instr_timer),
    .X(_01294_));
 sky130_fd_sc_hd__mux2_1 _41296_ (.A0(_01293_),
    .A1(_01294_),
    .S(\cpu_state[2] ),
    .X(_02431_));
 sky130_fd_sc_hd__mux2_1 _41297_ (.A0(_01290_),
    .A1(\cpuregs_rs1[27] ),
    .S(instr_timer),
    .X(_01291_));
 sky130_fd_sc_hd__mux2_1 _41298_ (.A0(_01290_),
    .A1(_01291_),
    .S(\cpu_state[2] ),
    .X(_02430_));
 sky130_fd_sc_hd__mux2_1 _41299_ (.A0(_01287_),
    .A1(\cpuregs_rs1[26] ),
    .S(instr_timer),
    .X(_01288_));
 sky130_fd_sc_hd__mux2_1 _41300_ (.A0(_01287_),
    .A1(_01288_),
    .S(\cpu_state[2] ),
    .X(_02429_));
 sky130_fd_sc_hd__mux2_1 _41301_ (.A0(_01284_),
    .A1(\cpuregs_rs1[25] ),
    .S(instr_timer),
    .X(_01285_));
 sky130_fd_sc_hd__mux2_1 _41302_ (.A0(_01284_),
    .A1(_01285_),
    .S(\cpu_state[2] ),
    .X(_02428_));
 sky130_fd_sc_hd__mux2_1 _41303_ (.A0(_01281_),
    .A1(\cpuregs_rs1[24] ),
    .S(instr_timer),
    .X(_01282_));
 sky130_fd_sc_hd__mux2_1 _41304_ (.A0(_01281_),
    .A1(_01282_),
    .S(\cpu_state[2] ),
    .X(_02427_));
 sky130_fd_sc_hd__mux2_1 _41305_ (.A0(_01278_),
    .A1(\cpuregs_rs1[23] ),
    .S(instr_timer),
    .X(_01279_));
 sky130_fd_sc_hd__mux2_1 _41306_ (.A0(_01278_),
    .A1(_01279_),
    .S(\cpu_state[2] ),
    .X(_02426_));
 sky130_fd_sc_hd__mux2_1 _41307_ (.A0(_01275_),
    .A1(\cpuregs_rs1[22] ),
    .S(instr_timer),
    .X(_01276_));
 sky130_fd_sc_hd__mux2_1 _41308_ (.A0(_01275_),
    .A1(_01276_),
    .S(\cpu_state[2] ),
    .X(_02425_));
 sky130_fd_sc_hd__mux2_1 _41309_ (.A0(_01272_),
    .A1(\cpuregs_rs1[21] ),
    .S(instr_timer),
    .X(_01273_));
 sky130_fd_sc_hd__mux2_1 _41310_ (.A0(_01272_),
    .A1(_01273_),
    .S(\cpu_state[2] ),
    .X(_02424_));
 sky130_fd_sc_hd__mux2_1 _41311_ (.A0(_01269_),
    .A1(\cpuregs_rs1[20] ),
    .S(instr_timer),
    .X(_01270_));
 sky130_fd_sc_hd__mux2_1 _41312_ (.A0(_01269_),
    .A1(_01270_),
    .S(\cpu_state[2] ),
    .X(_02423_));
 sky130_fd_sc_hd__mux2_1 _41313_ (.A0(_01266_),
    .A1(\cpuregs_rs1[19] ),
    .S(instr_timer),
    .X(_01267_));
 sky130_fd_sc_hd__mux2_1 _41314_ (.A0(_01266_),
    .A1(_01267_),
    .S(\cpu_state[2] ),
    .X(_02421_));
 sky130_fd_sc_hd__mux2_1 _41315_ (.A0(_01263_),
    .A1(\cpuregs_rs1[18] ),
    .S(instr_timer),
    .X(_01264_));
 sky130_fd_sc_hd__mux2_1 _41316_ (.A0(_01263_),
    .A1(_01264_),
    .S(\cpu_state[2] ),
    .X(_02420_));
 sky130_fd_sc_hd__mux2_1 _41317_ (.A0(_01260_),
    .A1(\cpuregs_rs1[17] ),
    .S(instr_timer),
    .X(_01261_));
 sky130_fd_sc_hd__mux2_1 _41318_ (.A0(_01260_),
    .A1(_01261_),
    .S(\cpu_state[2] ),
    .X(_02419_));
 sky130_fd_sc_hd__mux2_1 _41319_ (.A0(_01257_),
    .A1(\cpuregs_rs1[16] ),
    .S(instr_timer),
    .X(_01258_));
 sky130_fd_sc_hd__mux2_1 _41320_ (.A0(_01257_),
    .A1(_01258_),
    .S(\cpu_state[2] ),
    .X(_02418_));
 sky130_fd_sc_hd__mux2_1 _41321_ (.A0(_01254_),
    .A1(\cpuregs_rs1[15] ),
    .S(instr_timer),
    .X(_01255_));
 sky130_fd_sc_hd__mux2_1 _41322_ (.A0(_01254_),
    .A1(_01255_),
    .S(\cpu_state[2] ),
    .X(_02417_));
 sky130_fd_sc_hd__mux2_1 _41323_ (.A0(_01251_),
    .A1(\cpuregs_rs1[14] ),
    .S(instr_timer),
    .X(_01252_));
 sky130_fd_sc_hd__mux2_1 _41324_ (.A0(_01251_),
    .A1(_01252_),
    .S(\cpu_state[2] ),
    .X(_02416_));
 sky130_fd_sc_hd__mux2_1 _41325_ (.A0(_01248_),
    .A1(\cpuregs_rs1[13] ),
    .S(instr_timer),
    .X(_01249_));
 sky130_fd_sc_hd__mux2_1 _41326_ (.A0(_01248_),
    .A1(_01249_),
    .S(\cpu_state[2] ),
    .X(_02415_));
 sky130_fd_sc_hd__mux2_1 _41327_ (.A0(_01245_),
    .A1(\cpuregs_rs1[12] ),
    .S(instr_timer),
    .X(_01246_));
 sky130_fd_sc_hd__mux2_1 _41328_ (.A0(_01245_),
    .A1(_01246_),
    .S(\cpu_state[2] ),
    .X(_02414_));
 sky130_fd_sc_hd__mux2_1 _41329_ (.A0(_01242_),
    .A1(\cpuregs_rs1[11] ),
    .S(instr_timer),
    .X(_01243_));
 sky130_fd_sc_hd__mux2_1 _41330_ (.A0(_01242_),
    .A1(_01243_),
    .S(\cpu_state[2] ),
    .X(_02413_));
 sky130_fd_sc_hd__mux2_1 _41331_ (.A0(_01239_),
    .A1(\cpuregs_rs1[10] ),
    .S(instr_timer),
    .X(_01240_));
 sky130_fd_sc_hd__mux2_1 _41332_ (.A0(_01239_),
    .A1(_01240_),
    .S(\cpu_state[2] ),
    .X(_02412_));
 sky130_fd_sc_hd__mux2_1 _41333_ (.A0(_01236_),
    .A1(\cpuregs_rs1[9] ),
    .S(instr_timer),
    .X(_01237_));
 sky130_fd_sc_hd__mux2_1 _41334_ (.A0(_01236_),
    .A1(_01237_),
    .S(\cpu_state[2] ),
    .X(_02442_));
 sky130_fd_sc_hd__mux2_1 _41335_ (.A0(_01233_),
    .A1(\cpuregs_rs1[8] ),
    .S(instr_timer),
    .X(_01234_));
 sky130_fd_sc_hd__mux2_1 _41336_ (.A0(_01233_),
    .A1(_01234_),
    .S(\cpu_state[2] ),
    .X(_02441_));
 sky130_fd_sc_hd__mux2_1 _41337_ (.A0(_01230_),
    .A1(\cpuregs_rs1[7] ),
    .S(instr_timer),
    .X(_01231_));
 sky130_fd_sc_hd__mux2_1 _41338_ (.A0(_01230_),
    .A1(_01231_),
    .S(\cpu_state[2] ),
    .X(_02440_));
 sky130_fd_sc_hd__mux2_1 _41339_ (.A0(_01227_),
    .A1(\cpuregs_rs1[6] ),
    .S(instr_timer),
    .X(_01228_));
 sky130_fd_sc_hd__mux2_1 _41340_ (.A0(_01227_),
    .A1(_01228_),
    .S(\cpu_state[2] ),
    .X(_02439_));
 sky130_fd_sc_hd__mux2_1 _41341_ (.A0(_01224_),
    .A1(\cpuregs_rs1[5] ),
    .S(instr_timer),
    .X(_01225_));
 sky130_fd_sc_hd__mux2_1 _41342_ (.A0(_01224_),
    .A1(_01225_),
    .S(\cpu_state[2] ),
    .X(_02438_));
 sky130_fd_sc_hd__mux2_1 _41343_ (.A0(_01221_),
    .A1(\cpuregs_rs1[4] ),
    .S(instr_timer),
    .X(_01222_));
 sky130_fd_sc_hd__mux2_1 _41344_ (.A0(_01221_),
    .A1(_01222_),
    .S(\cpu_state[2] ),
    .X(_02437_));
 sky130_fd_sc_hd__mux2_1 _41345_ (.A0(_01218_),
    .A1(\cpuregs_rs1[3] ),
    .S(instr_timer),
    .X(_01219_));
 sky130_fd_sc_hd__mux2_1 _41346_ (.A0(_01218_),
    .A1(_01219_),
    .S(\cpu_state[2] ),
    .X(_02436_));
 sky130_fd_sc_hd__mux2_1 _41347_ (.A0(_01215_),
    .A1(\cpuregs_rs1[2] ),
    .S(instr_timer),
    .X(_01216_));
 sky130_fd_sc_hd__mux2_1 _41348_ (.A0(_01215_),
    .A1(_01216_),
    .S(\cpu_state[2] ),
    .X(_02433_));
 sky130_fd_sc_hd__mux2_1 _41349_ (.A0(_01212_),
    .A1(\cpuregs_rs1[1] ),
    .S(instr_timer),
    .X(_01213_));
 sky130_fd_sc_hd__mux2_1 _41350_ (.A0(_01212_),
    .A1(_01213_),
    .S(\cpu_state[2] ),
    .X(_02422_));
 sky130_fd_sc_hd__mux2_1 _41351_ (.A0(_01209_),
    .A1(\cpuregs_rs1[0] ),
    .S(instr_timer),
    .X(_01210_));
 sky130_fd_sc_hd__mux2_1 _41352_ (.A0(_01209_),
    .A1(_01210_),
    .S(\cpu_state[2] ),
    .X(_02411_));
 sky130_fd_sc_hd__mux4_1 _41353_ (.A0(_01202_),
    .A1(_01203_),
    .A2(_01204_),
    .A3(_01205_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01206_));
 sky130_fd_sc_hd__mux4_1 _41354_ (.A0(_01181_),
    .A1(_01182_),
    .A2(_01183_),
    .A3(_01184_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01185_));
 sky130_fd_sc_hd__mux4_1 _41355_ (.A0(_01186_),
    .A1(_01187_),
    .A2(_01188_),
    .A3(_01189_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01190_));
 sky130_fd_sc_hd__mux4_1 _41356_ (.A0(_01191_),
    .A1(_01192_),
    .A2(_01193_),
    .A3(_01194_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01195_));
 sky130_fd_sc_hd__mux4_1 _41357_ (.A0(_01196_),
    .A1(_01197_),
    .A2(_01198_),
    .A3(_01199_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01200_));
 sky130_fd_sc_hd__mux4_1 _41358_ (.A0(_01185_),
    .A1(_01190_),
    .A2(_01195_),
    .A3(_01200_),
    .S0(_00360_),
    .S1(_00362_),
    .X(_01201_));
 sky130_fd_sc_hd__mux4_1 _41359_ (.A0(_01175_),
    .A1(_01176_),
    .A2(_01177_),
    .A3(_01178_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01179_));
 sky130_fd_sc_hd__mux4_1 _41360_ (.A0(_01154_),
    .A1(_01155_),
    .A2(_01156_),
    .A3(_01157_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01158_));
 sky130_fd_sc_hd__mux4_1 _41361_ (.A0(_01159_),
    .A1(_01160_),
    .A2(_01161_),
    .A3(_01162_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01163_));
 sky130_fd_sc_hd__mux4_1 _41362_ (.A0(_01164_),
    .A1(_01165_),
    .A2(_01166_),
    .A3(_01167_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01168_));
 sky130_fd_sc_hd__mux4_1 _41363_ (.A0(_01169_),
    .A1(_01170_),
    .A2(_01171_),
    .A3(_01172_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01173_));
 sky130_fd_sc_hd__mux4_1 _41364_ (.A0(_01158_),
    .A1(_01163_),
    .A2(_01168_),
    .A3(_01173_),
    .S0(_00360_),
    .S1(_00362_),
    .X(_01174_));
 sky130_fd_sc_hd__mux4_1 _41365_ (.A0(_01148_),
    .A1(_01149_),
    .A2(_01150_),
    .A3(_01151_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01152_));
 sky130_fd_sc_hd__mux4_1 _41366_ (.A0(_01127_),
    .A1(_01128_),
    .A2(_01129_),
    .A3(_01130_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01131_));
 sky130_fd_sc_hd__mux4_1 _41367_ (.A0(_01132_),
    .A1(_01133_),
    .A2(_01134_),
    .A3(_01135_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01136_));
 sky130_fd_sc_hd__mux4_1 _41368_ (.A0(_01137_),
    .A1(_01138_),
    .A2(_01139_),
    .A3(_01140_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01141_));
 sky130_fd_sc_hd__mux4_1 _41369_ (.A0(_01142_),
    .A1(_01143_),
    .A2(_01144_),
    .A3(_01145_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01146_));
 sky130_fd_sc_hd__mux4_1 _41370_ (.A0(_01131_),
    .A1(_01136_),
    .A2(_01141_),
    .A3(_01146_),
    .S0(_00360_),
    .S1(_00362_),
    .X(_01147_));
 sky130_fd_sc_hd__mux4_1 _41371_ (.A0(_01121_),
    .A1(_01122_),
    .A2(_01123_),
    .A3(_01124_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01125_));
 sky130_fd_sc_hd__mux4_1 _41372_ (.A0(_01100_),
    .A1(_01101_),
    .A2(_01102_),
    .A3(_01103_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01104_));
 sky130_fd_sc_hd__mux4_1 _41373_ (.A0(_01105_),
    .A1(_01106_),
    .A2(_01107_),
    .A3(_01108_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01109_));
 sky130_fd_sc_hd__mux4_1 _41374_ (.A0(_01110_),
    .A1(_01111_),
    .A2(_01112_),
    .A3(_01113_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01114_));
 sky130_fd_sc_hd__mux4_1 _41375_ (.A0(_01115_),
    .A1(_01116_),
    .A2(_01117_),
    .A3(_01118_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01119_));
 sky130_fd_sc_hd__mux4_1 _41376_ (.A0(_01104_),
    .A1(_01109_),
    .A2(_01114_),
    .A3(_01119_),
    .S0(_00360_),
    .S1(_00362_),
    .X(_01120_));
 sky130_fd_sc_hd__mux4_1 _41377_ (.A0(_01094_),
    .A1(_01095_),
    .A2(_01096_),
    .A3(_01097_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01098_));
 sky130_fd_sc_hd__mux4_1 _41378_ (.A0(_01073_),
    .A1(_01074_),
    .A2(_01075_),
    .A3(_01076_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01077_));
 sky130_fd_sc_hd__mux4_1 _41379_ (.A0(_01078_),
    .A1(_01079_),
    .A2(_01080_),
    .A3(_01081_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01082_));
 sky130_fd_sc_hd__mux4_1 _41380_ (.A0(_01083_),
    .A1(_01084_),
    .A2(_01085_),
    .A3(_01086_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01087_));
 sky130_fd_sc_hd__mux4_1 _41381_ (.A0(_01088_),
    .A1(_01089_),
    .A2(_01090_),
    .A3(_01091_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01092_));
 sky130_fd_sc_hd__mux4_1 _41382_ (.A0(_01077_),
    .A1(_01082_),
    .A2(_01087_),
    .A3(_01092_),
    .S0(_00360_),
    .S1(_00362_),
    .X(_01093_));
 sky130_fd_sc_hd__mux4_1 _41383_ (.A0(_01067_),
    .A1(_01068_),
    .A2(_01069_),
    .A3(_01070_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01071_));
 sky130_fd_sc_hd__mux4_1 _41384_ (.A0(_01046_),
    .A1(_01047_),
    .A2(_01048_),
    .A3(_01049_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01050_));
 sky130_fd_sc_hd__mux4_1 _41385_ (.A0(_01051_),
    .A1(_01052_),
    .A2(_01053_),
    .A3(_01054_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01055_));
 sky130_fd_sc_hd__mux4_1 _41386_ (.A0(_01056_),
    .A1(_01057_),
    .A2(_01058_),
    .A3(_01059_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01060_));
 sky130_fd_sc_hd__mux4_1 _41387_ (.A0(_01061_),
    .A1(_01062_),
    .A2(_01063_),
    .A3(_01064_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01065_));
 sky130_fd_sc_hd__mux4_1 _41388_ (.A0(_01050_),
    .A1(_01055_),
    .A2(_01060_),
    .A3(_01065_),
    .S0(_00360_),
    .S1(_00362_),
    .X(_01066_));
 sky130_fd_sc_hd__mux4_1 _41389_ (.A0(_01040_),
    .A1(_01041_),
    .A2(_01042_),
    .A3(_01043_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01044_));
 sky130_fd_sc_hd__mux4_1 _41390_ (.A0(_01019_),
    .A1(_01020_),
    .A2(_01021_),
    .A3(_01022_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01023_));
 sky130_fd_sc_hd__mux4_1 _41391_ (.A0(_01024_),
    .A1(_01025_),
    .A2(_01026_),
    .A3(_01027_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01028_));
 sky130_fd_sc_hd__mux4_1 _41392_ (.A0(_01029_),
    .A1(_01030_),
    .A2(_01031_),
    .A3(_01032_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01033_));
 sky130_fd_sc_hd__mux4_1 _41393_ (.A0(_01034_),
    .A1(_01035_),
    .A2(_01036_),
    .A3(_01037_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01038_));
 sky130_fd_sc_hd__mux4_1 _41394_ (.A0(_01023_),
    .A1(_01028_),
    .A2(_01033_),
    .A3(_01038_),
    .S0(_00360_),
    .S1(_00362_),
    .X(_01039_));
 sky130_fd_sc_hd__mux4_1 _41395_ (.A0(_01013_),
    .A1(_01014_),
    .A2(_01015_),
    .A3(_01016_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01017_));
 sky130_fd_sc_hd__mux4_1 _41396_ (.A0(_00992_),
    .A1(_00993_),
    .A2(_00994_),
    .A3(_00995_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00996_));
 sky130_fd_sc_hd__mux4_1 _41397_ (.A0(_00997_),
    .A1(_00998_),
    .A2(_00999_),
    .A3(_01000_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01001_));
 sky130_fd_sc_hd__mux4_1 _41398_ (.A0(_01002_),
    .A1(_01003_),
    .A2(_01004_),
    .A3(_01005_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01006_));
 sky130_fd_sc_hd__mux4_1 _41399_ (.A0(_01007_),
    .A1(_01008_),
    .A2(_01009_),
    .A3(_01010_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01011_));
 sky130_fd_sc_hd__mux4_1 _41400_ (.A0(_00996_),
    .A1(_01001_),
    .A2(_01006_),
    .A3(_01011_),
    .S0(_00360_),
    .S1(_00362_),
    .X(_01012_));
 sky130_fd_sc_hd__mux4_1 _41401_ (.A0(_00986_),
    .A1(_00987_),
    .A2(_00988_),
    .A3(_00989_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00990_));
 sky130_fd_sc_hd__mux4_1 _41402_ (.A0(_00965_),
    .A1(_00966_),
    .A2(_00967_),
    .A3(_00968_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00969_));
 sky130_fd_sc_hd__mux4_1 _41403_ (.A0(_00970_),
    .A1(_00971_),
    .A2(_00972_),
    .A3(_00973_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00974_));
 sky130_fd_sc_hd__mux4_1 _41404_ (.A0(_00975_),
    .A1(_00976_),
    .A2(_00977_),
    .A3(_00978_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00979_));
 sky130_fd_sc_hd__mux4_1 _41405_ (.A0(_00980_),
    .A1(_00981_),
    .A2(_00982_),
    .A3(_00983_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00984_));
 sky130_fd_sc_hd__mux4_1 _41406_ (.A0(_00969_),
    .A1(_00974_),
    .A2(_00979_),
    .A3(_00984_),
    .S0(_00360_),
    .S1(_00362_),
    .X(_00985_));
 sky130_fd_sc_hd__mux4_1 _41407_ (.A0(_00959_),
    .A1(_00960_),
    .A2(_00961_),
    .A3(_00962_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00963_));
 sky130_fd_sc_hd__mux4_1 _41408_ (.A0(_00938_),
    .A1(_00939_),
    .A2(_00940_),
    .A3(_00941_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00942_));
 sky130_fd_sc_hd__mux4_1 _41409_ (.A0(_00943_),
    .A1(_00944_),
    .A2(_00945_),
    .A3(_00946_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00947_));
 sky130_fd_sc_hd__mux4_1 _41410_ (.A0(_00948_),
    .A1(_00949_),
    .A2(_00950_),
    .A3(_00951_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00952_));
 sky130_fd_sc_hd__mux4_1 _41411_ (.A0(_00953_),
    .A1(_00954_),
    .A2(_00955_),
    .A3(_00956_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00957_));
 sky130_fd_sc_hd__mux4_1 _41412_ (.A0(_00942_),
    .A1(_00947_),
    .A2(_00952_),
    .A3(_00957_),
    .S0(_00360_),
    .S1(_00362_),
    .X(_00958_));
 sky130_fd_sc_hd__mux4_1 _41413_ (.A0(_00932_),
    .A1(_00933_),
    .A2(_00934_),
    .A3(_00935_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00936_));
 sky130_fd_sc_hd__mux4_1 _41414_ (.A0(_00911_),
    .A1(_00912_),
    .A2(_00913_),
    .A3(_00914_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00915_));
 sky130_fd_sc_hd__mux4_1 _41415_ (.A0(_00916_),
    .A1(_00917_),
    .A2(_00918_),
    .A3(_00919_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00920_));
 sky130_fd_sc_hd__mux4_1 _41416_ (.A0(_00921_),
    .A1(_00922_),
    .A2(_00923_),
    .A3(_00924_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00925_));
 sky130_fd_sc_hd__mux4_1 _41417_ (.A0(_00926_),
    .A1(_00927_),
    .A2(_00928_),
    .A3(_00929_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00930_));
 sky130_fd_sc_hd__mux4_1 _41418_ (.A0(_00915_),
    .A1(_00920_),
    .A2(_00925_),
    .A3(_00930_),
    .S0(_00360_),
    .S1(_00362_),
    .X(_00931_));
 sky130_fd_sc_hd__mux4_1 _41419_ (.A0(_00905_),
    .A1(_00906_),
    .A2(_00907_),
    .A3(_00908_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00909_));
 sky130_fd_sc_hd__mux4_1 _41420_ (.A0(_00884_),
    .A1(_00885_),
    .A2(_00886_),
    .A3(_00887_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00888_));
 sky130_fd_sc_hd__mux4_1 _41421_ (.A0(_00889_),
    .A1(_00890_),
    .A2(_00891_),
    .A3(_00892_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00893_));
 sky130_fd_sc_hd__mux4_1 _41422_ (.A0(_00894_),
    .A1(_00895_),
    .A2(_00896_),
    .A3(_00897_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00898_));
 sky130_fd_sc_hd__mux4_1 _41423_ (.A0(_00899_),
    .A1(_00900_),
    .A2(_00901_),
    .A3(_00902_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00903_));
 sky130_fd_sc_hd__mux4_1 _41424_ (.A0(_00888_),
    .A1(_00893_),
    .A2(_00898_),
    .A3(_00903_),
    .S0(_00360_),
    .S1(_00362_),
    .X(_00904_));
 sky130_fd_sc_hd__mux4_1 _41425_ (.A0(_00878_),
    .A1(_00879_),
    .A2(_00880_),
    .A3(_00881_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00882_));
 sky130_fd_sc_hd__mux4_1 _41426_ (.A0(_00857_),
    .A1(_00858_),
    .A2(_00859_),
    .A3(_00860_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00861_));
 sky130_fd_sc_hd__mux4_1 _41427_ (.A0(_00862_),
    .A1(_00863_),
    .A2(_00864_),
    .A3(_00865_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00866_));
 sky130_fd_sc_hd__mux4_1 _41428_ (.A0(_00867_),
    .A1(_00868_),
    .A2(_00869_),
    .A3(_00870_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00871_));
 sky130_fd_sc_hd__mux4_1 _41429_ (.A0(_00872_),
    .A1(_00873_),
    .A2(_00874_),
    .A3(_00875_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00876_));
 sky130_fd_sc_hd__mux4_1 _41430_ (.A0(_00861_),
    .A1(_00866_),
    .A2(_00871_),
    .A3(_00876_),
    .S0(_00360_),
    .S1(_00362_),
    .X(_00877_));
 sky130_fd_sc_hd__mux4_1 _41431_ (.A0(_00851_),
    .A1(_00852_),
    .A2(_00853_),
    .A3(_00854_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00855_));
 sky130_fd_sc_hd__mux4_1 _41432_ (.A0(_00830_),
    .A1(_00831_),
    .A2(_00832_),
    .A3(_00833_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00834_));
 sky130_fd_sc_hd__mux4_1 _41433_ (.A0(_00835_),
    .A1(_00836_),
    .A2(_00837_),
    .A3(_00838_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00839_));
 sky130_fd_sc_hd__mux4_1 _41434_ (.A0(_00840_),
    .A1(_00841_),
    .A2(_00842_),
    .A3(_00843_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00844_));
 sky130_fd_sc_hd__mux4_1 _41435_ (.A0(_00845_),
    .A1(_00846_),
    .A2(_00847_),
    .A3(_00848_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00849_));
 sky130_fd_sc_hd__mux4_1 _41436_ (.A0(_00834_),
    .A1(_00839_),
    .A2(_00844_),
    .A3(_00849_),
    .S0(_00360_),
    .S1(_00362_),
    .X(_00850_));
 sky130_fd_sc_hd__mux4_1 _41437_ (.A0(_00824_),
    .A1(_00825_),
    .A2(_00826_),
    .A3(_00827_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00828_));
 sky130_fd_sc_hd__mux4_1 _41438_ (.A0(_00803_),
    .A1(_00804_),
    .A2(_00805_),
    .A3(_00806_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00807_));
 sky130_fd_sc_hd__mux4_1 _41439_ (.A0(_00808_),
    .A1(_00809_),
    .A2(_00810_),
    .A3(_00811_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00812_));
 sky130_fd_sc_hd__mux4_1 _41440_ (.A0(_00813_),
    .A1(_00814_),
    .A2(_00815_),
    .A3(_00816_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00817_));
 sky130_fd_sc_hd__mux4_1 _41441_ (.A0(_00818_),
    .A1(_00819_),
    .A2(_00820_),
    .A3(_00821_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00822_));
 sky130_fd_sc_hd__mux4_1 _41442_ (.A0(_00807_),
    .A1(_00812_),
    .A2(_00817_),
    .A3(_00822_),
    .S0(_00360_),
    .S1(_00362_),
    .X(_00823_));
 sky130_fd_sc_hd__mux4_1 _41443_ (.A0(_00797_),
    .A1(_00798_),
    .A2(_00799_),
    .A3(_00800_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00801_));
 sky130_fd_sc_hd__mux4_1 _41444_ (.A0(_00776_),
    .A1(_00777_),
    .A2(_00778_),
    .A3(_00779_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00780_));
 sky130_fd_sc_hd__mux4_1 _41445_ (.A0(_00781_),
    .A1(_00782_),
    .A2(_00783_),
    .A3(_00784_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00785_));
 sky130_fd_sc_hd__mux4_1 _41446_ (.A0(_00786_),
    .A1(_00787_),
    .A2(_00788_),
    .A3(_00789_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00790_));
 sky130_fd_sc_hd__mux4_1 _41447_ (.A0(_00791_),
    .A1(_00792_),
    .A2(_00793_),
    .A3(_00794_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00795_));
 sky130_fd_sc_hd__mux4_1 _41448_ (.A0(_00780_),
    .A1(_00785_),
    .A2(_00790_),
    .A3(_00795_),
    .S0(_00360_),
    .S1(_00362_),
    .X(_00796_));
 sky130_fd_sc_hd__mux4_1 _41449_ (.A0(_00770_),
    .A1(_00771_),
    .A2(_00772_),
    .A3(_00773_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00774_));
 sky130_fd_sc_hd__mux4_1 _41450_ (.A0(_00749_),
    .A1(_00750_),
    .A2(_00751_),
    .A3(_00752_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00753_));
 sky130_fd_sc_hd__mux4_1 _41451_ (.A0(_00754_),
    .A1(_00755_),
    .A2(_00756_),
    .A3(_00757_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00758_));
 sky130_fd_sc_hd__mux4_1 _41452_ (.A0(_00759_),
    .A1(_00760_),
    .A2(_00761_),
    .A3(_00762_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00763_));
 sky130_fd_sc_hd__mux4_1 _41453_ (.A0(_00764_),
    .A1(_00765_),
    .A2(_00766_),
    .A3(_00767_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00768_));
 sky130_fd_sc_hd__mux4_1 _41454_ (.A0(_00753_),
    .A1(_00758_),
    .A2(_00763_),
    .A3(_00768_),
    .S0(_00360_),
    .S1(_00362_),
    .X(_00769_));
 sky130_fd_sc_hd__mux4_1 _41455_ (.A0(_00743_),
    .A1(_00744_),
    .A2(_00745_),
    .A3(_00746_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00747_));
 sky130_fd_sc_hd__mux4_1 _41456_ (.A0(_00722_),
    .A1(_00723_),
    .A2(_00724_),
    .A3(_00725_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00726_));
 sky130_fd_sc_hd__mux4_1 _41457_ (.A0(_00727_),
    .A1(_00728_),
    .A2(_00729_),
    .A3(_00730_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00731_));
 sky130_fd_sc_hd__mux4_1 _41458_ (.A0(_00732_),
    .A1(_00733_),
    .A2(_00734_),
    .A3(_00735_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00736_));
 sky130_fd_sc_hd__mux4_1 _41459_ (.A0(_00737_),
    .A1(_00738_),
    .A2(_00739_),
    .A3(_00740_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00741_));
 sky130_fd_sc_hd__mux4_1 _41460_ (.A0(_00726_),
    .A1(_00731_),
    .A2(_00736_),
    .A3(_00741_),
    .S0(_00360_),
    .S1(_00362_),
    .X(_00742_));
 sky130_fd_sc_hd__mux4_1 _41461_ (.A0(_00716_),
    .A1(_00717_),
    .A2(_00718_),
    .A3(_00719_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00720_));
 sky130_fd_sc_hd__mux4_1 _41462_ (.A0(_00695_),
    .A1(_00696_),
    .A2(_00697_),
    .A3(_00698_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00699_));
 sky130_fd_sc_hd__mux4_1 _41463_ (.A0(_00700_),
    .A1(_00701_),
    .A2(_00702_),
    .A3(_00703_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00704_));
 sky130_fd_sc_hd__mux4_1 _41464_ (.A0(_00705_),
    .A1(_00706_),
    .A2(_00707_),
    .A3(_00708_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00709_));
 sky130_fd_sc_hd__mux4_1 _41465_ (.A0(_00710_),
    .A1(_00711_),
    .A2(_00712_),
    .A3(_00713_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00714_));
 sky130_fd_sc_hd__mux4_1 _41466_ (.A0(_00699_),
    .A1(_00704_),
    .A2(_00709_),
    .A3(_00714_),
    .S0(_00360_),
    .S1(_00362_),
    .X(_00715_));
 sky130_fd_sc_hd__mux4_1 _41467_ (.A0(_00689_),
    .A1(_00690_),
    .A2(_00691_),
    .A3(_00692_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00693_));
 sky130_fd_sc_hd__mux4_1 _41468_ (.A0(_00668_),
    .A1(_00669_),
    .A2(_00670_),
    .A3(_00671_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00672_));
 sky130_fd_sc_hd__mux4_1 _41469_ (.A0(_00673_),
    .A1(_00674_),
    .A2(_00675_),
    .A3(_00676_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00677_));
 sky130_fd_sc_hd__mux4_1 _41470_ (.A0(_00678_),
    .A1(_00679_),
    .A2(_00680_),
    .A3(_00681_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00682_));
 sky130_fd_sc_hd__mux4_1 _41471_ (.A0(_00683_),
    .A1(_00684_),
    .A2(_00685_),
    .A3(_00686_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00687_));
 sky130_fd_sc_hd__mux4_1 _41472_ (.A0(_00672_),
    .A1(_00677_),
    .A2(_00682_),
    .A3(_00687_),
    .S0(_00360_),
    .S1(_00362_),
    .X(_00688_));
 sky130_fd_sc_hd__mux4_1 _41473_ (.A0(_00662_),
    .A1(_00663_),
    .A2(_00664_),
    .A3(_00665_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00666_));
 sky130_fd_sc_hd__mux4_1 _41474_ (.A0(_00641_),
    .A1(_00642_),
    .A2(_00643_),
    .A3(_00644_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00645_));
 sky130_fd_sc_hd__mux4_1 _41475_ (.A0(_00646_),
    .A1(_00647_),
    .A2(_00648_),
    .A3(_00649_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00650_));
 sky130_fd_sc_hd__mux4_1 _41476_ (.A0(_00651_),
    .A1(_00652_),
    .A2(_00653_),
    .A3(_00654_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00655_));
 sky130_fd_sc_hd__mux4_1 _41477_ (.A0(_00656_),
    .A1(_00657_),
    .A2(_00658_),
    .A3(_00659_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00660_));
 sky130_fd_sc_hd__mux4_1 _41478_ (.A0(_00645_),
    .A1(_00650_),
    .A2(_00655_),
    .A3(_00660_),
    .S0(_00360_),
    .S1(_00362_),
    .X(_00661_));
 sky130_fd_sc_hd__mux4_1 _41479_ (.A0(_00635_),
    .A1(_00636_),
    .A2(_00637_),
    .A3(_00638_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00639_));
 sky130_fd_sc_hd__mux4_1 _41480_ (.A0(_00614_),
    .A1(_00615_),
    .A2(_00616_),
    .A3(_00617_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00618_));
 sky130_fd_sc_hd__mux4_1 _41481_ (.A0(_00619_),
    .A1(_00620_),
    .A2(_00621_),
    .A3(_00622_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00623_));
 sky130_fd_sc_hd__mux4_1 _41482_ (.A0(_00624_),
    .A1(_00625_),
    .A2(_00626_),
    .A3(_00627_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00628_));
 sky130_fd_sc_hd__mux4_1 _41483_ (.A0(_00629_),
    .A1(_00630_),
    .A2(_00631_),
    .A3(_00632_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00633_));
 sky130_fd_sc_hd__mux4_1 _41484_ (.A0(_00618_),
    .A1(_00623_),
    .A2(_00628_),
    .A3(_00633_),
    .S0(_00360_),
    .S1(_00362_),
    .X(_00634_));
 sky130_fd_sc_hd__mux4_1 _41485_ (.A0(_00608_),
    .A1(_00609_),
    .A2(_00610_),
    .A3(_00611_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00612_));
 sky130_fd_sc_hd__mux4_1 _41486_ (.A0(_00587_),
    .A1(_00588_),
    .A2(_00589_),
    .A3(_00590_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00591_));
 sky130_fd_sc_hd__mux4_1 _41487_ (.A0(_00592_),
    .A1(_00593_),
    .A2(_00594_),
    .A3(_00595_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00596_));
 sky130_fd_sc_hd__mux4_1 _41488_ (.A0(_00597_),
    .A1(_00598_),
    .A2(_00599_),
    .A3(_00600_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00601_));
 sky130_fd_sc_hd__mux4_1 _41489_ (.A0(_00602_),
    .A1(_00603_),
    .A2(_00604_),
    .A3(_00605_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00606_));
 sky130_fd_sc_hd__mux4_1 _41490_ (.A0(_00591_),
    .A1(_00596_),
    .A2(_00601_),
    .A3(_00606_),
    .S0(_00360_),
    .S1(_00362_),
    .X(_00607_));
 sky130_fd_sc_hd__mux4_1 _41491_ (.A0(_00581_),
    .A1(_00582_),
    .A2(_00583_),
    .A3(_00584_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00585_));
 sky130_fd_sc_hd__mux4_1 _41492_ (.A0(_00560_),
    .A1(_00561_),
    .A2(_00562_),
    .A3(_00563_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00564_));
 sky130_fd_sc_hd__mux4_1 _41493_ (.A0(_00565_),
    .A1(_00566_),
    .A2(_00567_),
    .A3(_00568_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00569_));
 sky130_fd_sc_hd__mux4_1 _41494_ (.A0(_00570_),
    .A1(_00571_),
    .A2(_00572_),
    .A3(_00573_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00574_));
 sky130_fd_sc_hd__mux4_1 _41495_ (.A0(_00575_),
    .A1(_00576_),
    .A2(_00577_),
    .A3(_00578_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00579_));
 sky130_fd_sc_hd__mux4_1 _41496_ (.A0(_00564_),
    .A1(_00569_),
    .A2(_00574_),
    .A3(_00579_),
    .S0(_00360_),
    .S1(_00362_),
    .X(_00580_));
 sky130_fd_sc_hd__mux4_1 _41497_ (.A0(_00554_),
    .A1(_00555_),
    .A2(_00556_),
    .A3(_00557_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00558_));
 sky130_fd_sc_hd__mux4_1 _41498_ (.A0(_00533_),
    .A1(_00534_),
    .A2(_00535_),
    .A3(_00536_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00537_));
 sky130_fd_sc_hd__mux4_1 _41499_ (.A0(_00538_),
    .A1(_00539_),
    .A2(_00540_),
    .A3(_00541_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00542_));
 sky130_fd_sc_hd__mux4_1 _41500_ (.A0(_00543_),
    .A1(_00544_),
    .A2(_00545_),
    .A3(_00546_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00547_));
 sky130_fd_sc_hd__mux4_1 _41501_ (.A0(_00548_),
    .A1(_00549_),
    .A2(_00550_),
    .A3(_00551_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00552_));
 sky130_fd_sc_hd__mux4_1 _41502_ (.A0(_00537_),
    .A1(_00542_),
    .A2(_00547_),
    .A3(_00552_),
    .S0(_00360_),
    .S1(_00362_),
    .X(_00553_));
 sky130_fd_sc_hd__mux4_1 _41503_ (.A0(_00527_),
    .A1(_00528_),
    .A2(_00529_),
    .A3(_00530_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00531_));
 sky130_fd_sc_hd__mux4_1 _41504_ (.A0(_00506_),
    .A1(_00507_),
    .A2(_00508_),
    .A3(_00509_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00510_));
 sky130_fd_sc_hd__mux4_1 _41505_ (.A0(_00511_),
    .A1(_00512_),
    .A2(_00513_),
    .A3(_00514_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00515_));
 sky130_fd_sc_hd__mux4_1 _41506_ (.A0(_00516_),
    .A1(_00517_),
    .A2(_00518_),
    .A3(_00519_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00520_));
 sky130_fd_sc_hd__mux4_1 _41507_ (.A0(_00521_),
    .A1(_00522_),
    .A2(_00523_),
    .A3(_00524_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00525_));
 sky130_fd_sc_hd__mux4_1 _41508_ (.A0(_00510_),
    .A1(_00515_),
    .A2(_00520_),
    .A3(_00525_),
    .S0(_00360_),
    .S1(_00362_),
    .X(_00526_));
 sky130_fd_sc_hd__mux4_1 _41509_ (.A0(_00500_),
    .A1(_00501_),
    .A2(_00502_),
    .A3(_00503_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00504_));
 sky130_fd_sc_hd__mux4_1 _41510_ (.A0(_00479_),
    .A1(_00480_),
    .A2(_00481_),
    .A3(_00482_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00483_));
 sky130_fd_sc_hd__mux4_1 _41511_ (.A0(_00484_),
    .A1(_00485_),
    .A2(_00486_),
    .A3(_00487_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00488_));
 sky130_fd_sc_hd__mux4_1 _41512_ (.A0(_00489_),
    .A1(_00490_),
    .A2(_00491_),
    .A3(_00492_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00493_));
 sky130_fd_sc_hd__mux4_1 _41513_ (.A0(_00494_),
    .A1(_00495_),
    .A2(_00496_),
    .A3(_00497_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00498_));
 sky130_fd_sc_hd__mux4_1 _41514_ (.A0(_00483_),
    .A1(_00488_),
    .A2(_00493_),
    .A3(_00498_),
    .S0(_00360_),
    .S1(_00362_),
    .X(_00499_));
 sky130_fd_sc_hd__mux4_1 _41515_ (.A0(_00473_),
    .A1(_00474_),
    .A2(_00475_),
    .A3(_00476_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00477_));
 sky130_fd_sc_hd__mux4_1 _41516_ (.A0(_00452_),
    .A1(_00453_),
    .A2(_00454_),
    .A3(_00455_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00456_));
 sky130_fd_sc_hd__mux4_1 _41517_ (.A0(_00457_),
    .A1(_00458_),
    .A2(_00459_),
    .A3(_00460_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00461_));
 sky130_fd_sc_hd__mux4_1 _41518_ (.A0(_00462_),
    .A1(_00463_),
    .A2(_00464_),
    .A3(_00465_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00466_));
 sky130_fd_sc_hd__mux4_1 _41519_ (.A0(_00467_),
    .A1(_00468_),
    .A2(_00469_),
    .A3(_00470_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00471_));
 sky130_fd_sc_hd__mux4_1 _41520_ (.A0(_00456_),
    .A1(_00461_),
    .A2(_00466_),
    .A3(_00471_),
    .S0(_00360_),
    .S1(_00362_),
    .X(_00472_));
 sky130_fd_sc_hd__mux4_1 _41521_ (.A0(_00446_),
    .A1(_00447_),
    .A2(_00448_),
    .A3(_00449_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00450_));
 sky130_fd_sc_hd__mux4_1 _41522_ (.A0(_00425_),
    .A1(_00426_),
    .A2(_00427_),
    .A3(_00428_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00429_));
 sky130_fd_sc_hd__mux4_1 _41523_ (.A0(_00430_),
    .A1(_00431_),
    .A2(_00432_),
    .A3(_00433_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00434_));
 sky130_fd_sc_hd__mux4_1 _41524_ (.A0(_00435_),
    .A1(_00436_),
    .A2(_00437_),
    .A3(_00438_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00439_));
 sky130_fd_sc_hd__mux4_1 _41525_ (.A0(_00440_),
    .A1(_00441_),
    .A2(_00442_),
    .A3(_00443_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00444_));
 sky130_fd_sc_hd__mux4_1 _41526_ (.A0(_00429_),
    .A1(_00434_),
    .A2(_00439_),
    .A3(_00444_),
    .S0(_00360_),
    .S1(_00362_),
    .X(_00445_));
 sky130_fd_sc_hd__mux4_1 _41527_ (.A0(_00419_),
    .A1(_00420_),
    .A2(_00421_),
    .A3(_00422_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00423_));
 sky130_fd_sc_hd__mux4_1 _41528_ (.A0(_00398_),
    .A1(_00399_),
    .A2(_00400_),
    .A3(_00401_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00402_));
 sky130_fd_sc_hd__mux4_1 _41529_ (.A0(_00403_),
    .A1(_00404_),
    .A2(_00405_),
    .A3(_00406_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00407_));
 sky130_fd_sc_hd__mux4_1 _41530_ (.A0(_00408_),
    .A1(_00409_),
    .A2(_00410_),
    .A3(_00411_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00412_));
 sky130_fd_sc_hd__mux4_1 _41531_ (.A0(_00413_),
    .A1(_00414_),
    .A2(_00415_),
    .A3(_00416_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00417_));
 sky130_fd_sc_hd__mux4_1 _41532_ (.A0(_00402_),
    .A1(_00407_),
    .A2(_00412_),
    .A3(_00417_),
    .S0(_00360_),
    .S1(_00362_),
    .X(_00418_));
 sky130_fd_sc_hd__mux4_1 _41533_ (.A0(_00392_),
    .A1(_00393_),
    .A2(_00394_),
    .A3(_00395_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00396_));
 sky130_fd_sc_hd__mux4_1 _41534_ (.A0(_00371_),
    .A1(_00372_),
    .A2(_00373_),
    .A3(_00374_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00375_));
 sky130_fd_sc_hd__mux4_1 _41535_ (.A0(_00376_),
    .A1(_00377_),
    .A2(_00378_),
    .A3(_00379_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00380_));
 sky130_fd_sc_hd__mux4_1 _41536_ (.A0(_00381_),
    .A1(_00382_),
    .A2(_00383_),
    .A3(_00384_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00385_));
 sky130_fd_sc_hd__mux4_1 _41537_ (.A0(_00386_),
    .A1(_00387_),
    .A2(_00388_),
    .A3(_00389_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00390_));
 sky130_fd_sc_hd__mux4_1 _41538_ (.A0(_00375_),
    .A1(_00380_),
    .A2(_00385_),
    .A3(_00390_),
    .S0(_00360_),
    .S1(_00362_),
    .X(_00391_));
 sky130_fd_sc_hd__mux4_1 _41539_ (.A0(\cpuregs[16][0] ),
    .A1(\cpuregs[17][0] ),
    .A2(\cpuregs[18][0] ),
    .A3(\cpuregs[19][0] ),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00369_));
 sky130_fd_sc_hd__mux4_1 _41540_ (.A0(\cpuregs[0][0] ),
    .A1(\cpuregs[1][0] ),
    .A2(\cpuregs[2][0] ),
    .A3(\cpuregs[3][0] ),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00359_));
 sky130_fd_sc_hd__mux4_1 _41541_ (.A0(\cpuregs[4][0] ),
    .A1(\cpuregs[5][0] ),
    .A2(\cpuregs[6][0] ),
    .A3(\cpuregs[7][0] ),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00361_));
 sky130_fd_sc_hd__mux4_1 _41542_ (.A0(\cpuregs[8][0] ),
    .A1(\cpuregs[9][0] ),
    .A2(\cpuregs[10][0] ),
    .A3(\cpuregs[11][0] ),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00363_));
 sky130_fd_sc_hd__mux4_1 _41543_ (.A0(\cpuregs[12][0] ),
    .A1(\cpuregs[13][0] ),
    .A2(\cpuregs[14][0] ),
    .A3(\cpuregs[15][0] ),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00364_));
 sky130_fd_sc_hd__mux4_1 _41544_ (.A0(_00359_),
    .A1(_00361_),
    .A2(_00363_),
    .A3(_00364_),
    .S0(_00360_),
    .S1(_00362_),
    .X(_00365_));
 sky130_fd_sc_hd__mux4_1 _41545_ (.A0(_02581_),
    .A1(_01681_),
    .A2(_01679_),
    .A3(_02581_),
    .S0(_20586_),
    .S1(_00309_),
    .X(_01682_));
 sky130_fd_sc_hd__mux4_1 _41546_ (.A0(_02580_),
    .A1(_01677_),
    .A2(_01675_),
    .A3(_02580_),
    .S0(_20586_),
    .S1(_00309_),
    .X(_01678_));
 sky130_fd_sc_hd__mux4_1 _41547_ (.A0(_02579_),
    .A1(_01673_),
    .A2(_01671_),
    .A3(_02579_),
    .S0(_20586_),
    .S1(_00309_),
    .X(_01674_));
 sky130_fd_sc_hd__mux4_1 _41548_ (.A0(_02578_),
    .A1(_01669_),
    .A2(_01667_),
    .A3(_02578_),
    .S0(_20586_),
    .S1(_00309_),
    .X(_01670_));
 sky130_fd_sc_hd__mux4_1 _41549_ (.A0(_02577_),
    .A1(_01665_),
    .A2(_01663_),
    .A3(_02577_),
    .S0(_20586_),
    .S1(_00309_),
    .X(_01666_));
 sky130_fd_sc_hd__mux4_1 _41550_ (.A0(_02576_),
    .A1(_01661_),
    .A2(_01659_),
    .A3(_02576_),
    .S0(_20586_),
    .S1(_00309_),
    .X(_01662_));
 sky130_fd_sc_hd__mux4_1 _41551_ (.A0(_02575_),
    .A1(_01657_),
    .A2(_01655_),
    .A3(_02575_),
    .S0(_20586_),
    .S1(_00309_),
    .X(_01658_));
 sky130_fd_sc_hd__mux4_1 _41552_ (.A0(_02574_),
    .A1(_01653_),
    .A2(_01651_),
    .A3(_02574_),
    .S0(_20586_),
    .S1(_00309_),
    .X(_01654_));
 sky130_fd_sc_hd__mux4_1 _41553_ (.A0(_02573_),
    .A1(_01649_),
    .A2(_01647_),
    .A3(_02573_),
    .S0(_20586_),
    .S1(_00309_),
    .X(_01650_));
 sky130_fd_sc_hd__mux4_1 _41554_ (.A0(_02572_),
    .A1(_01645_),
    .A2(_01643_),
    .A3(_02572_),
    .S0(_20586_),
    .S1(_00309_),
    .X(_01646_));
 sky130_fd_sc_hd__mux4_1 _41555_ (.A0(_02570_),
    .A1(_01641_),
    .A2(_01639_),
    .A3(_02570_),
    .S0(_20586_),
    .S1(_00309_),
    .X(_01642_));
 sky130_fd_sc_hd__mux4_1 _41556_ (.A0(_02569_),
    .A1(_01637_),
    .A2(_01635_),
    .A3(_02569_),
    .S0(_20586_),
    .S1(_00309_),
    .X(_01638_));
 sky130_fd_sc_hd__mux4_1 _41557_ (.A0(_02568_),
    .A1(_01633_),
    .A2(_01631_),
    .A3(_02568_),
    .S0(_20586_),
    .S1(_00309_),
    .X(_01634_));
 sky130_fd_sc_hd__mux4_1 _41558_ (.A0(_02567_),
    .A1(_01629_),
    .A2(_01627_),
    .A3(_02567_),
    .S0(_20586_),
    .S1(_00309_),
    .X(_01630_));
 sky130_fd_sc_hd__mux4_1 _41559_ (.A0(_02566_),
    .A1(_01625_),
    .A2(_01623_),
    .A3(_02566_),
    .S0(_20586_),
    .S1(_00309_),
    .X(_01626_));
 sky130_fd_sc_hd__mux4_1 _41560_ (.A0(_02565_),
    .A1(_01621_),
    .A2(_01619_),
    .A3(_02565_),
    .S0(_20586_),
    .S1(_00309_),
    .X(_01622_));
 sky130_fd_sc_hd__mux4_1 _41561_ (.A0(_02564_),
    .A1(_01617_),
    .A2(_01615_),
    .A3(_02564_),
    .S0(_20586_),
    .S1(_00309_),
    .X(_01618_));
 sky130_fd_sc_hd__mux4_1 _41562_ (.A0(_02563_),
    .A1(_01613_),
    .A2(_01611_),
    .A3(_02563_),
    .S0(_20586_),
    .S1(_00309_),
    .X(_01614_));
 sky130_fd_sc_hd__mux4_1 _41563_ (.A0(_02562_),
    .A1(_01609_),
    .A2(_01607_),
    .A3(_02562_),
    .S0(_20586_),
    .S1(_00309_),
    .X(_01610_));
 sky130_fd_sc_hd__mux4_1 _41564_ (.A0(_02561_),
    .A1(_01605_),
    .A2(_01603_),
    .A3(_02561_),
    .S0(_20586_),
    .S1(_00309_),
    .X(_01606_));
 sky130_fd_sc_hd__mux4_1 _41565_ (.A0(_02589_),
    .A1(_01601_),
    .A2(_01599_),
    .A3(_02589_),
    .S0(_20586_),
    .S1(_00309_),
    .X(_01602_));
 sky130_fd_sc_hd__mux4_1 _41566_ (.A0(_02588_),
    .A1(_01597_),
    .A2(_01595_),
    .A3(_02588_),
    .S0(_20586_),
    .S1(_00309_),
    .X(_01598_));
 sky130_fd_sc_hd__mux4_1 _41567_ (.A0(_02587_),
    .A1(_01593_),
    .A2(_01591_),
    .A3(_02587_),
    .S0(_20586_),
    .S1(_00309_),
    .X(_01594_));
 sky130_fd_sc_hd__mux4_1 _41568_ (.A0(_02586_),
    .A1(_01589_),
    .A2(_01587_),
    .A3(_02586_),
    .S0(_20586_),
    .S1(_00309_),
    .X(_01590_));
 sky130_fd_sc_hd__mux4_1 _41569_ (.A0(_02585_),
    .A1(_01585_),
    .A2(_01583_),
    .A3(_02585_),
    .S0(_20586_),
    .S1(_00309_),
    .X(_01586_));
 sky130_fd_sc_hd__mux4_1 _41570_ (.A0(_02584_),
    .A1(_01581_),
    .A2(_01579_),
    .A3(_02584_),
    .S0(_20586_),
    .S1(_00309_),
    .X(_01582_));
 sky130_fd_sc_hd__mux4_1 _41571_ (.A0(_02583_),
    .A1(_01577_),
    .A2(_01575_),
    .A3(_02583_),
    .S0(_20586_),
    .S1(_00309_),
    .X(_01578_));
 sky130_fd_sc_hd__mux4_1 _41572_ (.A0(_02582_),
    .A1(_01573_),
    .A2(_01571_),
    .A3(_02582_),
    .S0(_20586_),
    .S1(_00309_),
    .X(_01574_));
 sky130_fd_sc_hd__mux4_1 _41573_ (.A0(_02571_),
    .A1(_01569_),
    .A2(_01567_),
    .A3(_02571_),
    .S0(_20586_),
    .S1(_00309_),
    .X(_01570_));
 sky130_fd_sc_hd__dfxtp_2 _41574_ (.D(_02687_),
    .Q(\alu_shl[0] ),
    .CLK(clknet_leaf_112_clk));
 sky130_fd_sc_hd__dfxtp_2 _41575_ (.D(_02688_),
    .Q(\alu_shl[1] ),
    .CLK(clknet_leaf_111_clk));
 sky130_fd_sc_hd__dfxtp_2 _41576_ (.D(_02689_),
    .Q(\alu_shl[2] ),
    .CLK(clknet_leaf_111_clk));
 sky130_fd_sc_hd__dfxtp_2 _41577_ (.D(_02690_),
    .Q(\alu_shl[3] ),
    .CLK(clknet_leaf_122_clk));
 sky130_fd_sc_hd__dfxtp_2 _41578_ (.D(_02691_),
    .Q(\alu_shl[4] ),
    .CLK(clknet_leaf_115_clk));
 sky130_fd_sc_hd__dfxtp_2 _41579_ (.D(_02692_),
    .Q(\alu_shl[5] ),
    .CLK(clknet_leaf_120_clk));
 sky130_fd_sc_hd__dfxtp_2 _41580_ (.D(_02693_),
    .Q(\alu_shl[6] ),
    .CLK(clknet_leaf_115_clk));
 sky130_fd_sc_hd__dfxtp_2 _41581_ (.D(_02694_),
    .Q(\alu_shl[7] ),
    .CLK(clknet_leaf_120_clk));
 sky130_fd_sc_hd__dfxtp_2 _41582_ (.D(_02695_),
    .Q(\alu_shl[8] ),
    .CLK(clknet_leaf_115_clk));
 sky130_fd_sc_hd__dfxtp_2 _41583_ (.D(_02696_),
    .Q(\alu_shl[9] ),
    .CLK(clknet_leaf_115_clk));
 sky130_fd_sc_hd__dfxtp_2 _41584_ (.D(_02697_),
    .Q(\alu_shl[10] ),
    .CLK(clknet_leaf_117_clk));
 sky130_fd_sc_hd__dfxtp_2 _41585_ (.D(_02698_),
    .Q(\alu_shl[11] ),
    .CLK(clknet_leaf_116_clk));
 sky130_fd_sc_hd__dfxtp_2 _41586_ (.D(_02699_),
    .Q(\alu_shl[12] ),
    .CLK(clknet_leaf_116_clk));
 sky130_fd_sc_hd__dfxtp_2 _41587_ (.D(_02700_),
    .Q(\alu_shl[13] ),
    .CLK(clknet_leaf_135_clk));
 sky130_fd_sc_hd__dfxtp_2 _41588_ (.D(_02701_),
    .Q(\alu_shl[14] ),
    .CLK(clknet_leaf_163_clk));
 sky130_fd_sc_hd__dfxtp_2 _41589_ (.D(_02702_),
    .Q(\alu_shl[15] ),
    .CLK(clknet_leaf_117_clk));
 sky130_fd_sc_hd__dfxtp_2 _41590_ (.D(_02703_),
    .Q(alu_wait),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__dfxtp_2 _41591_ (.D(_02704_),
    .Q(\latched_rd[3] ),
    .CLK(clknet_leaf_201_clk));
 sky130_fd_sc_hd__dfxtp_2 _41592_ (.D(_02705_),
    .Q(\latched_rd[2] ),
    .CLK(clknet_leaf_201_clk));
 sky130_fd_sc_hd__dfxtp_2 _41593_ (.D(_02706_),
    .Q(\latched_rd[1] ),
    .CLK(clknet_leaf_203_clk));
 sky130_fd_sc_hd__dfxtp_2 _41594_ (.D(_02707_),
    .Q(\latched_rd[0] ),
    .CLK(clknet_leaf_201_clk));
 sky130_fd_sc_hd__dfxtp_2 _41595_ (.D(_02708_),
    .Q(\decoded_imm[31] ),
    .CLK(clknet_leaf_214_clk));
 sky130_fd_sc_hd__dfxtp_2 _41596_ (.D(_02709_),
    .Q(\decoded_imm[30] ),
    .CLK(clknet_leaf_214_clk));
 sky130_fd_sc_hd__dfxtp_2 _41597_ (.D(_02710_),
    .Q(\decoded_imm[29] ),
    .CLK(clknet_leaf_202_clk));
 sky130_fd_sc_hd__dfxtp_2 _41598_ (.D(_02711_),
    .Q(\decoded_imm[28] ),
    .CLK(clknet_leaf_206_clk));
 sky130_fd_sc_hd__dfxtp_2 _41599_ (.D(_02712_),
    .Q(\decoded_imm[27] ),
    .CLK(clknet_leaf_202_clk));
 sky130_fd_sc_hd__dfxtp_2 _41600_ (.D(_02713_),
    .Q(\decoded_imm[26] ),
    .CLK(clknet_leaf_202_clk));
 sky130_fd_sc_hd__dfxtp_2 _41601_ (.D(_02714_),
    .Q(\decoded_imm[25] ),
    .CLK(clknet_leaf_206_clk));
 sky130_fd_sc_hd__dfxtp_2 _41602_ (.D(_02715_),
    .Q(\decoded_imm[24] ),
    .CLK(clknet_leaf_202_clk));
 sky130_fd_sc_hd__dfxtp_2 _41603_ (.D(_02716_),
    .Q(\decoded_imm[23] ),
    .CLK(clknet_leaf_202_clk));
 sky130_fd_sc_hd__dfxtp_2 _41604_ (.D(_02717_),
    .Q(\decoded_imm[22] ),
    .CLK(clknet_leaf_202_clk));
 sky130_fd_sc_hd__dfxtp_2 _41605_ (.D(_02718_),
    .Q(\decoded_imm[21] ),
    .CLK(clknet_leaf_205_clk));
 sky130_fd_sc_hd__dfxtp_2 _41606_ (.D(_02719_),
    .Q(\decoded_imm[20] ),
    .CLK(clknet_leaf_205_clk));
 sky130_fd_sc_hd__dfxtp_2 _41607_ (.D(_02720_),
    .Q(\decoded_imm[19] ),
    .CLK(clknet_leaf_215_clk));
 sky130_fd_sc_hd__dfxtp_2 _41608_ (.D(_02721_),
    .Q(\decoded_imm[18] ),
    .CLK(clknet_leaf_200_clk));
 sky130_fd_sc_hd__dfxtp_2 _41609_ (.D(_02722_),
    .Q(\decoded_imm[17] ),
    .CLK(clknet_leaf_230_clk));
 sky130_fd_sc_hd__dfxtp_2 _41610_ (.D(_02723_),
    .Q(\decoded_imm[16] ),
    .CLK(clknet_leaf_230_clk));
 sky130_fd_sc_hd__dfxtp_2 _41611_ (.D(_02724_),
    .Q(\decoded_imm[15] ),
    .CLK(clknet_leaf_186_clk));
 sky130_fd_sc_hd__dfxtp_2 _41612_ (.D(_02725_),
    .Q(\decoded_imm[14] ),
    .CLK(clknet_leaf_229_clk));
 sky130_fd_sc_hd__dfxtp_2 _41613_ (.D(_02726_),
    .Q(\decoded_imm[13] ),
    .CLK(clknet_leaf_186_clk));
 sky130_fd_sc_hd__dfxtp_2 _41614_ (.D(_02727_),
    .Q(\decoded_imm[12] ),
    .CLK(clknet_leaf_187_clk));
 sky130_fd_sc_hd__dfxtp_2 _41615_ (.D(_02728_),
    .Q(\decoded_imm[11] ),
    .CLK(clknet_leaf_201_clk));
 sky130_fd_sc_hd__dfxtp_2 _41616_ (.D(_02729_),
    .Q(\decoded_imm[10] ),
    .CLK(clknet_leaf_201_clk));
 sky130_fd_sc_hd__dfxtp_2 _41617_ (.D(_02730_),
    .Q(\decoded_imm[9] ),
    .CLK(clknet_leaf_215_clk));
 sky130_fd_sc_hd__dfxtp_2 _41618_ (.D(_02731_),
    .Q(\decoded_imm[8] ),
    .CLK(clknet_leaf_201_clk));
 sky130_fd_sc_hd__dfxtp_2 _41619_ (.D(_02732_),
    .Q(\decoded_imm[7] ),
    .CLK(clknet_leaf_201_clk));
 sky130_fd_sc_hd__dfxtp_2 _41620_ (.D(_02733_),
    .Q(\decoded_imm[6] ),
    .CLK(clknet_leaf_201_clk));
 sky130_fd_sc_hd__dfxtp_2 _41621_ (.D(_02734_),
    .Q(\decoded_imm[5] ),
    .CLK(clknet_leaf_214_clk));
 sky130_fd_sc_hd__dfxtp_2 _41622_ (.D(_02735_),
    .Q(\decoded_imm[4] ),
    .CLK(clknet_leaf_205_clk));
 sky130_fd_sc_hd__dfxtp_2 _41623_ (.D(_02736_),
    .Q(\decoded_imm[3] ),
    .CLK(clknet_leaf_205_clk));
 sky130_fd_sc_hd__dfxtp_2 _41624_ (.D(_02737_),
    .Q(\decoded_imm[2] ),
    .CLK(clknet_leaf_205_clk));
 sky130_fd_sc_hd__dfxtp_2 _41625_ (.D(_02738_),
    .Q(\decoded_imm[1] ),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__dfxtp_2 _41626_ (.D(_02739_),
    .Q(\irq_pending[31] ),
    .CLK(clknet_leaf_222_clk));
 sky130_fd_sc_hd__dfxtp_2 _41627_ (.D(_02740_),
    .Q(\irq_pending[30] ),
    .CLK(clknet_leaf_222_clk));
 sky130_fd_sc_hd__dfxtp_2 _41628_ (.D(_02741_),
    .Q(\irq_pending[29] ),
    .CLK(clknet_leaf_222_clk));
 sky130_fd_sc_hd__dfxtp_2 _41629_ (.D(_02742_),
    .Q(\irq_pending[28] ),
    .CLK(clknet_leaf_222_clk));
 sky130_fd_sc_hd__dfxtp_2 _41630_ (.D(_02743_),
    .Q(\irq_pending[27] ),
    .CLK(clknet_leaf_247_clk));
 sky130_fd_sc_hd__dfxtp_2 _41631_ (.D(_02744_),
    .Q(\irq_pending[26] ),
    .CLK(clknet_leaf_252_clk));
 sky130_fd_sc_hd__dfxtp_2 _41632_ (.D(_02745_),
    .Q(\irq_pending[25] ),
    .CLK(clknet_leaf_244_clk));
 sky130_fd_sc_hd__dfxtp_2 _41633_ (.D(_02746_),
    .Q(\irq_pending[24] ),
    .CLK(clknet_leaf_256_clk));
 sky130_fd_sc_hd__dfxtp_2 _41634_ (.D(_02747_),
    .Q(\irq_pending[23] ),
    .CLK(clknet_leaf_246_clk));
 sky130_fd_sc_hd__dfxtp_2 _41635_ (.D(_02748_),
    .Q(\irq_pending[22] ),
    .CLK(clknet_leaf_257_clk));
 sky130_fd_sc_hd__dfxtp_2 _41636_ (.D(_02749_),
    .Q(\irq_pending[21] ),
    .CLK(clknet_leaf_245_clk));
 sky130_fd_sc_hd__dfxtp_2 _41637_ (.D(_02750_),
    .Q(\irq_pending[20] ),
    .CLK(clknet_leaf_246_clk));
 sky130_fd_sc_hd__dfxtp_2 _41638_ (.D(_02751_),
    .Q(\irq_pending[19] ),
    .CLK(clknet_leaf_257_clk));
 sky130_fd_sc_hd__dfxtp_2 _41639_ (.D(_02752_),
    .Q(\irq_pending[18] ),
    .CLK(clknet_leaf_256_clk));
 sky130_fd_sc_hd__dfxtp_2 _41640_ (.D(_02753_),
    .Q(\irq_pending[17] ),
    .CLK(clknet_leaf_246_clk));
 sky130_fd_sc_hd__dfxtp_2 _41641_ (.D(_02754_),
    .Q(\irq_pending[16] ),
    .CLK(clknet_leaf_239_clk));
 sky130_fd_sc_hd__dfxtp_2 _41642_ (.D(_02755_),
    .Q(\irq_pending[15] ),
    .CLK(clknet_leaf_249_clk));
 sky130_fd_sc_hd__dfxtp_2 _41643_ (.D(_02756_),
    .Q(\irq_pending[14] ),
    .CLK(clknet_leaf_252_clk));
 sky130_fd_sc_hd__dfxtp_2 _41644_ (.D(_02757_),
    .Q(\irq_pending[13] ),
    .CLK(clknet_leaf_249_clk));
 sky130_fd_sc_hd__dfxtp_2 _41645_ (.D(_02758_),
    .Q(\irq_pending[12] ),
    .CLK(clknet_leaf_252_clk));
 sky130_fd_sc_hd__dfxtp_2 _41646_ (.D(_02759_),
    .Q(\irq_pending[11] ),
    .CLK(clknet_leaf_247_clk));
 sky130_fd_sc_hd__dfxtp_2 _41647_ (.D(_02760_),
    .Q(\irq_pending[10] ),
    .CLK(clknet_leaf_247_clk));
 sky130_fd_sc_hd__dfxtp_2 _41648_ (.D(_02761_),
    .Q(\irq_pending[9] ),
    .CLK(clknet_leaf_250_clk));
 sky130_fd_sc_hd__dfxtp_2 _41649_ (.D(_02762_),
    .Q(\irq_pending[8] ),
    .CLK(clknet_leaf_250_clk));
 sky130_fd_sc_hd__dfxtp_2 _41650_ (.D(_02763_),
    .Q(\irq_pending[7] ),
    .CLK(clknet_leaf_251_clk));
 sky130_fd_sc_hd__dfxtp_2 _41651_ (.D(_02764_),
    .Q(\irq_pending[6] ),
    .CLK(clknet_leaf_250_clk));
 sky130_fd_sc_hd__dfxtp_2 _41652_ (.D(_02765_),
    .Q(\irq_pending[5] ),
    .CLK(clknet_leaf_250_clk));
 sky130_fd_sc_hd__dfxtp_2 _41653_ (.D(_02766_),
    .Q(\irq_pending[4] ),
    .CLK(clknet_leaf_250_clk));
 sky130_fd_sc_hd__dfxtp_2 _41654_ (.D(_02767_),
    .Q(\irq_pending[3] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__dfxtp_2 _41655_ (.D(_02768_),
    .Q(\irq_pending[1] ),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfxtp_2 _41656_ (.D(_02769_),
    .Q(\irq_pending[0] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__dfxtp_2 _41657_ (.D(_02770_),
    .Q(\reg_next_pc[0] ),
    .CLK(clknet_leaf_224_clk));
 sky130_fd_sc_hd__dfxtp_2 _41658_ (.D(_00045_),
    .Q(\mem_wordsize[0] ),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__dfxtp_2 _41659_ (.D(_00046_),
    .Q(\mem_wordsize[1] ),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__dfxtp_2 _41660_ (.D(_00047_),
    .Q(\mem_wordsize[2] ),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__dfxtp_2 _41661_ (.D(_20588_),
    .Q(\reg_out[0] ),
    .CLK(clknet_leaf_221_clk));
 sky130_fd_sc_hd__dfxtp_2 _41662_ (.D(_20599_),
    .Q(\reg_out[1] ),
    .CLK(clknet_leaf_219_clk));
 sky130_fd_sc_hd__dfxtp_2 _41663_ (.D(_20610_),
    .Q(\reg_out[2] ),
    .CLK(clknet_5_30_0_clk));
 sky130_fd_sc_hd__dfxtp_2 _41664_ (.D(_20613_),
    .Q(\reg_out[3] ),
    .CLK(clknet_leaf_216_clk));
 sky130_fd_sc_hd__dfxtp_2 _41665_ (.D(_20614_),
    .Q(\reg_out[4] ),
    .CLK(clknet_leaf_216_clk));
 sky130_fd_sc_hd__dfxtp_2 _41666_ (.D(_20615_),
    .Q(\reg_out[5] ),
    .CLK(clknet_leaf_228_clk));
 sky130_fd_sc_hd__dfxtp_2 _41667_ (.D(_20616_),
    .Q(\reg_out[6] ),
    .CLK(clknet_leaf_224_clk));
 sky130_fd_sc_hd__dfxtp_2 _41668_ (.D(_20617_),
    .Q(\reg_out[7] ),
    .CLK(clknet_leaf_229_clk));
 sky130_fd_sc_hd__dfxtp_2 _41669_ (.D(_20618_),
    .Q(\reg_out[8] ),
    .CLK(clknet_leaf_230_clk));
 sky130_fd_sc_hd__dfxtp_2 _41670_ (.D(_20619_),
    .Q(\reg_out[9] ),
    .CLK(clknet_leaf_227_clk));
 sky130_fd_sc_hd__dfxtp_2 _41671_ (.D(_20589_),
    .Q(\reg_out[10] ),
    .CLK(clknet_leaf_225_clk));
 sky130_fd_sc_hd__dfxtp_2 _41672_ (.D(_20590_),
    .Q(\reg_out[11] ),
    .CLK(clknet_leaf_226_clk));
 sky130_fd_sc_hd__dfxtp_2 _41673_ (.D(_20591_),
    .Q(\reg_out[12] ),
    .CLK(clknet_leaf_230_clk));
 sky130_fd_sc_hd__dfxtp_2 _41674_ (.D(_20592_),
    .Q(\reg_out[13] ),
    .CLK(clknet_leaf_230_clk));
 sky130_fd_sc_hd__dfxtp_2 _41675_ (.D(_20593_),
    .Q(\reg_out[14] ),
    .CLK(clknet_leaf_231_clk));
 sky130_fd_sc_hd__dfxtp_2 _41676_ (.D(_20594_),
    .Q(\reg_out[15] ),
    .CLK(clknet_leaf_226_clk));
 sky130_fd_sc_hd__dfxtp_2 _41677_ (.D(_20595_),
    .Q(\reg_out[16] ),
    .CLK(clknet_leaf_231_clk));
 sky130_fd_sc_hd__dfxtp_2 _41678_ (.D(_20596_),
    .Q(\reg_out[17] ),
    .CLK(clknet_5_28_0_clk));
 sky130_fd_sc_hd__dfxtp_2 _41679_ (.D(_20597_),
    .Q(\reg_out[18] ),
    .CLK(clknet_leaf_231_clk));
 sky130_fd_sc_hd__dfxtp_2 _41680_ (.D(_20598_),
    .Q(\reg_out[19] ),
    .CLK(clknet_leaf_238_clk));
 sky130_fd_sc_hd__dfxtp_2 _41681_ (.D(_20600_),
    .Q(\reg_out[20] ),
    .CLK(clknet_leaf_233_clk));
 sky130_fd_sc_hd__dfxtp_2 _41682_ (.D(_20601_),
    .Q(\reg_out[21] ),
    .CLK(clknet_leaf_238_clk));
 sky130_fd_sc_hd__dfxtp_2 _41683_ (.D(_20602_),
    .Q(\reg_out[22] ),
    .CLK(clknet_leaf_234_clk));
 sky130_fd_sc_hd__dfxtp_2 _41684_ (.D(_20603_),
    .Q(\reg_out[23] ),
    .CLK(clknet_leaf_238_clk));
 sky130_fd_sc_hd__dfxtp_2 _41685_ (.D(_20604_),
    .Q(\reg_out[24] ),
    .CLK(clknet_leaf_234_clk));
 sky130_fd_sc_hd__dfxtp_2 _41686_ (.D(_20605_),
    .Q(\reg_out[25] ),
    .CLK(clknet_leaf_246_clk));
 sky130_fd_sc_hd__dfxtp_2 _41687_ (.D(_20606_),
    .Q(\reg_out[26] ),
    .CLK(clknet_leaf_225_clk));
 sky130_fd_sc_hd__dfxtp_2 _41688_ (.D(_20607_),
    .Q(\reg_out[27] ),
    .CLK(clknet_leaf_224_clk));
 sky130_fd_sc_hd__dfxtp_2 _41689_ (.D(_20608_),
    .Q(\reg_out[28] ),
    .CLK(clknet_leaf_247_clk));
 sky130_fd_sc_hd__dfxtp_2 _41690_ (.D(_20609_),
    .Q(\reg_out[29] ),
    .CLK(clknet_leaf_223_clk));
 sky130_fd_sc_hd__dfxtp_2 _41691_ (.D(_20611_),
    .Q(\reg_out[30] ),
    .CLK(clknet_leaf_224_clk));
 sky130_fd_sc_hd__dfxtp_2 _41692_ (.D(_20612_),
    .Q(\reg_out[31] ),
    .CLK(clknet_leaf_225_clk));
 sky130_fd_sc_hd__dfxtp_2 _41693_ (.D(_00004_),
    .Q(\irq_pending[2] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__dfxtp_2 _41694_ (.D(_00003_),
    .Q(decoder_trigger),
    .CLK(clknet_leaf_221_clk));
 sky130_fd_sc_hd__dfxtp_2 _41695_ (.D(\alu_out[0] ),
    .Q(\alu_out_q[0] ),
    .CLK(clknet_leaf_195_clk));
 sky130_fd_sc_hd__dfxtp_2 _41696_ (.D(\alu_out[1] ),
    .Q(\alu_out_q[1] ),
    .CLK(clknet_leaf_115_clk));
 sky130_fd_sc_hd__dfxtp_2 _41697_ (.D(\alu_out[2] ),
    .Q(\alu_out_q[2] ),
    .CLK(clknet_leaf_115_clk));
 sky130_fd_sc_hd__dfxtp_2 _41698_ (.D(\alu_out[3] ),
    .Q(\alu_out_q[3] ),
    .CLK(clknet_leaf_115_clk));
 sky130_fd_sc_hd__dfxtp_2 _41699_ (.D(\alu_out[4] ),
    .Q(\alu_out_q[4] ),
    .CLK(clknet_leaf_195_clk));
 sky130_fd_sc_hd__dfxtp_2 _41700_ (.D(\alu_out[5] ),
    .Q(\alu_out_q[5] ),
    .CLK(clknet_leaf_194_clk));
 sky130_fd_sc_hd__dfxtp_2 _41701_ (.D(\alu_out[6] ),
    .Q(\alu_out_q[6] ),
    .CLK(clknet_leaf_194_clk));
 sky130_fd_sc_hd__dfxtp_2 _41702_ (.D(\alu_out[7] ),
    .Q(\alu_out_q[7] ),
    .CLK(clknet_leaf_188_clk));
 sky130_fd_sc_hd__dfxtp_2 _41703_ (.D(\alu_out[8] ),
    .Q(\alu_out_q[8] ),
    .CLK(clknet_leaf_164_clk));
 sky130_fd_sc_hd__dfxtp_2 _41704_ (.D(\alu_out[9] ),
    .Q(\alu_out_q[9] ),
    .CLK(clknet_leaf_164_clk));
 sky130_fd_sc_hd__dfxtp_2 _41705_ (.D(\alu_out[10] ),
    .Q(\alu_out_q[10] ),
    .CLK(clknet_leaf_164_clk));
 sky130_fd_sc_hd__dfxtp_2 _41706_ (.D(\alu_out[11] ),
    .Q(\alu_out_q[11] ),
    .CLK(clknet_leaf_164_clk));
 sky130_fd_sc_hd__dfxtp_2 _41707_ (.D(\alu_out[12] ),
    .Q(\alu_out_q[12] ),
    .CLK(clknet_leaf_164_clk));
 sky130_fd_sc_hd__dfxtp_2 _41708_ (.D(\alu_out[13] ),
    .Q(\alu_out_q[13] ),
    .CLK(clknet_leaf_162_clk));
 sky130_fd_sc_hd__dfxtp_2 _41709_ (.D(\alu_out[14] ),
    .Q(\alu_out_q[14] ),
    .CLK(clknet_leaf_158_clk));
 sky130_fd_sc_hd__dfxtp_2 _41710_ (.D(\alu_out[15] ),
    .Q(\alu_out_q[15] ),
    .CLK(clknet_leaf_158_clk));
 sky130_fd_sc_hd__dfxtp_2 _41711_ (.D(\alu_out[16] ),
    .Q(\alu_out_q[16] ),
    .CLK(clknet_leaf_165_clk));
 sky130_fd_sc_hd__dfxtp_2 _41712_ (.D(\alu_out[17] ),
    .Q(\alu_out_q[17] ),
    .CLK(clknet_leaf_168_clk));
 sky130_fd_sc_hd__dfxtp_2 _41713_ (.D(\alu_out[18] ),
    .Q(\alu_out_q[18] ),
    .CLK(clknet_leaf_168_clk));
 sky130_fd_sc_hd__dfxtp_2 _41714_ (.D(\alu_out[19] ),
    .Q(\alu_out_q[19] ),
    .CLK(clknet_leaf_167_clk));
 sky130_fd_sc_hd__dfxtp_2 _41715_ (.D(\alu_out[20] ),
    .Q(\alu_out_q[20] ),
    .CLK(clknet_leaf_167_clk));
 sky130_fd_sc_hd__dfxtp_2 _41716_ (.D(\alu_out[21] ),
    .Q(\alu_out_q[21] ),
    .CLK(clknet_leaf_166_clk));
 sky130_fd_sc_hd__dfxtp_2 _41717_ (.D(\alu_out[22] ),
    .Q(\alu_out_q[22] ),
    .CLK(clknet_leaf_182_clk));
 sky130_fd_sc_hd__dfxtp_2 _41718_ (.D(\alu_out[23] ),
    .Q(\alu_out_q[23] ),
    .CLK(clknet_leaf_183_clk));
 sky130_fd_sc_hd__dfxtp_2 _41719_ (.D(\alu_out[24] ),
    .Q(\alu_out_q[24] ),
    .CLK(clknet_leaf_166_clk));
 sky130_fd_sc_hd__dfxtp_2 _41720_ (.D(\alu_out[25] ),
    .Q(\alu_out_q[25] ),
    .CLK(clknet_leaf_166_clk));
 sky130_fd_sc_hd__dfxtp_2 _41721_ (.D(\alu_out[26] ),
    .Q(\alu_out_q[26] ),
    .CLK(clknet_leaf_190_clk));
 sky130_fd_sc_hd__dfxtp_2 _41722_ (.D(\alu_out[27] ),
    .Q(\alu_out_q[27] ),
    .CLK(clknet_leaf_192_clk));
 sky130_fd_sc_hd__dfxtp_2 _41723_ (.D(\alu_out[28] ),
    .Q(\alu_out_q[28] ),
    .CLK(clknet_leaf_166_clk));
 sky130_fd_sc_hd__dfxtp_2 _41724_ (.D(\alu_out[29] ),
    .Q(\alu_out_q[29] ),
    .CLK(clknet_leaf_194_clk));
 sky130_fd_sc_hd__dfxtp_2 _41725_ (.D(\alu_out[30] ),
    .Q(\alu_out_q[30] ),
    .CLK(clknet_leaf_194_clk));
 sky130_fd_sc_hd__dfxtp_2 _41726_ (.D(\alu_out[31] ),
    .Q(\alu_out_q[31] ),
    .CLK(clknet_leaf_190_clk));
 sky130_fd_sc_hd__dfxtp_2 _41727_ (.D(_00005_),
    .Q(is_lui_auipc_jal),
    .CLK(clknet_leaf_201_clk));
 sky130_fd_sc_hd__dfxtp_2 _41728_ (.D(_00006_),
    .Q(is_slti_blt_slt),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__dfxtp_2 _41729_ (.D(_00007_),
    .Q(is_sltiu_bltu_sltu),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__dfxtp_2 _41730_ (.D(_02591_),
    .Q(\alu_add_sub[0] ),
    .CLK(clknet_5_15_0_clk));
 sky130_fd_sc_hd__dfxtp_2 _41731_ (.D(_02602_),
    .Q(\alu_add_sub[1] ),
    .CLK(clknet_leaf_111_clk));
 sky130_fd_sc_hd__dfxtp_2 _41732_ (.D(_02613_),
    .Q(\alu_add_sub[2] ),
    .CLK(clknet_leaf_111_clk));
 sky130_fd_sc_hd__dfxtp_2 _41733_ (.D(_02616_),
    .Q(\alu_add_sub[3] ),
    .CLK(clknet_leaf_111_clk));
 sky130_fd_sc_hd__dfxtp_2 _41734_ (.D(_02617_),
    .Q(\alu_add_sub[4] ),
    .CLK(clknet_leaf_112_clk));
 sky130_fd_sc_hd__dfxtp_2 _41735_ (.D(_02618_),
    .Q(\alu_add_sub[5] ),
    .CLK(clknet_leaf_112_clk));
 sky130_fd_sc_hd__dfxtp_2 _41736_ (.D(_02619_),
    .Q(\alu_add_sub[6] ),
    .CLK(clknet_leaf_196_clk));
 sky130_fd_sc_hd__dfxtp_2 _41737_ (.D(_02620_),
    .Q(\alu_add_sub[7] ),
    .CLK(clknet_leaf_196_clk));
 sky130_fd_sc_hd__dfxtp_2 _41738_ (.D(_02621_),
    .Q(\alu_add_sub[8] ),
    .CLK(clknet_leaf_116_clk));
 sky130_fd_sc_hd__dfxtp_2 _41739_ (.D(_02622_),
    .Q(\alu_add_sub[9] ),
    .CLK(clknet_leaf_116_clk));
 sky130_fd_sc_hd__dfxtp_2 _41740_ (.D(_02592_),
    .Q(\alu_add_sub[10] ),
    .CLK(clknet_leaf_117_clk));
 sky130_fd_sc_hd__dfxtp_2 _41741_ (.D(_02593_),
    .Q(\alu_add_sub[11] ),
    .CLK(clknet_5_9_0_clk));
 sky130_fd_sc_hd__dfxtp_2 _41742_ (.D(_02594_),
    .Q(\alu_add_sub[12] ),
    .CLK(clknet_leaf_163_clk));
 sky130_fd_sc_hd__dfxtp_2 _41743_ (.D(_02595_),
    .Q(\alu_add_sub[13] ),
    .CLK(clknet_leaf_164_clk));
 sky130_fd_sc_hd__dfxtp_2 _41744_ (.D(_02596_),
    .Q(\alu_add_sub[14] ),
    .CLK(clknet_leaf_162_clk));
 sky130_fd_sc_hd__dfxtp_2 _41745_ (.D(_02597_),
    .Q(\alu_add_sub[15] ),
    .CLK(clknet_leaf_162_clk));
 sky130_fd_sc_hd__dfxtp_2 _41746_ (.D(_02598_),
    .Q(\alu_add_sub[16] ),
    .CLK(clknet_leaf_165_clk));
 sky130_fd_sc_hd__dfxtp_2 _41747_ (.D(_02599_),
    .Q(\alu_add_sub[17] ),
    .CLK(clknet_leaf_168_clk));
 sky130_fd_sc_hd__dfxtp_2 _41748_ (.D(_02600_),
    .Q(\alu_add_sub[18] ),
    .CLK(clknet_leaf_168_clk));
 sky130_fd_sc_hd__dfxtp_2 _41749_ (.D(_02601_),
    .Q(\alu_add_sub[19] ),
    .CLK(clknet_leaf_167_clk));
 sky130_fd_sc_hd__dfxtp_2 _41750_ (.D(_02603_),
    .Q(\alu_add_sub[20] ),
    .CLK(clknet_leaf_167_clk));
 sky130_fd_sc_hd__dfxtp_2 _41751_ (.D(_02604_),
    .Q(\alu_add_sub[21] ),
    .CLK(clknet_leaf_166_clk));
 sky130_fd_sc_hd__dfxtp_2 _41752_ (.D(_02605_),
    .Q(\alu_add_sub[22] ),
    .CLK(clknet_leaf_166_clk));
 sky130_fd_sc_hd__dfxtp_2 _41753_ (.D(_02606_),
    .Q(\alu_add_sub[23] ),
    .CLK(clknet_leaf_166_clk));
 sky130_fd_sc_hd__dfxtp_2 _41754_ (.D(_02607_),
    .Q(\alu_add_sub[24] ),
    .CLK(clknet_leaf_191_clk));
 sky130_fd_sc_hd__dfxtp_2 _41755_ (.D(_02608_),
    .Q(\alu_add_sub[25] ),
    .CLK(clknet_leaf_191_clk));
 sky130_fd_sc_hd__dfxtp_2 _41756_ (.D(_02609_),
    .Q(\alu_add_sub[26] ),
    .CLK(clknet_leaf_192_clk));
 sky130_fd_sc_hd__dfxtp_2 _41757_ (.D(_02610_),
    .Q(\alu_add_sub[27] ),
    .CLK(clknet_leaf_192_clk));
 sky130_fd_sc_hd__dfxtp_2 _41758_ (.D(_02611_),
    .Q(\alu_add_sub[28] ),
    .CLK(clknet_leaf_194_clk));
 sky130_fd_sc_hd__dfxtp_2 _41759_ (.D(_02612_),
    .Q(\alu_add_sub[29] ),
    .CLK(clknet_leaf_194_clk));
 sky130_fd_sc_hd__dfxtp_2 _41760_ (.D(_02614_),
    .Q(\alu_add_sub[30] ),
    .CLK(clknet_leaf_195_clk));
 sky130_fd_sc_hd__dfxtp_2 _41761_ (.D(_02615_),
    .Q(\alu_add_sub[31] ),
    .CLK(clknet_leaf_195_clk));
 sky130_fd_sc_hd__dfxtp_2 _41762_ (.D(_20623_),
    .Q(\alu_shl[16] ),
    .CLK(clknet_leaf_115_clk));
 sky130_fd_sc_hd__dfxtp_2 _41763_ (.D(_20624_),
    .Q(\alu_shl[17] ),
    .CLK(clknet_leaf_122_clk));
 sky130_fd_sc_hd__dfxtp_2 _41764_ (.D(_20625_),
    .Q(\alu_shl[18] ),
    .CLK(clknet_leaf_163_clk));
 sky130_fd_sc_hd__dfxtp_2 _41765_ (.D(_20626_),
    .Q(\alu_shl[19] ),
    .CLK(clknet_leaf_121_clk));
 sky130_fd_sc_hd__dfxtp_2 _41766_ (.D(_20627_),
    .Q(\alu_shl[20] ),
    .CLK(clknet_leaf_116_clk));
 sky130_fd_sc_hd__dfxtp_2 _41767_ (.D(_20628_),
    .Q(\alu_shl[21] ),
    .CLK(clknet_leaf_120_clk));
 sky130_fd_sc_hd__dfxtp_2 _41768_ (.D(_20629_),
    .Q(\alu_shl[22] ),
    .CLK(clknet_leaf_163_clk));
 sky130_fd_sc_hd__dfxtp_2 _41769_ (.D(_20630_),
    .Q(\alu_shl[23] ),
    .CLK(clknet_leaf_136_clk));
 sky130_fd_sc_hd__dfxtp_2 _41770_ (.D(_20631_),
    .Q(\alu_shl[24] ),
    .CLK(clknet_leaf_115_clk));
 sky130_fd_sc_hd__dfxtp_2 _41771_ (.D(_20632_),
    .Q(\alu_shl[25] ),
    .CLK(clknet_leaf_118_clk));
 sky130_fd_sc_hd__dfxtp_2 _41772_ (.D(_20633_),
    .Q(\alu_shl[26] ),
    .CLK(clknet_5_14_0_clk));
 sky130_fd_sc_hd__dfxtp_2 _41773_ (.D(_20634_),
    .Q(\alu_shl[27] ),
    .CLK(clknet_leaf_120_clk));
 sky130_fd_sc_hd__dfxtp_2 _41774_ (.D(_20635_),
    .Q(\alu_shl[28] ),
    .CLK(clknet_leaf_116_clk));
 sky130_fd_sc_hd__dfxtp_2 _41775_ (.D(_20636_),
    .Q(\alu_shl[29] ),
    .CLK(clknet_leaf_118_clk));
 sky130_fd_sc_hd__dfxtp_2 _41776_ (.D(_20637_),
    .Q(\alu_shl[30] ),
    .CLK(clknet_leaf_117_clk));
 sky130_fd_sc_hd__dfxtp_2 _41777_ (.D(_20638_),
    .Q(\alu_shl[31] ),
    .CLK(clknet_leaf_118_clk));
 sky130_fd_sc_hd__dfxtp_2 _41778_ (.D(_20639_),
    .Q(\alu_shr[0] ),
    .CLK(clknet_leaf_136_clk));
 sky130_fd_sc_hd__dfxtp_2 _41779_ (.D(_20650_),
    .Q(\alu_shr[1] ),
    .CLK(clknet_leaf_118_clk));
 sky130_fd_sc_hd__dfxtp_2 _41780_ (.D(_20661_),
    .Q(\alu_shr[2] ),
    .CLK(clknet_leaf_162_clk));
 sky130_fd_sc_hd__dfxtp_2 _41781_ (.D(_20664_),
    .Q(\alu_shr[3] ),
    .CLK(clknet_leaf_118_clk));
 sky130_fd_sc_hd__dfxtp_2 _41782_ (.D(_20665_),
    .Q(\alu_shr[4] ),
    .CLK(clknet_leaf_163_clk));
 sky130_fd_sc_hd__dfxtp_2 _41783_ (.D(_20666_),
    .Q(\alu_shr[5] ),
    .CLK(clknet_leaf_117_clk));
 sky130_fd_sc_hd__dfxtp_2 _41784_ (.D(_20667_),
    .Q(\alu_shr[6] ),
    .CLK(clknet_leaf_163_clk));
 sky130_fd_sc_hd__dfxtp_2 _41785_ (.D(_20668_),
    .Q(\alu_shr[7] ),
    .CLK(clknet_leaf_117_clk));
 sky130_fd_sc_hd__dfxtp_2 _41786_ (.D(_20669_),
    .Q(\alu_shr[8] ),
    .CLK(clknet_leaf_135_clk));
 sky130_fd_sc_hd__dfxtp_2 _41787_ (.D(_20670_),
    .Q(\alu_shr[9] ),
    .CLK(clknet_5_9_0_clk));
 sky130_fd_sc_hd__dfxtp_2 _41788_ (.D(_20640_),
    .Q(\alu_shr[10] ),
    .CLK(clknet_leaf_162_clk));
 sky130_fd_sc_hd__dfxtp_2 _41789_ (.D(_20641_),
    .Q(\alu_shr[11] ),
    .CLK(clknet_leaf_117_clk));
 sky130_fd_sc_hd__dfxtp_2 _41790_ (.D(_20642_),
    .Q(\alu_shr[12] ),
    .CLK(clknet_leaf_135_clk));
 sky130_fd_sc_hd__dfxtp_2 _41791_ (.D(_20643_),
    .Q(\alu_shr[13] ),
    .CLK(clknet_leaf_163_clk));
 sky130_fd_sc_hd__dfxtp_2 _41792_ (.D(_20644_),
    .Q(\alu_shr[14] ),
    .CLK(clknet_leaf_163_clk));
 sky130_fd_sc_hd__dfxtp_2 _41793_ (.D(_20645_),
    .Q(\alu_shr[15] ),
    .CLK(clknet_leaf_117_clk));
 sky130_fd_sc_hd__dfxtp_2 _41794_ (.D(_20646_),
    .Q(\alu_shr[16] ),
    .CLK(clknet_leaf_163_clk));
 sky130_fd_sc_hd__dfxtp_2 _41795_ (.D(_20647_),
    .Q(\alu_shr[17] ),
    .CLK(clknet_leaf_135_clk));
 sky130_fd_sc_hd__dfxtp_2 _41796_ (.D(_20648_),
    .Q(\alu_shr[18] ),
    .CLK(clknet_leaf_162_clk));
 sky130_fd_sc_hd__dfxtp_2 _41797_ (.D(_20649_),
    .Q(\alu_shr[19] ),
    .CLK(clknet_leaf_135_clk));
 sky130_fd_sc_hd__dfxtp_2 _41798_ (.D(_20651_),
    .Q(\alu_shr[20] ),
    .CLK(clknet_leaf_163_clk));
 sky130_fd_sc_hd__dfxtp_2 _41799_ (.D(_20652_),
    .Q(\alu_shr[21] ),
    .CLK(clknet_leaf_162_clk));
 sky130_fd_sc_hd__dfxtp_2 _41800_ (.D(_20653_),
    .Q(\alu_shr[22] ),
    .CLK(clknet_leaf_162_clk));
 sky130_fd_sc_hd__dfxtp_2 _41801_ (.D(_20654_),
    .Q(\alu_shr[23] ),
    .CLK(clknet_leaf_135_clk));
 sky130_fd_sc_hd__dfxtp_2 _41802_ (.D(_20655_),
    .Q(\alu_shr[24] ),
    .CLK(clknet_leaf_135_clk));
 sky130_fd_sc_hd__dfxtp_2 _41803_ (.D(_20656_),
    .Q(\alu_shr[25] ),
    .CLK(clknet_leaf_135_clk));
 sky130_fd_sc_hd__dfxtp_2 _41804_ (.D(_20657_),
    .Q(\alu_shr[26] ),
    .CLK(clknet_leaf_162_clk));
 sky130_fd_sc_hd__dfxtp_2 _41805_ (.D(_20658_),
    .Q(\alu_shr[27] ),
    .CLK(clknet_leaf_135_clk));
 sky130_fd_sc_hd__dfxtp_2 _41806_ (.D(_20659_),
    .Q(\alu_shr[28] ),
    .CLK(clknet_leaf_163_clk));
 sky130_fd_sc_hd__dfxtp_2 _41807_ (.D(_20660_),
    .Q(\alu_shr[29] ),
    .CLK(clknet_leaf_117_clk));
 sky130_fd_sc_hd__dfxtp_2 _41808_ (.D(_20662_),
    .Q(\alu_shr[30] ),
    .CLK(clknet_leaf_163_clk));
 sky130_fd_sc_hd__dfxtp_2 _41809_ (.D(_20663_),
    .Q(\alu_shr[31] ),
    .CLK(clknet_leaf_117_clk));
 sky130_fd_sc_hd__dfxtp_2 _41810_ (.D(_00000_),
    .Q(alu_eq),
    .CLK(clknet_leaf_109_clk));
 sky130_fd_sc_hd__dfxtp_2 _41811_ (.D(_00002_),
    .Q(alu_ltu),
    .CLK(clknet_leaf_109_clk));
 sky130_fd_sc_hd__dfxtp_2 _41812_ (.D(_00001_),
    .Q(alu_lts),
    .CLK(clknet_leaf_109_clk));
 sky130_fd_sc_hd__dfxtp_2 _41813_ (.D(_02623_),
    .Q(\pcpi_mul.rd[0] ),
    .CLK(clknet_leaf_207_clk));
 sky130_fd_sc_hd__dfxtp_2 _41814_ (.D(_02624_),
    .Q(\pcpi_mul.rd[1] ),
    .CLK(clknet_leaf_208_clk));
 sky130_fd_sc_hd__dfxtp_2 _41815_ (.D(_02625_),
    .Q(\pcpi_mul.rd[2] ),
    .CLK(clknet_leaf_207_clk));
 sky130_fd_sc_hd__dfxtp_2 _41816_ (.D(_02626_),
    .Q(\pcpi_mul.rd[3] ),
    .CLK(clknet_leaf_207_clk));
 sky130_fd_sc_hd__dfxtp_2 _41817_ (.D(_02627_),
    .Q(\pcpi_mul.rd[4] ),
    .CLK(clknet_leaf_208_clk));
 sky130_fd_sc_hd__dfxtp_2 _41818_ (.D(_02628_),
    .Q(\pcpi_mul.rd[5] ),
    .CLK(clknet_leaf_208_clk));
 sky130_fd_sc_hd__dfxtp_2 _41819_ (.D(_02683_),
    .Q(\pcpi_mul.rd[6] ),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__dfxtp_2 _41820_ (.D(_02684_),
    .Q(\pcpi_mul.rd[7] ),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__dfxtp_2 _41821_ (.D(_02685_),
    .Q(\pcpi_mul.rd[8] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__dfxtp_2 _41822_ (.D(_02686_),
    .Q(\pcpi_mul.rd[9] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__dfxtp_2 _41823_ (.D(_02629_),
    .Q(\pcpi_mul.rd[10] ),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__dfxtp_2 _41824_ (.D(_02630_),
    .Q(\pcpi_mul.rd[11] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__dfxtp_2 _41825_ (.D(_02631_),
    .Q(\pcpi_mul.rd[12] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__dfxtp_2 _41826_ (.D(_02632_),
    .Q(\pcpi_mul.rd[13] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__dfxtp_2 _41827_ (.D(_02633_),
    .Q(\pcpi_mul.rd[14] ),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__dfxtp_2 _41828_ (.D(_02634_),
    .Q(\pcpi_mul.rd[15] ),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__dfxtp_2 _41829_ (.D(_02635_),
    .Q(\pcpi_mul.rd[16] ),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__dfxtp_2 _41830_ (.D(_02636_),
    .Q(\pcpi_mul.rd[17] ),
    .CLK(clknet_5_20_0_clk));
 sky130_fd_sc_hd__dfxtp_2 _41831_ (.D(_02637_),
    .Q(\pcpi_mul.rd[18] ),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__dfxtp_2 _41832_ (.D(_02638_),
    .Q(\pcpi_mul.rd[19] ),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__dfxtp_2 _41833_ (.D(_02639_),
    .Q(\pcpi_mul.rd[20] ),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__dfxtp_2 _41834_ (.D(_02640_),
    .Q(\pcpi_mul.rd[21] ),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__dfxtp_2 _41835_ (.D(_02641_),
    .Q(\pcpi_mul.rd[22] ),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__dfxtp_2 _41836_ (.D(_02642_),
    .Q(\pcpi_mul.rd[23] ),
    .CLK(clknet_5_21_0_clk));
 sky130_fd_sc_hd__dfxtp_2 _41837_ (.D(_02643_),
    .Q(\pcpi_mul.rd[24] ),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__dfxtp_2 _41838_ (.D(_02644_),
    .Q(\pcpi_mul.rd[25] ),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__dfxtp_2 _41839_ (.D(_02645_),
    .Q(\pcpi_mul.rd[26] ),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__dfxtp_2 _41840_ (.D(_02646_),
    .Q(\pcpi_mul.rd[27] ),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__dfxtp_2 _41841_ (.D(_02647_),
    .Q(\pcpi_mul.rd[28] ),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__dfxtp_2 _41842_ (.D(_02648_),
    .Q(\pcpi_mul.rd[29] ),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__dfxtp_2 _41843_ (.D(_02649_),
    .Q(\pcpi_mul.rd[30] ),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__dfxtp_2 _41844_ (.D(_02650_),
    .Q(\pcpi_mul.rd[31] ),
    .CLK(clknet_opt_27_clk));
 sky130_fd_sc_hd__dfxtp_2 _41845_ (.D(_02651_),
    .Q(\pcpi_mul.rd[32] ),
    .CLK(clknet_leaf_207_clk));
 sky130_fd_sc_hd__dfxtp_2 _41846_ (.D(_02652_),
    .Q(\pcpi_mul.rd[33] ),
    .CLK(clknet_leaf_207_clk));
 sky130_fd_sc_hd__dfxtp_2 _41847_ (.D(_02653_),
    .Q(\pcpi_mul.rd[34] ),
    .CLK(clknet_leaf_122_clk));
 sky130_fd_sc_hd__dfxtp_2 _41848_ (.D(_02654_),
    .Q(\pcpi_mul.rd[35] ),
    .CLK(clknet_leaf_122_clk));
 sky130_fd_sc_hd__dfxtp_2 _41849_ (.D(_02655_),
    .Q(\pcpi_mul.rd[36] ),
    .CLK(clknet_leaf_123_clk));
 sky130_fd_sc_hd__dfxtp_2 _41850_ (.D(_02656_),
    .Q(\pcpi_mul.rd[37] ),
    .CLK(clknet_leaf_123_clk));
 sky130_fd_sc_hd__dfxtp_2 _41851_ (.D(_02657_),
    .Q(\pcpi_mul.rd[38] ),
    .CLK(clknet_leaf_125_clk));
 sky130_fd_sc_hd__dfxtp_2 _41852_ (.D(_02658_),
    .Q(\pcpi_mul.rd[39] ),
    .CLK(clknet_leaf_125_clk));
 sky130_fd_sc_hd__dfxtp_2 _41853_ (.D(_02659_),
    .Q(\pcpi_mul.rd[40] ),
    .CLK(clknet_leaf_124_clk));
 sky130_fd_sc_hd__dfxtp_2 _41854_ (.D(_02660_),
    .Q(\pcpi_mul.rd[41] ),
    .CLK(clknet_leaf_124_clk));
 sky130_fd_sc_hd__dfxtp_2 _41855_ (.D(_02661_),
    .Q(\pcpi_mul.rd[42] ),
    .CLK(clknet_leaf_124_clk));
 sky130_fd_sc_hd__dfxtp_2 _41856_ (.D(_02662_),
    .Q(\pcpi_mul.rd[43] ),
    .CLK(clknet_leaf_124_clk));
 sky130_fd_sc_hd__dfxtp_2 _41857_ (.D(_02663_),
    .Q(\pcpi_mul.rd[44] ),
    .CLK(clknet_leaf_124_clk));
 sky130_fd_sc_hd__dfxtp_2 _41858_ (.D(_02664_),
    .Q(\pcpi_mul.rd[45] ),
    .CLK(clknet_leaf_124_clk));
 sky130_fd_sc_hd__dfxtp_2 _41859_ (.D(_02665_),
    .Q(\pcpi_mul.rd[46] ),
    .CLK(clknet_5_12_0_clk));
 sky130_fd_sc_hd__dfxtp_2 _41860_ (.D(_02666_),
    .Q(\pcpi_mul.rd[47] ),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__dfxtp_2 _41861_ (.D(_02667_),
    .Q(\pcpi_mul.rd[48] ),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__dfxtp_2 _41862_ (.D(_02668_),
    .Q(\pcpi_mul.rd[49] ),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__dfxtp_2 _41863_ (.D(_02669_),
    .Q(\pcpi_mul.rd[50] ),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__dfxtp_2 _41864_ (.D(_02670_),
    .Q(\pcpi_mul.rd[51] ),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__dfxtp_2 _41865_ (.D(_02671_),
    .Q(\pcpi_mul.rd[52] ),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__dfxtp_2 _41866_ (.D(_02672_),
    .Q(\pcpi_mul.rd[53] ),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__dfxtp_2 _41867_ (.D(_02673_),
    .Q(\pcpi_mul.rd[54] ),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__dfxtp_2 _41868_ (.D(_02674_),
    .Q(\pcpi_mul.rd[55] ),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__dfxtp_2 _41869_ (.D(_02675_),
    .Q(\pcpi_mul.rd[56] ),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__dfxtp_2 _41870_ (.D(_02676_),
    .Q(\pcpi_mul.rd[57] ),
    .CLK(clknet_opt_28_clk));
 sky130_fd_sc_hd__dfxtp_2 _41871_ (.D(_02677_),
    .Q(\pcpi_mul.rd[58] ),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__dfxtp_2 _41872_ (.D(_02678_),
    .Q(\pcpi_mul.rd[59] ),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__dfxtp_2 _41873_ (.D(_02679_),
    .Q(\pcpi_mul.rd[60] ),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__dfxtp_2 _41874_ (.D(_02680_),
    .Q(\pcpi_mul.rd[61] ),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__dfxtp_2 _41875_ (.D(_02681_),
    .Q(\pcpi_mul.rd[62] ),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__dfxtp_2 _41876_ (.D(_02682_),
    .Q(\pcpi_mul.rd[63] ),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__dfxtp_2 _41877_ (.D(\pcpi_mul.instr_any_mulh ),
    .Q(\pcpi_mul.shift_out ),
    .CLK(clknet_leaf_209_clk));
 sky130_fd_sc_hd__dfxtp_2 _41878_ (.D(_00038_),
    .Q(\cpu_state[0] ),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfxtp_2 _41879_ (.D(_00039_),
    .Q(\cpu_state[1] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__dfxtp_2 _41880_ (.D(_00040_),
    .Q(\cpu_state[2] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__dfxtp_2 _41881_ (.D(_00041_),
    .Q(\cpu_state[3] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__dfxtp_2 _41882_ (.D(_00042_),
    .Q(\cpu_state[4] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__dfxtp_2 _41883_ (.D(_00043_),
    .Q(\cpu_state[5] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__dfxtp_2 _41884_ (.D(_00044_),
    .Q(\cpu_state[6] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__dfxtp_2 _41885_ (.D(_02771_),
    .Q(\cpuregs[8][0] ),
    .CLK(clknet_leaf_243_clk));
 sky130_fd_sc_hd__dfxtp_2 _41886_ (.D(_02772_),
    .Q(\cpuregs[8][1] ),
    .CLK(clknet_leaf_241_clk));
 sky130_fd_sc_hd__dfxtp_2 _41887_ (.D(_02773_),
    .Q(\cpuregs[8][2] ),
    .CLK(clknet_leaf_138_clk));
 sky130_fd_sc_hd__dfxtp_2 _41888_ (.D(_02774_),
    .Q(\cpuregs[8][3] ),
    .CLK(clknet_leaf_142_clk));
 sky130_fd_sc_hd__dfxtp_2 _41889_ (.D(_02775_),
    .Q(\cpuregs[8][4] ),
    .CLK(clknet_leaf_128_clk));
 sky130_fd_sc_hd__dfxtp_2 _41890_ (.D(_02776_),
    .Q(\cpuregs[8][5] ),
    .CLK(clknet_leaf_130_clk));
 sky130_fd_sc_hd__dfxtp_2 _41891_ (.D(_02777_),
    .Q(\cpuregs[8][6] ),
    .CLK(clknet_leaf_132_clk));
 sky130_fd_sc_hd__dfxtp_2 _41892_ (.D(_02778_),
    .Q(\cpuregs[8][7] ),
    .CLK(clknet_leaf_142_clk));
 sky130_fd_sc_hd__dfxtp_2 _41893_ (.D(_02779_),
    .Q(\cpuregs[8][8] ),
    .CLK(clknet_leaf_160_clk));
 sky130_fd_sc_hd__dfxtp_2 _41894_ (.D(_02780_),
    .Q(\cpuregs[8][9] ),
    .CLK(clknet_leaf_146_clk));
 sky130_fd_sc_hd__dfxtp_2 _41895_ (.D(_02781_),
    .Q(\cpuregs[8][10] ),
    .CLK(clknet_leaf_147_clk));
 sky130_fd_sc_hd__dfxtp_2 _41896_ (.D(_02782_),
    .Q(\cpuregs[8][11] ),
    .CLK(clknet_leaf_152_clk));
 sky130_fd_sc_hd__dfxtp_2 _41897_ (.D(_02783_),
    .Q(\cpuregs[8][12] ),
    .CLK(clknet_leaf_158_clk));
 sky130_fd_sc_hd__dfxtp_2 _41898_ (.D(_02784_),
    .Q(\cpuregs[8][13] ),
    .CLK(clknet_leaf_159_clk));
 sky130_fd_sc_hd__dfxtp_2 _41899_ (.D(_02785_),
    .Q(\cpuregs[8][14] ),
    .CLK(clknet_leaf_263_clk));
 sky130_fd_sc_hd__dfxtp_2 _41900_ (.D(_02786_),
    .Q(\cpuregs[8][15] ),
    .CLK(clknet_leaf_263_clk));
 sky130_fd_sc_hd__dfxtp_2 _41901_ (.D(_02787_),
    .Q(\cpuregs[8][16] ),
    .CLK(clknet_leaf_265_clk));
 sky130_fd_sc_hd__dfxtp_2 _41902_ (.D(_02788_),
    .Q(\cpuregs[8][17] ),
    .CLK(clknet_leaf_255_clk));
 sky130_fd_sc_hd__dfxtp_2 _41903_ (.D(_02789_),
    .Q(\cpuregs[8][18] ),
    .CLK(clknet_leaf_269_clk));
 sky130_fd_sc_hd__dfxtp_2 _41904_ (.D(_02790_),
    .Q(\cpuregs[8][19] ),
    .CLK(clknet_leaf_269_clk));
 sky130_fd_sc_hd__dfxtp_2 _41905_ (.D(_02791_),
    .Q(\cpuregs[8][20] ),
    .CLK(clknet_leaf_169_clk));
 sky130_fd_sc_hd__dfxtp_2 _41906_ (.D(_02792_),
    .Q(\cpuregs[8][21] ),
    .CLK(clknet_leaf_174_clk));
 sky130_fd_sc_hd__dfxtp_2 _41907_ (.D(_02793_),
    .Q(\cpuregs[8][22] ),
    .CLK(clknet_leaf_176_clk));
 sky130_fd_sc_hd__dfxtp_2 _41908_ (.D(_02794_),
    .Q(\cpuregs[8][23] ),
    .CLK(clknet_leaf_174_clk));
 sky130_fd_sc_hd__dfxtp_2 _41909_ (.D(_02795_),
    .Q(\cpuregs[8][24] ),
    .CLK(clknet_leaf_176_clk));
 sky130_fd_sc_hd__dfxtp_2 _41910_ (.D(_02796_),
    .Q(\cpuregs[8][25] ),
    .CLK(clknet_leaf_169_clk));
 sky130_fd_sc_hd__dfxtp_2 _41911_ (.D(_02797_),
    .Q(\cpuregs[8][26] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__dfxtp_2 _41912_ (.D(_02798_),
    .Q(\cpuregs[8][27] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__dfxtp_2 _41913_ (.D(_02799_),
    .Q(\cpuregs[8][28] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__dfxtp_2 _41914_ (.D(_02800_),
    .Q(\cpuregs[8][29] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__dfxtp_2 _41915_ (.D(_02801_),
    .Q(\cpuregs[8][30] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__dfxtp_2 _41916_ (.D(_02802_),
    .Q(\cpuregs[8][31] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__dfxtp_2 _41917_ (.D(_02803_),
    .Q(\cpuregs[14][0] ),
    .CLK(clknet_leaf_243_clk));
 sky130_fd_sc_hd__dfxtp_2 _41918_ (.D(_02804_),
    .Q(\cpuregs[14][1] ),
    .CLK(clknet_leaf_241_clk));
 sky130_fd_sc_hd__dfxtp_2 _41919_ (.D(_02805_),
    .Q(\cpuregs[14][2] ),
    .CLK(clknet_leaf_138_clk));
 sky130_fd_sc_hd__dfxtp_2 _41920_ (.D(_02806_),
    .Q(\cpuregs[14][3] ),
    .CLK(clknet_leaf_145_clk));
 sky130_fd_sc_hd__dfxtp_2 _41921_ (.D(_02807_),
    .Q(\cpuregs[14][4] ),
    .CLK(clknet_leaf_128_clk));
 sky130_fd_sc_hd__dfxtp_2 _41922_ (.D(_02808_),
    .Q(\cpuregs[14][5] ),
    .CLK(clknet_leaf_128_clk));
 sky130_fd_sc_hd__dfxtp_2 _41923_ (.D(_02809_),
    .Q(\cpuregs[14][6] ),
    .CLK(clknet_leaf_133_clk));
 sky130_fd_sc_hd__dfxtp_2 _41924_ (.D(_02810_),
    .Q(\cpuregs[14][7] ),
    .CLK(clknet_leaf_142_clk));
 sky130_fd_sc_hd__dfxtp_2 _41925_ (.D(_02811_),
    .Q(\cpuregs[14][8] ),
    .CLK(clknet_leaf_153_clk));
 sky130_fd_sc_hd__dfxtp_2 _41926_ (.D(_02812_),
    .Q(\cpuregs[14][9] ),
    .CLK(clknet_leaf_151_clk));
 sky130_fd_sc_hd__dfxtp_2 _41927_ (.D(_02813_),
    .Q(\cpuregs[14][10] ),
    .CLK(clknet_leaf_151_clk));
 sky130_fd_sc_hd__dfxtp_2 _41928_ (.D(_02814_),
    .Q(\cpuregs[14][11] ),
    .CLK(clknet_leaf_152_clk));
 sky130_fd_sc_hd__dfxtp_2 _41929_ (.D(_02815_),
    .Q(\cpuregs[14][12] ),
    .CLK(clknet_leaf_157_clk));
 sky130_fd_sc_hd__dfxtp_2 _41930_ (.D(_02816_),
    .Q(\cpuregs[14][13] ),
    .CLK(clknet_leaf_153_clk));
 sky130_fd_sc_hd__dfxtp_2 _41931_ (.D(_02817_),
    .Q(\cpuregs[14][14] ),
    .CLK(clknet_leaf_262_clk));
 sky130_fd_sc_hd__dfxtp_2 _41932_ (.D(_02818_),
    .Q(\cpuregs[14][15] ),
    .CLK(clknet_leaf_260_clk));
 sky130_fd_sc_hd__dfxtp_2 _41933_ (.D(_02819_),
    .Q(\cpuregs[14][16] ),
    .CLK(clknet_leaf_266_clk));
 sky130_fd_sc_hd__dfxtp_2 _41934_ (.D(_02820_),
    .Q(\cpuregs[14][17] ),
    .CLK(clknet_leaf_259_clk));
 sky130_fd_sc_hd__dfxtp_2 _41935_ (.D(_02821_),
    .Q(\cpuregs[14][18] ),
    .CLK(clknet_leaf_267_clk));
 sky130_fd_sc_hd__dfxtp_2 _41936_ (.D(_02822_),
    .Q(\cpuregs[14][19] ),
    .CLK(clknet_leaf_267_clk));
 sky130_fd_sc_hd__dfxtp_2 _41937_ (.D(_02823_),
    .Q(\cpuregs[14][20] ),
    .CLK(clknet_leaf_169_clk));
 sky130_fd_sc_hd__dfxtp_2 _41938_ (.D(_02824_),
    .Q(\cpuregs[14][21] ),
    .CLK(clknet_leaf_174_clk));
 sky130_fd_sc_hd__dfxtp_2 _41939_ (.D(_02825_),
    .Q(\cpuregs[14][22] ),
    .CLK(clknet_leaf_176_clk));
 sky130_fd_sc_hd__dfxtp_2 _41940_ (.D(_02826_),
    .Q(\cpuregs[14][23] ),
    .CLK(clknet_leaf_172_clk));
 sky130_fd_sc_hd__dfxtp_2 _41941_ (.D(_02827_),
    .Q(\cpuregs[14][24] ),
    .CLK(clknet_leaf_178_clk));
 sky130_fd_sc_hd__dfxtp_2 _41942_ (.D(_02828_),
    .Q(\cpuregs[14][25] ),
    .CLK(clknet_leaf_169_clk));
 sky130_fd_sc_hd__dfxtp_2 _41943_ (.D(_02829_),
    .Q(\cpuregs[14][26] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__dfxtp_2 _41944_ (.D(_02830_),
    .Q(\cpuregs[14][27] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__dfxtp_2 _41945_ (.D(_02831_),
    .Q(\cpuregs[14][28] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__dfxtp_2 _41946_ (.D(_02832_),
    .Q(\cpuregs[14][29] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__dfxtp_2 _41947_ (.D(_02833_),
    .Q(\cpuregs[14][30] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__dfxtp_2 _41948_ (.D(_02834_),
    .Q(\cpuregs[14][31] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__dfxtp_2 _41949_ (.D(_02835_),
    .Q(\cpuregs[0][0] ),
    .CLK(clknet_leaf_259_clk));
 sky130_fd_sc_hd__dfxtp_2 _41950_ (.D(_02836_),
    .Q(\cpuregs[0][1] ),
    .CLK(clknet_leaf_242_clk));
 sky130_fd_sc_hd__dfxtp_2 _41951_ (.D(_02837_),
    .Q(\cpuregs[0][2] ),
    .CLK(clknet_leaf_138_clk));
 sky130_fd_sc_hd__dfxtp_2 _41952_ (.D(_02838_),
    .Q(\cpuregs[0][3] ),
    .CLK(clknet_leaf_145_clk));
 sky130_fd_sc_hd__dfxtp_2 _41953_ (.D(_02839_),
    .Q(\cpuregs[0][4] ),
    .CLK(clknet_leaf_126_clk));
 sky130_fd_sc_hd__dfxtp_2 _41954_ (.D(_02840_),
    .Q(\cpuregs[0][5] ),
    .CLK(clknet_leaf_131_clk));
 sky130_fd_sc_hd__dfxtp_2 _41955_ (.D(_02841_),
    .Q(\cpuregs[0][6] ),
    .CLK(clknet_leaf_131_clk));
 sky130_fd_sc_hd__dfxtp_2 _41956_ (.D(_02842_),
    .Q(\cpuregs[0][7] ),
    .CLK(clknet_leaf_143_clk));
 sky130_fd_sc_hd__dfxtp_2 _41957_ (.D(_02843_),
    .Q(\cpuregs[0][8] ),
    .CLK(clknet_leaf_153_clk));
 sky130_fd_sc_hd__dfxtp_2 _41958_ (.D(_02844_),
    .Q(\cpuregs[0][9] ),
    .CLK(clknet_leaf_148_clk));
 sky130_fd_sc_hd__dfxtp_2 _41959_ (.D(_02845_),
    .Q(\cpuregs[0][10] ),
    .CLK(clknet_leaf_148_clk));
 sky130_fd_sc_hd__dfxtp_2 _41960_ (.D(_02846_),
    .Q(\cpuregs[0][11] ),
    .CLK(clknet_leaf_149_clk));
 sky130_fd_sc_hd__dfxtp_2 _41961_ (.D(_02847_),
    .Q(\cpuregs[0][12] ),
    .CLK(clknet_leaf_157_clk));
 sky130_fd_sc_hd__dfxtp_2 _41962_ (.D(_02848_),
    .Q(\cpuregs[0][13] ),
    .CLK(clknet_leaf_157_clk));
 sky130_fd_sc_hd__dfxtp_2 _41963_ (.D(_02849_),
    .Q(\cpuregs[0][14] ),
    .CLK(clknet_leaf_266_clk));
 sky130_fd_sc_hd__dfxtp_2 _41964_ (.D(_02850_),
    .Q(\cpuregs[0][15] ),
    .CLK(clknet_leaf_261_clk));
 sky130_fd_sc_hd__dfxtp_2 _41965_ (.D(_02851_),
    .Q(\cpuregs[0][16] ),
    .CLK(clknet_leaf_267_clk));
 sky130_fd_sc_hd__dfxtp_2 _41966_ (.D(_02852_),
    .Q(\cpuregs[0][17] ),
    .CLK(clknet_leaf_259_clk));
 sky130_fd_sc_hd__dfxtp_2 _41967_ (.D(_02853_),
    .Q(\cpuregs[0][18] ),
    .CLK(clknet_leaf_268_clk));
 sky130_fd_sc_hd__dfxtp_2 _41968_ (.D(_02854_),
    .Q(\cpuregs[0][19] ),
    .CLK(clknet_leaf_269_clk));
 sky130_fd_sc_hd__dfxtp_2 _41969_ (.D(_02855_),
    .Q(\cpuregs[0][20] ),
    .CLK(clknet_leaf_156_clk));
 sky130_fd_sc_hd__dfxtp_2 _41970_ (.D(_02856_),
    .Q(\cpuregs[0][21] ),
    .CLK(clknet_leaf_173_clk));
 sky130_fd_sc_hd__dfxtp_2 _41971_ (.D(_02857_),
    .Q(\cpuregs[0][22] ),
    .CLK(clknet_leaf_181_clk));
 sky130_fd_sc_hd__dfxtp_2 _41972_ (.D(_02858_),
    .Q(\cpuregs[0][23] ),
    .CLK(clknet_leaf_172_clk));
 sky130_fd_sc_hd__dfxtp_2 _41973_ (.D(_02859_),
    .Q(\cpuregs[0][24] ),
    .CLK(clknet_leaf_179_clk));
 sky130_fd_sc_hd__dfxtp_2 _41974_ (.D(_02860_),
    .Q(\cpuregs[0][25] ),
    .CLK(clknet_leaf_157_clk));
 sky130_fd_sc_hd__dfxtp_2 _41975_ (.D(_02861_),
    .Q(\cpuregs[0][26] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__dfxtp_2 _41976_ (.D(_02862_),
    .Q(\cpuregs[0][27] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__dfxtp_2 _41977_ (.D(_02863_),
    .Q(\cpuregs[0][28] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__dfxtp_2 _41978_ (.D(_02864_),
    .Q(\cpuregs[0][29] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__dfxtp_2 _41979_ (.D(_02865_),
    .Q(\cpuregs[0][30] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__dfxtp_2 _41980_ (.D(_02866_),
    .Q(\cpuregs[0][31] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfxtp_2 _41981_ (.D(_02867_),
    .Q(\cpuregs[10][0] ),
    .CLK(clknet_leaf_243_clk));
 sky130_fd_sc_hd__dfxtp_2 _41982_ (.D(_02868_),
    .Q(\cpuregs[10][1] ),
    .CLK(clknet_leaf_241_clk));
 sky130_fd_sc_hd__dfxtp_2 _41983_ (.D(_02869_),
    .Q(\cpuregs[10][2] ),
    .CLK(clknet_leaf_137_clk));
 sky130_fd_sc_hd__dfxtp_2 _41984_ (.D(_02870_),
    .Q(\cpuregs[10][3] ),
    .CLK(clknet_leaf_145_clk));
 sky130_fd_sc_hd__dfxtp_2 _41985_ (.D(_02871_),
    .Q(\cpuregs[10][4] ),
    .CLK(clknet_leaf_126_clk));
 sky130_fd_sc_hd__dfxtp_2 _41986_ (.D(_02872_),
    .Q(\cpuregs[10][5] ),
    .CLK(clknet_leaf_130_clk));
 sky130_fd_sc_hd__dfxtp_2 _41987_ (.D(_02873_),
    .Q(\cpuregs[10][6] ),
    .CLK(clknet_leaf_132_clk));
 sky130_fd_sc_hd__dfxtp_2 _41988_ (.D(_02874_),
    .Q(\cpuregs[10][7] ),
    .CLK(clknet_leaf_142_clk));
 sky130_fd_sc_hd__dfxtp_2 _41989_ (.D(_02875_),
    .Q(\cpuregs[10][8] ),
    .CLK(clknet_leaf_160_clk));
 sky130_fd_sc_hd__dfxtp_2 _41990_ (.D(_02876_),
    .Q(\cpuregs[10][9] ),
    .CLK(clknet_leaf_145_clk));
 sky130_fd_sc_hd__dfxtp_2 _41991_ (.D(_02877_),
    .Q(\cpuregs[10][10] ),
    .CLK(clknet_leaf_146_clk));
 sky130_fd_sc_hd__dfxtp_2 _41992_ (.D(_02878_),
    .Q(\cpuregs[10][11] ),
    .CLK(clknet_leaf_146_clk));
 sky130_fd_sc_hd__dfxtp_2 _41993_ (.D(_02879_),
    .Q(\cpuregs[10][12] ),
    .CLK(clknet_leaf_161_clk));
 sky130_fd_sc_hd__dfxtp_2 _41994_ (.D(_02880_),
    .Q(\cpuregs[10][13] ),
    .CLK(clknet_leaf_159_clk));
 sky130_fd_sc_hd__dfxtp_2 _41995_ (.D(_02881_),
    .Q(\cpuregs[10][14] ),
    .CLK(clknet_leaf_263_clk));
 sky130_fd_sc_hd__dfxtp_2 _41996_ (.D(_02882_),
    .Q(\cpuregs[10][15] ),
    .CLK(clknet_leaf_263_clk));
 sky130_fd_sc_hd__dfxtp_2 _41997_ (.D(_02883_),
    .Q(\cpuregs[10][16] ),
    .CLK(clknet_leaf_264_clk));
 sky130_fd_sc_hd__dfxtp_2 _41998_ (.D(_02884_),
    .Q(\cpuregs[10][17] ),
    .CLK(clknet_leaf_255_clk));
 sky130_fd_sc_hd__dfxtp_2 _41999_ (.D(_02885_),
    .Q(\cpuregs[10][18] ),
    .CLK(clknet_leaf_269_clk));
 sky130_fd_sc_hd__dfxtp_2 _42000_ (.D(_02886_),
    .Q(\cpuregs[10][19] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__dfxtp_2 _42001_ (.D(_02887_),
    .Q(\cpuregs[10][20] ),
    .CLK(clknet_leaf_170_clk));
 sky130_fd_sc_hd__dfxtp_2 _42002_ (.D(_02888_),
    .Q(\cpuregs[10][21] ),
    .CLK(clknet_leaf_174_clk));
 sky130_fd_sc_hd__dfxtp_2 _42003_ (.D(_02889_),
    .Q(\cpuregs[10][22] ),
    .CLK(clknet_leaf_175_clk));
 sky130_fd_sc_hd__dfxtp_2 _42004_ (.D(_02890_),
    .Q(\cpuregs[10][23] ),
    .CLK(clknet_leaf_167_clk));
 sky130_fd_sc_hd__dfxtp_2 _42005_ (.D(_02891_),
    .Q(\cpuregs[10][24] ),
    .CLK(clknet_leaf_177_clk));
 sky130_fd_sc_hd__dfxtp_2 _42006_ (.D(_02892_),
    .Q(\cpuregs[10][25] ),
    .CLK(clknet_leaf_169_clk));
 sky130_fd_sc_hd__dfxtp_2 _42007_ (.D(_02893_),
    .Q(\cpuregs[10][26] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__dfxtp_2 _42008_ (.D(_02894_),
    .Q(\cpuregs[10][27] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__dfxtp_2 _42009_ (.D(_02895_),
    .Q(\cpuregs[10][28] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__dfxtp_2 _42010_ (.D(_02896_),
    .Q(\cpuregs[10][29] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__dfxtp_2 _42011_ (.D(_02897_),
    .Q(\cpuregs[10][30] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__dfxtp_2 _42012_ (.D(_02898_),
    .Q(\cpuregs[10][31] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__dfxtp_2 _42013_ (.D(_02899_),
    .Q(\cpuregs[18][0] ),
    .CLK(clknet_leaf_258_clk));
 sky130_fd_sc_hd__dfxtp_2 _42014_ (.D(_02900_),
    .Q(\cpuregs[18][1] ),
    .CLK(clknet_leaf_243_clk));
 sky130_fd_sc_hd__dfxtp_2 _42015_ (.D(_02901_),
    .Q(\cpuregs[18][2] ),
    .CLK(clknet_leaf_137_clk));
 sky130_fd_sc_hd__dfxtp_2 _42016_ (.D(_02902_),
    .Q(\cpuregs[18][3] ),
    .CLK(clknet_leaf_140_clk));
 sky130_fd_sc_hd__dfxtp_2 _42017_ (.D(_02903_),
    .Q(\cpuregs[18][4] ),
    .CLK(clknet_leaf_128_clk));
 sky130_fd_sc_hd__dfxtp_2 _42018_ (.D(_02904_),
    .Q(\cpuregs[18][5] ),
    .CLK(clknet_leaf_129_clk));
 sky130_fd_sc_hd__dfxtp_2 _42019_ (.D(_02905_),
    .Q(\cpuregs[18][6] ),
    .CLK(clknet_leaf_133_clk));
 sky130_fd_sc_hd__dfxtp_2 _42020_ (.D(_02906_),
    .Q(\cpuregs[18][7] ),
    .CLK(clknet_leaf_142_clk));
 sky130_fd_sc_hd__dfxtp_2 _42021_ (.D(_02907_),
    .Q(\cpuregs[18][8] ),
    .CLK(clknet_leaf_160_clk));
 sky130_fd_sc_hd__dfxtp_2 _42022_ (.D(_02908_),
    .Q(\cpuregs[18][9] ),
    .CLK(clknet_leaf_146_clk));
 sky130_fd_sc_hd__dfxtp_2 _42023_ (.D(_02909_),
    .Q(\cpuregs[18][10] ),
    .CLK(clknet_leaf_146_clk));
 sky130_fd_sc_hd__dfxtp_2 _42024_ (.D(_02910_),
    .Q(\cpuregs[18][11] ),
    .CLK(clknet_leaf_160_clk));
 sky130_fd_sc_hd__dfxtp_2 _42025_ (.D(_02911_),
    .Q(\cpuregs[18][12] ),
    .CLK(clknet_leaf_161_clk));
 sky130_fd_sc_hd__dfxtp_2 _42026_ (.D(_02912_),
    .Q(\cpuregs[18][13] ),
    .CLK(clknet_leaf_161_clk));
 sky130_fd_sc_hd__dfxtp_2 _42027_ (.D(_02913_),
    .Q(\cpuregs[18][14] ),
    .CLK(clknet_leaf_264_clk));
 sky130_fd_sc_hd__dfxtp_2 _42028_ (.D(_02914_),
    .Q(\cpuregs[18][15] ),
    .CLK(clknet_leaf_254_clk));
 sky130_fd_sc_hd__dfxtp_2 _42029_ (.D(_02915_),
    .Q(\cpuregs[18][16] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__dfxtp_2 _42030_ (.D(_02916_),
    .Q(\cpuregs[18][17] ),
    .CLK(clknet_leaf_255_clk));
 sky130_fd_sc_hd__dfxtp_2 _42031_ (.D(_02917_),
    .Q(\cpuregs[18][18] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__dfxtp_2 _42032_ (.D(_02918_),
    .Q(\cpuregs[18][19] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__dfxtp_2 _42033_ (.D(_02919_),
    .Q(\cpuregs[18][20] ),
    .CLK(clknet_leaf_157_clk));
 sky130_fd_sc_hd__dfxtp_2 _42034_ (.D(_02920_),
    .Q(\cpuregs[18][21] ),
    .CLK(clknet_leaf_174_clk));
 sky130_fd_sc_hd__dfxtp_2 _42035_ (.D(_02921_),
    .Q(\cpuregs[18][22] ),
    .CLK(clknet_leaf_176_clk));
 sky130_fd_sc_hd__dfxtp_2 _42036_ (.D(_02922_),
    .Q(\cpuregs[18][23] ),
    .CLK(clknet_leaf_167_clk));
 sky130_fd_sc_hd__dfxtp_2 _42037_ (.D(_02923_),
    .Q(\cpuregs[18][24] ),
    .CLK(clknet_leaf_175_clk));
 sky130_fd_sc_hd__dfxtp_2 _42038_ (.D(_02924_),
    .Q(\cpuregs[18][25] ),
    .CLK(clknet_leaf_158_clk));
 sky130_fd_sc_hd__dfxtp_2 _42039_ (.D(_02925_),
    .Q(\cpuregs[18][26] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__dfxtp_2 _42040_ (.D(_02926_),
    .Q(\cpuregs[18][27] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__dfxtp_2 _42041_ (.D(_02927_),
    .Q(\cpuregs[18][28] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__dfxtp_2 _42042_ (.D(_02928_),
    .Q(\cpuregs[18][29] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__dfxtp_2 _42043_ (.D(_02929_),
    .Q(\cpuregs[18][30] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__dfxtp_2 _42044_ (.D(_02930_),
    .Q(\cpuregs[18][31] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__dfxtp_2 _42045_ (.D(_02931_),
    .Q(\mem_rdata_q[0] ),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__dfxtp_2 _42046_ (.D(_02932_),
    .Q(\mem_rdata_q[1] ),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__dfxtp_2 _42047_ (.D(_02933_),
    .Q(\mem_rdata_q[2] ),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__dfxtp_2 _42048_ (.D(_02934_),
    .Q(\mem_rdata_q[3] ),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__dfxtp_2 _42049_ (.D(_02935_),
    .Q(\mem_rdata_q[4] ),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__dfxtp_2 _42050_ (.D(_02936_),
    .Q(\mem_rdata_q[5] ),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__dfxtp_2 _42051_ (.D(_02937_),
    .Q(\mem_rdata_q[6] ),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__dfxtp_2 _42052_ (.D(_02938_),
    .Q(\mem_rdata_q[7] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__dfxtp_2 _42053_ (.D(_02939_),
    .Q(\mem_rdata_q[8] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__dfxtp_2 _42054_ (.D(_02940_),
    .Q(\mem_rdata_q[9] ),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__dfxtp_2 _42055_ (.D(_02941_),
    .Q(\mem_rdata_q[10] ),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__dfxtp_2 _42056_ (.D(_02942_),
    .Q(\mem_rdata_q[11] ),
    .CLK(clknet_leaf_209_clk));
 sky130_fd_sc_hd__dfxtp_2 _42057_ (.D(_02943_),
    .Q(\mem_rdata_q[12] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__dfxtp_2 _42058_ (.D(_02944_),
    .Q(\mem_rdata_q[13] ),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__dfxtp_2 _42059_ (.D(_02945_),
    .Q(\mem_rdata_q[14] ),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__dfxtp_2 _42060_ (.D(_02946_),
    .Q(\mem_rdata_q[15] ),
    .CLK(clknet_leaf_211_clk));
 sky130_fd_sc_hd__dfxtp_2 _42061_ (.D(_02947_),
    .Q(\mem_rdata_q[16] ),
    .CLK(clknet_leaf_211_clk));
 sky130_fd_sc_hd__dfxtp_2 _42062_ (.D(_02948_),
    .Q(\mem_rdata_q[17] ),
    .CLK(clknet_leaf_211_clk));
 sky130_fd_sc_hd__dfxtp_2 _42063_ (.D(_02949_),
    .Q(\mem_rdata_q[18] ),
    .CLK(clknet_leaf_212_clk));
 sky130_fd_sc_hd__dfxtp_2 _42064_ (.D(_02950_),
    .Q(\mem_rdata_q[19] ),
    .CLK(clknet_leaf_209_clk));
 sky130_fd_sc_hd__dfxtp_2 _42065_ (.D(_02951_),
    .Q(\mem_rdata_q[20] ),
    .CLK(clknet_leaf_213_clk));
 sky130_fd_sc_hd__dfxtp_2 _42066_ (.D(_02952_),
    .Q(\mem_rdata_q[21] ),
    .CLK(clknet_leaf_211_clk));
 sky130_fd_sc_hd__dfxtp_2 _42067_ (.D(_02953_),
    .Q(\mem_rdata_q[22] ),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__dfxtp_2 _42068_ (.D(_02954_),
    .Q(\mem_rdata_q[23] ),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__dfxtp_2 _42069_ (.D(_02955_),
    .Q(\mem_rdata_q[24] ),
    .CLK(clknet_leaf_211_clk));
 sky130_fd_sc_hd__dfxtp_2 _42070_ (.D(_02956_),
    .Q(\mem_rdata_q[25] ),
    .CLK(clknet_leaf_211_clk));
 sky130_fd_sc_hd__dfxtp_2 _42071_ (.D(_02957_),
    .Q(\mem_rdata_q[26] ),
    .CLK(clknet_leaf_211_clk));
 sky130_fd_sc_hd__dfxtp_2 _42072_ (.D(_02958_),
    .Q(\mem_rdata_q[27] ),
    .CLK(clknet_leaf_213_clk));
 sky130_fd_sc_hd__dfxtp_2 _42073_ (.D(_02959_),
    .Q(\mem_rdata_q[28] ),
    .CLK(clknet_leaf_219_clk));
 sky130_fd_sc_hd__dfxtp_2 _42074_ (.D(_02960_),
    .Q(\mem_rdata_q[29] ),
    .CLK(clknet_leaf_215_clk));
 sky130_fd_sc_hd__dfxtp_2 _42075_ (.D(_02961_),
    .Q(\mem_rdata_q[30] ),
    .CLK(clknet_leaf_209_clk));
 sky130_fd_sc_hd__dfxtp_2 _42076_ (.D(_02962_),
    .Q(\mem_rdata_q[31] ),
    .CLK(clknet_leaf_214_clk));
 sky130_fd_sc_hd__dfxtp_2 _42077_ (.D(_02963_),
    .Q(\cpuregs[2][0] ),
    .CLK(clknet_leaf_258_clk));
 sky130_fd_sc_hd__dfxtp_2 _42078_ (.D(_02964_),
    .Q(\cpuregs[2][1] ),
    .CLK(clknet_leaf_242_clk));
 sky130_fd_sc_hd__dfxtp_2 _42079_ (.D(_02965_),
    .Q(\cpuregs[2][2] ),
    .CLK(clknet_leaf_138_clk));
 sky130_fd_sc_hd__dfxtp_2 _42080_ (.D(_02966_),
    .Q(\cpuregs[2][3] ),
    .CLK(clknet_leaf_145_clk));
 sky130_fd_sc_hd__dfxtp_2 _42081_ (.D(_02967_),
    .Q(\cpuregs[2][4] ),
    .CLK(clknet_leaf_126_clk));
 sky130_fd_sc_hd__dfxtp_2 _42082_ (.D(_02968_),
    .Q(\cpuregs[2][5] ),
    .CLK(clknet_leaf_130_clk));
 sky130_fd_sc_hd__dfxtp_2 _42083_ (.D(_02969_),
    .Q(\cpuregs[2][6] ),
    .CLK(clknet_leaf_131_clk));
 sky130_fd_sc_hd__dfxtp_2 _42084_ (.D(_02970_),
    .Q(\cpuregs[2][7] ),
    .CLK(clknet_leaf_127_clk));
 sky130_fd_sc_hd__dfxtp_2 _42085_ (.D(_02971_),
    .Q(\cpuregs[2][8] ),
    .CLK(clknet_leaf_154_clk));
 sky130_fd_sc_hd__dfxtp_2 _42086_ (.D(_02972_),
    .Q(\cpuregs[2][9] ),
    .CLK(clknet_leaf_147_clk));
 sky130_fd_sc_hd__dfxtp_2 _42087_ (.D(_02973_),
    .Q(\cpuregs[2][10] ),
    .CLK(clknet_leaf_149_clk));
 sky130_fd_sc_hd__dfxtp_2 _42088_ (.D(_02974_),
    .Q(\cpuregs[2][11] ),
    .CLK(clknet_leaf_149_clk));
 sky130_fd_sc_hd__dfxtp_2 _42089_ (.D(_02975_),
    .Q(\cpuregs[2][12] ),
    .CLK(clknet_leaf_157_clk));
 sky130_fd_sc_hd__dfxtp_2 _42090_ (.D(_02976_),
    .Q(\cpuregs[2][13] ),
    .CLK(clknet_leaf_159_clk));
 sky130_fd_sc_hd__dfxtp_2 _42091_ (.D(_02977_),
    .Q(\cpuregs[2][14] ),
    .CLK(clknet_leaf_261_clk));
 sky130_fd_sc_hd__dfxtp_2 _42092_ (.D(_02978_),
    .Q(\cpuregs[2][15] ),
    .CLK(clknet_leaf_260_clk));
 sky130_fd_sc_hd__dfxtp_2 _42093_ (.D(_02979_),
    .Q(\cpuregs[2][16] ),
    .CLK(clknet_leaf_266_clk));
 sky130_fd_sc_hd__dfxtp_2 _42094_ (.D(_02980_),
    .Q(\cpuregs[2][17] ),
    .CLK(clknet_leaf_259_clk));
 sky130_fd_sc_hd__dfxtp_2 _42095_ (.D(_02981_),
    .Q(\cpuregs[2][18] ),
    .CLK(clknet_leaf_268_clk));
 sky130_fd_sc_hd__dfxtp_2 _42096_ (.D(_02982_),
    .Q(\cpuregs[2][19] ),
    .CLK(clknet_leaf_268_clk));
 sky130_fd_sc_hd__dfxtp_2 _42097_ (.D(_02983_),
    .Q(\cpuregs[2][20] ),
    .CLK(clknet_leaf_156_clk));
 sky130_fd_sc_hd__dfxtp_2 _42098_ (.D(_02984_),
    .Q(\cpuregs[2][21] ),
    .CLK(clknet_leaf_172_clk));
 sky130_fd_sc_hd__dfxtp_2 _42099_ (.D(_02985_),
    .Q(\cpuregs[2][22] ),
    .CLK(clknet_leaf_179_clk));
 sky130_fd_sc_hd__dfxtp_2 _42100_ (.D(_02986_),
    .Q(\cpuregs[2][23] ),
    .CLK(clknet_leaf_172_clk));
 sky130_fd_sc_hd__dfxtp_2 _42101_ (.D(_02987_),
    .Q(\cpuregs[2][24] ),
    .CLK(clknet_leaf_179_clk));
 sky130_fd_sc_hd__dfxtp_2 _42102_ (.D(_02988_),
    .Q(\cpuregs[2][25] ),
    .CLK(clknet_leaf_156_clk));
 sky130_fd_sc_hd__dfxtp_2 _42103_ (.D(_02989_),
    .Q(\cpuregs[2][26] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__dfxtp_2 _42104_ (.D(_02990_),
    .Q(\cpuregs[2][27] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfxtp_2 _42105_ (.D(_02991_),
    .Q(\cpuregs[2][28] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__dfxtp_2 _42106_ (.D(_02992_),
    .Q(\cpuregs[2][29] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__dfxtp_2 _42107_ (.D(_02993_),
    .Q(\cpuregs[2][30] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__dfxtp_2 _42108_ (.D(_02994_),
    .Q(\cpuregs[2][31] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__dfxtp_2 _42109_ (.D(_02995_),
    .Q(\cpuregs[5][0] ),
    .CLK(clknet_leaf_258_clk));
 sky130_fd_sc_hd__dfxtp_2 _42110_ (.D(_02996_),
    .Q(\cpuregs[5][1] ),
    .CLK(clknet_leaf_242_clk));
 sky130_fd_sc_hd__dfxtp_2 _42111_ (.D(_02997_),
    .Q(\cpuregs[5][2] ),
    .CLK(clknet_leaf_139_clk));
 sky130_fd_sc_hd__dfxtp_2 _42112_ (.D(_02998_),
    .Q(\cpuregs[5][3] ),
    .CLK(clknet_leaf_143_clk));
 sky130_fd_sc_hd__dfxtp_2 _42113_ (.D(_02999_),
    .Q(\cpuregs[5][4] ),
    .CLK(clknet_leaf_127_clk));
 sky130_fd_sc_hd__dfxtp_2 _42114_ (.D(_03000_),
    .Q(\cpuregs[5][5] ),
    .CLK(clknet_leaf_129_clk));
 sky130_fd_sc_hd__dfxtp_2 _42115_ (.D(_03001_),
    .Q(\cpuregs[5][6] ),
    .CLK(clknet_leaf_132_clk));
 sky130_fd_sc_hd__dfxtp_2 _42116_ (.D(_03002_),
    .Q(\cpuregs[5][7] ),
    .CLK(clknet_leaf_142_clk));
 sky130_fd_sc_hd__dfxtp_2 _42117_ (.D(_03003_),
    .Q(\cpuregs[5][8] ),
    .CLK(clknet_leaf_153_clk));
 sky130_fd_sc_hd__dfxtp_2 _42118_ (.D(_03004_),
    .Q(\cpuregs[5][9] ),
    .CLK(clknet_leaf_150_clk));
 sky130_fd_sc_hd__dfxtp_2 _42119_ (.D(_03005_),
    .Q(\cpuregs[5][10] ),
    .CLK(clknet_leaf_150_clk));
 sky130_fd_sc_hd__dfxtp_2 _42120_ (.D(_03006_),
    .Q(\cpuregs[5][11] ),
    .CLK(clknet_leaf_154_clk));
 sky130_fd_sc_hd__dfxtp_2 _42121_ (.D(_03007_),
    .Q(\cpuregs[5][12] ),
    .CLK(clknet_leaf_157_clk));
 sky130_fd_sc_hd__dfxtp_2 _42122_ (.D(_03008_),
    .Q(\cpuregs[5][13] ),
    .CLK(clknet_leaf_155_clk));
 sky130_fd_sc_hd__dfxtp_2 _42123_ (.D(_03009_),
    .Q(\cpuregs[5][14] ),
    .CLK(clknet_leaf_261_clk));
 sky130_fd_sc_hd__dfxtp_2 _42124_ (.D(_03010_),
    .Q(\cpuregs[5][15] ),
    .CLK(clknet_leaf_261_clk));
 sky130_fd_sc_hd__dfxtp_2 _42125_ (.D(_03011_),
    .Q(\cpuregs[5][16] ),
    .CLK(clknet_leaf_266_clk));
 sky130_fd_sc_hd__dfxtp_2 _42126_ (.D(_03012_),
    .Q(\cpuregs[5][17] ),
    .CLK(clknet_leaf_259_clk));
 sky130_fd_sc_hd__dfxtp_2 _42127_ (.D(_03013_),
    .Q(\cpuregs[5][18] ),
    .CLK(clknet_leaf_268_clk));
 sky130_fd_sc_hd__dfxtp_2 _42128_ (.D(_03014_),
    .Q(\cpuregs[5][19] ),
    .CLK(clknet_leaf_268_clk));
 sky130_fd_sc_hd__dfxtp_2 _42129_ (.D(_03015_),
    .Q(\cpuregs[5][20] ),
    .CLK(clknet_leaf_171_clk));
 sky130_fd_sc_hd__dfxtp_2 _42130_ (.D(_03016_),
    .Q(\cpuregs[5][21] ),
    .CLK(clknet_leaf_173_clk));
 sky130_fd_sc_hd__dfxtp_2 _42131_ (.D(_03017_),
    .Q(\cpuregs[5][22] ),
    .CLK(clknet_leaf_178_clk));
 sky130_fd_sc_hd__dfxtp_2 _42132_ (.D(_03018_),
    .Q(\cpuregs[5][23] ),
    .CLK(clknet_leaf_172_clk));
 sky130_fd_sc_hd__dfxtp_2 _42133_ (.D(_03019_),
    .Q(\cpuregs[5][24] ),
    .CLK(clknet_leaf_179_clk));
 sky130_fd_sc_hd__dfxtp_2 _42134_ (.D(_03020_),
    .Q(\cpuregs[5][25] ),
    .CLK(clknet_leaf_171_clk));
 sky130_fd_sc_hd__dfxtp_2 _42135_ (.D(_03021_),
    .Q(\cpuregs[5][26] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__dfxtp_2 _42136_ (.D(_03022_),
    .Q(\cpuregs[5][27] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__dfxtp_2 _42137_ (.D(_03023_),
    .Q(\cpuregs[5][28] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__dfxtp_2 _42138_ (.D(_03024_),
    .Q(\cpuregs[5][29] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__dfxtp_2 _42139_ (.D(_03025_),
    .Q(\cpuregs[5][30] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__dfxtp_2 _42140_ (.D(_03026_),
    .Q(\cpuregs[5][31] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__dfxtp_2 _42141_ (.D(_03027_),
    .Q(\pcpi_mul.rs1[0] ),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__dfxtp_2 _42142_ (.D(_03028_),
    .Q(\pcpi_mul.rs1[1] ),
    .CLK(clknet_opt_26_clk));
 sky130_fd_sc_hd__dfxtp_2 _42143_ (.D(_03029_),
    .Q(\pcpi_mul.rs1[2] ),
    .CLK(clknet_leaf_105_clk));
 sky130_fd_sc_hd__dfxtp_2 _42144_ (.D(_03030_),
    .Q(\pcpi_mul.rs1[3] ),
    .CLK(clknet_leaf_105_clk));
 sky130_fd_sc_hd__dfxtp_2 _42145_ (.D(_03031_),
    .Q(\pcpi_mul.rs1[4] ),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__dfxtp_2 _42146_ (.D(_03032_),
    .Q(\pcpi_mul.rs1[5] ),
    .CLK(clknet_leaf_105_clk));
 sky130_fd_sc_hd__dfxtp_2 _42147_ (.D(_03033_),
    .Q(\pcpi_mul.rs1[6] ),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__dfxtp_2 _42148_ (.D(_03034_),
    .Q(\pcpi_mul.rs1[7] ),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__dfxtp_2 _42149_ (.D(_03035_),
    .Q(\pcpi_mul.rs1[8] ),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__dfxtp_2 _42150_ (.D(_03036_),
    .Q(\pcpi_mul.rs1[9] ),
    .CLK(clknet_5_22_0_clk));
 sky130_fd_sc_hd__dfxtp_2 _42151_ (.D(_03037_),
    .Q(\pcpi_mul.rs1[10] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__dfxtp_2 _42152_ (.D(_03038_),
    .Q(\pcpi_mul.rs1[11] ),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__dfxtp_2 _42153_ (.D(_03039_),
    .Q(\pcpi_mul.rs1[12] ),
    .CLK(clknet_leaf_87_clk));
 sky130_fd_sc_hd__dfxtp_2 _42154_ (.D(_03040_),
    .Q(\pcpi_mul.rs1[13] ),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__dfxtp_2 _42155_ (.D(_03041_),
    .Q(\pcpi_mul.rs1[14] ),
    .CLK(clknet_leaf_87_clk));
 sky130_fd_sc_hd__dfxtp_2 _42156_ (.D(_03042_),
    .Q(\pcpi_mul.rs1[15] ),
    .CLK(clknet_leaf_87_clk));
 sky130_fd_sc_hd__dfxtp_2 _42157_ (.D(_03043_),
    .Q(\pcpi_mul.rs1[16] ),
    .CLK(clknet_leaf_87_clk));
 sky130_fd_sc_hd__dfxtp_2 _42158_ (.D(_03044_),
    .Q(\pcpi_mul.rs1[17] ),
    .CLK(clknet_leaf_89_clk));
 sky130_fd_sc_hd__dfxtp_2 _42159_ (.D(_03045_),
    .Q(\pcpi_mul.rs1[18] ),
    .CLK(clknet_leaf_89_clk));
 sky130_fd_sc_hd__dfxtp_2 _42160_ (.D(_03046_),
    .Q(\pcpi_mul.rs1[19] ),
    .CLK(clknet_leaf_89_clk));
 sky130_fd_sc_hd__dfxtp_2 _42161_ (.D(_03047_),
    .Q(\pcpi_mul.rs1[20] ),
    .CLK(clknet_leaf_90_clk));
 sky130_fd_sc_hd__dfxtp_2 _42162_ (.D(_03048_),
    .Q(\pcpi_mul.rs1[21] ),
    .CLK(clknet_leaf_90_clk));
 sky130_fd_sc_hd__dfxtp_2 _42163_ (.D(_03049_),
    .Q(\pcpi_mul.rs1[22] ),
    .CLK(clknet_leaf_90_clk));
 sky130_fd_sc_hd__dfxtp_2 _42164_ (.D(_03050_),
    .Q(\pcpi_mul.rs1[23] ),
    .CLK(clknet_leaf_90_clk));
 sky130_fd_sc_hd__dfxtp_2 _42165_ (.D(_03051_),
    .Q(\pcpi_mul.rs1[24] ),
    .CLK(clknet_leaf_91_clk));
 sky130_fd_sc_hd__dfxtp_2 _42166_ (.D(_03052_),
    .Q(\pcpi_mul.rs1[25] ),
    .CLK(clknet_leaf_90_clk));
 sky130_fd_sc_hd__dfxtp_2 _42167_ (.D(_03053_),
    .Q(\pcpi_mul.rs1[26] ),
    .CLK(clknet_leaf_91_clk));
 sky130_fd_sc_hd__dfxtp_2 _42168_ (.D(_03054_),
    .Q(\pcpi_mul.rs1[27] ),
    .CLK(clknet_leaf_92_clk));
 sky130_fd_sc_hd__dfxtp_2 _42169_ (.D(_03055_),
    .Q(\pcpi_mul.rs1[28] ),
    .CLK(clknet_leaf_92_clk));
 sky130_fd_sc_hd__dfxtp_2 _42170_ (.D(_03056_),
    .Q(\pcpi_mul.rs1[29] ),
    .CLK(clknet_leaf_92_clk));
 sky130_fd_sc_hd__dfxtp_2 _42171_ (.D(_03057_),
    .Q(\pcpi_mul.rs1[30] ),
    .CLK(clknet_opt_2_clk));
 sky130_fd_sc_hd__dfxtp_2 _42172_ (.D(_03058_),
    .Q(\pcpi_mul.rs1[31] ),
    .CLK(clknet_leaf_91_clk));
 sky130_fd_sc_hd__dfxtp_2 _42173_ (.D(_03059_),
    .Q(mem_addr[2]),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__dfxtp_2 _42174_ (.D(_03060_),
    .Q(mem_addr[3]),
    .CLK(clknet_leaf_109_clk));
 sky130_fd_sc_hd__dfxtp_2 _42175_ (.D(_03061_),
    .Q(mem_addr[4]),
    .CLK(clknet_leaf_240_clk));
 sky130_fd_sc_hd__dfxtp_2 _42176_ (.D(_03062_),
    .Q(mem_addr[5]),
    .CLK(clknet_leaf_240_clk));
 sky130_fd_sc_hd__dfxtp_2 _42177_ (.D(_03063_),
    .Q(mem_addr[6]),
    .CLK(clknet_leaf_126_clk));
 sky130_fd_sc_hd__dfxtp_2 _42178_ (.D(_03064_),
    .Q(mem_addr[7]),
    .CLK(clknet_leaf_117_clk));
 sky130_fd_sc_hd__dfxtp_2 _42179_ (.D(_03065_),
    .Q(mem_addr[8]),
    .CLK(clknet_leaf_166_clk));
 sky130_fd_sc_hd__dfxtp_2 _42180_ (.D(_03066_),
    .Q(mem_addr[9]),
    .CLK(clknet_5_21_0_clk));
 sky130_fd_sc_hd__dfxtp_2 _42181_ (.D(_03067_),
    .Q(mem_addr[10]),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__dfxtp_2 _42182_ (.D(_03068_),
    .Q(mem_addr[11]),
    .CLK(clknet_leaf_149_clk));
 sky130_fd_sc_hd__dfxtp_2 _42183_ (.D(_03069_),
    .Q(mem_addr[12]),
    .CLK(clknet_leaf_125_clk));
 sky130_fd_sc_hd__dfxtp_2 _42184_ (.D(_03070_),
    .Q(mem_addr[13]),
    .CLK(clknet_leaf_125_clk));
 sky130_fd_sc_hd__dfxtp_2 _42185_ (.D(_03071_),
    .Q(mem_addr[14]),
    .CLK(clknet_leaf_240_clk));
 sky130_fd_sc_hd__dfxtp_2 _42186_ (.D(_03072_),
    .Q(mem_addr[15]),
    .CLK(clknet_leaf_180_clk));
 sky130_fd_sc_hd__dfxtp_2 _42187_ (.D(_03073_),
    .Q(mem_addr[16]),
    .CLK(clknet_opt_30_clk));
 sky130_fd_sc_hd__dfxtp_2 _42188_ (.D(_03074_),
    .Q(mem_addr[17]),
    .CLK(clknet_opt_21_clk));
 sky130_fd_sc_hd__dfxtp_2 _42189_ (.D(_03075_),
    .Q(mem_addr[18]),
    .CLK(clknet_leaf_161_clk));
 sky130_fd_sc_hd__dfxtp_2 _42190_ (.D(_03076_),
    .Q(mem_addr[19]),
    .CLK(clknet_leaf_240_clk));
 sky130_fd_sc_hd__dfxtp_2 _42191_ (.D(_03077_),
    .Q(mem_addr[20]),
    .CLK(clknet_leaf_122_clk));
 sky130_fd_sc_hd__dfxtp_2 _42192_ (.D(_03078_),
    .Q(mem_addr[21]),
    .CLK(clknet_leaf_138_clk));
 sky130_fd_sc_hd__dfxtp_2 _42193_ (.D(_03079_),
    .Q(mem_addr[22]),
    .CLK(clknet_opt_0_clk));
 sky130_fd_sc_hd__dfxtp_2 _42194_ (.D(_03080_),
    .Q(mem_addr[23]),
    .CLK(clknet_leaf_175_clk));
 sky130_fd_sc_hd__dfxtp_2 _42195_ (.D(_03081_),
    .Q(mem_addr[24]),
    .CLK(clknet_leaf_183_clk));
 sky130_fd_sc_hd__dfxtp_2 _42196_ (.D(_03082_),
    .Q(mem_addr[25]),
    .CLK(clknet_leaf_138_clk));
 sky130_fd_sc_hd__dfxtp_2 _42197_ (.D(_03083_),
    .Q(mem_addr[26]),
    .CLK(clknet_leaf_136_clk));
 sky130_fd_sc_hd__dfxtp_2 _42198_ (.D(_03084_),
    .Q(mem_addr[27]),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__dfxtp_2 _42199_ (.D(_03085_),
    .Q(mem_addr[28]),
    .CLK(clknet_leaf_148_clk));
 sky130_fd_sc_hd__dfxtp_2 _42200_ (.D(_03086_),
    .Q(mem_addr[29]),
    .CLK(clknet_leaf_124_clk));
 sky130_fd_sc_hd__dfxtp_2 _42201_ (.D(_03087_),
    .Q(mem_addr[30]),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__dfxtp_2 _42202_ (.D(_03088_),
    .Q(mem_addr[31]),
    .CLK(clknet_leaf_171_clk));
 sky130_fd_sc_hd__dfxtp_2 _42203_ (.D(_03089_),
    .Q(pcpi_rs1[0]),
    .CLK(clknet_leaf_202_clk));
 sky130_fd_sc_hd__dfxtp_2 _42204_ (.D(_03090_),
    .Q(pcpi_rs1[1]),
    .CLK(clknet_leaf_204_clk));
 sky130_fd_sc_hd__dfxtp_2 _42205_ (.D(_03091_),
    .Q(pcpi_rs1[2]),
    .CLK(clknet_leaf_204_clk));
 sky130_fd_sc_hd__dfxtp_2 _42206_ (.D(_03092_),
    .Q(pcpi_rs1[3]),
    .CLK(clknet_leaf_109_clk));
 sky130_fd_sc_hd__dfxtp_2 _42207_ (.D(_03093_),
    .Q(pcpi_rs1[4]),
    .CLK(clknet_leaf_113_clk));
 sky130_fd_sc_hd__dfxtp_2 _42208_ (.D(_03094_),
    .Q(pcpi_rs1[5]),
    .CLK(clknet_leaf_196_clk));
 sky130_fd_sc_hd__dfxtp_2 _42209_ (.D(_03095_),
    .Q(pcpi_rs1[6]),
    .CLK(clknet_leaf_196_clk));
 sky130_fd_sc_hd__dfxtp_2 _42210_ (.D(_03096_),
    .Q(pcpi_rs1[7]),
    .CLK(clknet_leaf_196_clk));
 sky130_fd_sc_hd__dfxtp_2 _42211_ (.D(_03097_),
    .Q(pcpi_rs1[8]),
    .CLK(clknet_leaf_195_clk));
 sky130_fd_sc_hd__dfxtp_2 _42212_ (.D(_03098_),
    .Q(pcpi_rs1[9]),
    .CLK(clknet_leaf_199_clk));
 sky130_fd_sc_hd__dfxtp_2 _42213_ (.D(_03099_),
    .Q(pcpi_rs1[10]),
    .CLK(clknet_leaf_199_clk));
 sky130_fd_sc_hd__dfxtp_2 _42214_ (.D(_03100_),
    .Q(pcpi_rs1[11]),
    .CLK(clknet_leaf_199_clk));
 sky130_fd_sc_hd__dfxtp_2 _42215_ (.D(_03101_),
    .Q(pcpi_rs1[12]),
    .CLK(clknet_leaf_187_clk));
 sky130_fd_sc_hd__dfxtp_2 _42216_ (.D(_03102_),
    .Q(pcpi_rs1[13]),
    .CLK(clknet_leaf_192_clk));
 sky130_fd_sc_hd__dfxtp_2 _42217_ (.D(_03103_),
    .Q(pcpi_rs1[14]),
    .CLK(clknet_leaf_182_clk));
 sky130_fd_sc_hd__dfxtp_2 _42218_ (.D(_03104_),
    .Q(pcpi_rs1[15]),
    .CLK(clknet_leaf_182_clk));
 sky130_fd_sc_hd__dfxtp_2 _42219_ (.D(_03105_),
    .Q(pcpi_rs1[16]),
    .CLK(clknet_leaf_183_clk));
 sky130_fd_sc_hd__dfxtp_2 _42220_ (.D(_03106_),
    .Q(pcpi_rs1[17]),
    .CLK(clknet_leaf_183_clk));
 sky130_fd_sc_hd__dfxtp_2 _42221_ (.D(_03107_),
    .Q(pcpi_rs1[18]),
    .CLK(clknet_leaf_184_clk));
 sky130_fd_sc_hd__dfxtp_2 _42222_ (.D(_03108_),
    .Q(pcpi_rs1[19]),
    .CLK(clknet_leaf_175_clk));
 sky130_fd_sc_hd__dfxtp_2 _42223_ (.D(_03109_),
    .Q(pcpi_rs1[20]),
    .CLK(clknet_leaf_166_clk));
 sky130_fd_sc_hd__dfxtp_2 _42224_ (.D(_03110_),
    .Q(pcpi_rs1[21]),
    .CLK(clknet_leaf_166_clk));
 sky130_fd_sc_hd__dfxtp_2 _42225_ (.D(_03111_),
    .Q(pcpi_rs1[22]),
    .CLK(clknet_leaf_190_clk));
 sky130_fd_sc_hd__dfxtp_2 _42226_ (.D(_03112_),
    .Q(pcpi_rs1[23]),
    .CLK(clknet_leaf_190_clk));
 sky130_fd_sc_hd__dfxtp_2 _42227_ (.D(_03113_),
    .Q(pcpi_rs1[24]),
    .CLK(clknet_leaf_191_clk));
 sky130_fd_sc_hd__dfxtp_2 _42228_ (.D(_03114_),
    .Q(pcpi_rs1[25]),
    .CLK(clknet_leaf_191_clk));
 sky130_fd_sc_hd__dfxtp_2 _42229_ (.D(_03115_),
    .Q(pcpi_rs1[26]),
    .CLK(clknet_leaf_188_clk));
 sky130_fd_sc_hd__dfxtp_2 _42230_ (.D(_03116_),
    .Q(pcpi_rs1[27]),
    .CLK(clknet_leaf_188_clk));
 sky130_fd_sc_hd__dfxtp_2 _42231_ (.D(_03117_),
    .Q(pcpi_rs1[28]),
    .CLK(clknet_leaf_198_clk));
 sky130_fd_sc_hd__dfxtp_2 _42232_ (.D(_03118_),
    .Q(pcpi_rs1[29]),
    .CLK(clknet_leaf_198_clk));
 sky130_fd_sc_hd__dfxtp_2 _42233_ (.D(_03119_),
    .Q(pcpi_rs1[30]),
    .CLK(clknet_leaf_197_clk));
 sky130_fd_sc_hd__dfxtp_2 _42234_ (.D(_03120_),
    .Q(pcpi_rs1[31]),
    .CLK(clknet_leaf_196_clk));
 sky130_fd_sc_hd__dfxtp_2 _42235_ (.D(_03121_),
    .Q(pcpi_insn[0]),
    .CLK(clknet_leaf_209_clk));
 sky130_fd_sc_hd__dfxtp_2 _42236_ (.D(_03122_),
    .Q(pcpi_insn[1]),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__dfxtp_2 _42237_ (.D(_03123_),
    .Q(pcpi_insn[2]),
    .CLK(clknet_leaf_209_clk));
 sky130_fd_sc_hd__dfxtp_2 _42238_ (.D(_03124_),
    .Q(pcpi_insn[3]),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__dfxtp_2 _42239_ (.D(_03125_),
    .Q(pcpi_insn[4]),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__dfxtp_2 _42240_ (.D(_03126_),
    .Q(pcpi_insn[5]),
    .CLK(clknet_leaf_209_clk));
 sky130_fd_sc_hd__dfxtp_2 _42241_ (.D(_03127_),
    .Q(pcpi_insn[6]),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__dfxtp_2 _42242_ (.D(_03128_),
    .Q(pcpi_insn[7]),
    .CLK(clknet_leaf_209_clk));
 sky130_fd_sc_hd__dfxtp_2 _42243_ (.D(_03129_),
    .Q(pcpi_insn[8]),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__dfxtp_2 _42244_ (.D(_03130_),
    .Q(pcpi_insn[9]),
    .CLK(clknet_leaf_208_clk));
 sky130_fd_sc_hd__dfxtp_2 _42245_ (.D(_03131_),
    .Q(pcpi_insn[10]),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__dfxtp_2 _42246_ (.D(_03132_),
    .Q(pcpi_insn[11]),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__dfxtp_2 _42247_ (.D(_03133_),
    .Q(pcpi_insn[12]),
    .CLK(clknet_leaf_209_clk));
 sky130_fd_sc_hd__dfxtp_2 _42248_ (.D(_03134_),
    .Q(pcpi_insn[13]),
    .CLK(clknet_leaf_208_clk));
 sky130_fd_sc_hd__dfxtp_2 _42249_ (.D(_03135_),
    .Q(pcpi_insn[14]),
    .CLK(clknet_leaf_208_clk));
 sky130_fd_sc_hd__dfxtp_2 _42250_ (.D(_03136_),
    .Q(pcpi_insn[15]),
    .CLK(clknet_leaf_216_clk));
 sky130_fd_sc_hd__dfxtp_2 _42251_ (.D(_03137_),
    .Q(pcpi_insn[16]),
    .CLK(clknet_leaf_217_clk));
 sky130_fd_sc_hd__dfxtp_2 _42252_ (.D(_03138_),
    .Q(pcpi_insn[17]),
    .CLK(clknet_leaf_205_clk));
 sky130_fd_sc_hd__dfxtp_2 _42253_ (.D(_03139_),
    .Q(pcpi_insn[18]),
    .CLK(clknet_leaf_205_clk));
 sky130_fd_sc_hd__dfxtp_2 _42254_ (.D(_03140_),
    .Q(pcpi_insn[19]),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__dfxtp_2 _42255_ (.D(_03141_),
    .Q(pcpi_insn[20]),
    .CLK(clknet_leaf_206_clk));
 sky130_fd_sc_hd__dfxtp_2 _42256_ (.D(_03142_),
    .Q(pcpi_insn[21]),
    .CLK(clknet_leaf_210_clk));
 sky130_fd_sc_hd__dfxtp_2 _42257_ (.D(_03143_),
    .Q(pcpi_insn[22]),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__dfxtp_2 _42258_ (.D(_03144_),
    .Q(pcpi_insn[23]),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__dfxtp_2 _42259_ (.D(_03145_),
    .Q(pcpi_insn[24]),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__dfxtp_2 _42260_ (.D(_03146_),
    .Q(pcpi_insn[25]),
    .CLK(clknet_leaf_209_clk));
 sky130_fd_sc_hd__dfxtp_2 _42261_ (.D(_03147_),
    .Q(pcpi_insn[26]),
    .CLK(clknet_leaf_209_clk));
 sky130_fd_sc_hd__dfxtp_2 _42262_ (.D(_03148_),
    .Q(pcpi_insn[27]),
    .CLK(clknet_leaf_206_clk));
 sky130_fd_sc_hd__dfxtp_2 _42263_ (.D(_03149_),
    .Q(pcpi_insn[28]),
    .CLK(clknet_leaf_210_clk));
 sky130_fd_sc_hd__dfxtp_2 _42264_ (.D(_03150_),
    .Q(pcpi_insn[29]),
    .CLK(clknet_leaf_206_clk));
 sky130_fd_sc_hd__dfxtp_2 _42265_ (.D(_03151_),
    .Q(pcpi_insn[30]),
    .CLK(clknet_leaf_209_clk));
 sky130_fd_sc_hd__dfxtp_2 _42266_ (.D(_03152_),
    .Q(pcpi_insn[31]),
    .CLK(clknet_leaf_210_clk));
 sky130_fd_sc_hd__dfxtp_2 _42267_ (.D(_03153_),
    .Q(instr_lui),
    .CLK(clknet_leaf_212_clk));
 sky130_fd_sc_hd__dfxtp_2 _42268_ (.D(_03154_),
    .Q(instr_auipc),
    .CLK(clknet_leaf_212_clk));
 sky130_fd_sc_hd__dfxtp_2 _42269_ (.D(_03155_),
    .Q(instr_jal),
    .CLK(clknet_leaf_219_clk));
 sky130_fd_sc_hd__dfxtp_2 _42270_ (.D(_03156_),
    .Q(instr_jalr),
    .CLK(clknet_leaf_219_clk));
 sky130_fd_sc_hd__dfxtp_2 _42271_ (.D(_03157_),
    .Q(instr_lb),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__dfxtp_2 _42272_ (.D(_03158_),
    .Q(instr_lh),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__dfxtp_2 _42273_ (.D(_03159_),
    .Q(instr_lw),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__dfxtp_2 _42274_ (.D(_03160_),
    .Q(instr_lbu),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__dfxtp_2 _42275_ (.D(_03161_),
    .Q(instr_lhu),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__dfxtp_2 _42276_ (.D(_03162_),
    .Q(instr_sb),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__dfxtp_2 _42277_ (.D(_03163_),
    .Q(instr_sh),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__dfxtp_2 _42278_ (.D(_03164_),
    .Q(instr_sw),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__dfxtp_2 _42279_ (.D(_03165_),
    .Q(instr_slli),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__dfxtp_2 _42280_ (.D(_03166_),
    .Q(instr_srli),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__dfxtp_2 _42281_ (.D(_03167_),
    .Q(instr_srai),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__dfxtp_2 _42282_ (.D(_03168_),
    .Q(instr_rdcycle),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__dfxtp_2 _42283_ (.D(_03169_),
    .Q(instr_rdcycleh),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__dfxtp_2 _42284_ (.D(_03170_),
    .Q(instr_rdinstr),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__dfxtp_2 _42285_ (.D(_03171_),
    .Q(instr_rdinstrh),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__dfxtp_2 _42286_ (.D(_03172_),
    .Q(instr_ecall_ebreak),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__dfxtp_2 _42287_ (.D(_03173_),
    .Q(instr_getq),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__dfxtp_2 _42288_ (.D(_03174_),
    .Q(instr_setq),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__dfxtp_2 _42289_ (.D(_03175_),
    .Q(instr_retirq),
    .CLK(clknet_leaf_222_clk));
 sky130_fd_sc_hd__dfxtp_2 _42290_ (.D(_03176_),
    .Q(instr_maskirq),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__dfxtp_2 _42291_ (.D(_03177_),
    .Q(instr_waitirq),
    .CLK(clknet_leaf_219_clk));
 sky130_fd_sc_hd__dfxtp_2 _42292_ (.D(_03178_),
    .Q(instr_timer),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__dfxtp_2 _42293_ (.D(_03179_),
    .Q(\decoded_rd[0] ),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__dfxtp_2 _42294_ (.D(_03180_),
    .Q(\decoded_rd[1] ),
    .CLK(clknet_leaf_207_clk));
 sky130_fd_sc_hd__dfxtp_2 _42295_ (.D(_03181_),
    .Q(\decoded_rd[2] ),
    .CLK(clknet_leaf_206_clk));
 sky130_fd_sc_hd__dfxtp_2 _42296_ (.D(_03182_),
    .Q(\decoded_rd[3] ),
    .CLK(clknet_leaf_202_clk));
 sky130_fd_sc_hd__dfxtp_2 _42297_ (.D(_03183_),
    .Q(\decoded_rd[4] ),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__dfxtp_2 _42298_ (.D(_03184_),
    .Q(\decoded_imm[0] ),
    .CLK(clknet_leaf_213_clk));
 sky130_fd_sc_hd__dfxtp_2 _42299_ (.D(_03185_),
    .Q(\decoded_imm_uj[1] ),
    .CLK(clknet_leaf_212_clk));
 sky130_fd_sc_hd__dfxtp_2 _42300_ (.D(_03186_),
    .Q(\decoded_imm_uj[2] ),
    .CLK(clknet_leaf_213_clk));
 sky130_fd_sc_hd__dfxtp_2 _42301_ (.D(_03187_),
    .Q(\decoded_imm_uj[3] ),
    .CLK(clknet_leaf_211_clk));
 sky130_fd_sc_hd__dfxtp_2 _42302_ (.D(_03188_),
    .Q(\decoded_imm_uj[4] ),
    .CLK(clknet_leaf_211_clk));
 sky130_fd_sc_hd__dfxtp_2 _42303_ (.D(_03189_),
    .Q(\decoded_imm_uj[5] ),
    .CLK(clknet_leaf_213_clk));
 sky130_fd_sc_hd__dfxtp_2 _42304_ (.D(_03190_),
    .Q(\decoded_imm_uj[6] ),
    .CLK(clknet_leaf_213_clk));
 sky130_fd_sc_hd__dfxtp_2 _42305_ (.D(_03191_),
    .Q(\decoded_imm_uj[7] ),
    .CLK(clknet_leaf_215_clk));
 sky130_fd_sc_hd__dfxtp_2 _42306_ (.D(_03192_),
    .Q(\decoded_imm_uj[8] ),
    .CLK(clknet_leaf_213_clk));
 sky130_fd_sc_hd__dfxtp_2 _42307_ (.D(_03193_),
    .Q(\decoded_imm_uj[9] ),
    .CLK(clknet_leaf_215_clk));
 sky130_fd_sc_hd__dfxtp_2 _42308_ (.D(_03194_),
    .Q(\decoded_imm_uj[10] ),
    .CLK(clknet_leaf_215_clk));
 sky130_fd_sc_hd__dfxtp_2 _42309_ (.D(_03195_),
    .Q(\decoded_imm_uj[11] ),
    .CLK(clknet_leaf_213_clk));
 sky130_fd_sc_hd__dfxtp_2 _42310_ (.D(_03196_),
    .Q(\decoded_imm_uj[12] ),
    .CLK(clknet_leaf_217_clk));
 sky130_fd_sc_hd__dfxtp_2 _42311_ (.D(_03197_),
    .Q(\decoded_imm_uj[13] ),
    .CLK(clknet_leaf_217_clk));
 sky130_fd_sc_hd__dfxtp_2 _42312_ (.D(_03198_),
    .Q(\decoded_imm_uj[14] ),
    .CLK(clknet_leaf_215_clk));
 sky130_fd_sc_hd__dfxtp_2 _42313_ (.D(_03199_),
    .Q(\decoded_imm_uj[15] ),
    .CLK(clknet_leaf_216_clk));
 sky130_fd_sc_hd__dfxtp_2 _42314_ (.D(_03200_),
    .Q(\decoded_imm_uj[16] ),
    .CLK(clknet_leaf_216_clk));
 sky130_fd_sc_hd__dfxtp_2 _42315_ (.D(_03201_),
    .Q(\decoded_imm_uj[17] ),
    .CLK(clknet_leaf_216_clk));
 sky130_fd_sc_hd__dfxtp_2 _42316_ (.D(_03202_),
    .Q(\decoded_imm_uj[18] ),
    .CLK(clknet_leaf_217_clk));
 sky130_fd_sc_hd__dfxtp_2 _42317_ (.D(_03203_),
    .Q(\decoded_imm_uj[19] ),
    .CLK(clknet_leaf_217_clk));
 sky130_fd_sc_hd__dfxtp_2 _42318_ (.D(_03204_),
    .Q(\decoded_imm_uj[20] ),
    .CLK(clknet_leaf_236_clk));
 sky130_fd_sc_hd__dfxtp_2 _42319_ (.D(_03205_),
    .Q(is_lb_lh_lw_lbu_lhu),
    .CLK(clknet_leaf_212_clk));
 sky130_fd_sc_hd__dfxtp_2 _42320_ (.D(_03206_),
    .Q(is_slli_srli_srai),
    .CLK(clknet_leaf_205_clk));
 sky130_fd_sc_hd__dfxtp_2 _42321_ (.D(_03207_),
    .Q(is_jalr_addi_slti_sltiu_xori_ori_andi),
    .CLK(clknet_leaf_206_clk));
 sky130_fd_sc_hd__dfxtp_2 _42322_ (.D(_03208_),
    .Q(is_sb_sh_sw),
    .CLK(clknet_leaf_220_clk));
 sky130_fd_sc_hd__dfxtp_2 _42323_ (.D(_03209_),
    .Q(\cpuregs[13][0] ),
    .CLK(clknet_leaf_244_clk));
 sky130_fd_sc_hd__dfxtp_2 _42324_ (.D(_03210_),
    .Q(\cpuregs[13][1] ),
    .CLK(clknet_leaf_239_clk));
 sky130_fd_sc_hd__dfxtp_2 _42325_ (.D(_03211_),
    .Q(\cpuregs[13][2] ),
    .CLK(clknet_leaf_139_clk));
 sky130_fd_sc_hd__dfxtp_2 _42326_ (.D(_03212_),
    .Q(\cpuregs[13][3] ),
    .CLK(clknet_leaf_140_clk));
 sky130_fd_sc_hd__dfxtp_2 _42327_ (.D(_03213_),
    .Q(\cpuregs[13][4] ),
    .CLK(clknet_leaf_128_clk));
 sky130_fd_sc_hd__dfxtp_2 _42328_ (.D(_03214_),
    .Q(\cpuregs[13][5] ),
    .CLK(clknet_leaf_129_clk));
 sky130_fd_sc_hd__dfxtp_2 _42329_ (.D(_03215_),
    .Q(\cpuregs[13][6] ),
    .CLK(clknet_leaf_133_clk));
 sky130_fd_sc_hd__dfxtp_2 _42330_ (.D(_03216_),
    .Q(\cpuregs[13][7] ),
    .CLK(clknet_leaf_142_clk));
 sky130_fd_sc_hd__dfxtp_2 _42331_ (.D(_03217_),
    .Q(\cpuregs[13][8] ),
    .CLK(clknet_leaf_159_clk));
 sky130_fd_sc_hd__dfxtp_2 _42332_ (.D(_03218_),
    .Q(\cpuregs[13][9] ),
    .CLK(clknet_leaf_152_clk));
 sky130_fd_sc_hd__dfxtp_2 _42333_ (.D(_03219_),
    .Q(\cpuregs[13][10] ),
    .CLK(clknet_leaf_152_clk));
 sky130_fd_sc_hd__dfxtp_2 _42334_ (.D(_03220_),
    .Q(\cpuregs[13][11] ),
    .CLK(clknet_leaf_152_clk));
 sky130_fd_sc_hd__dfxtp_2 _42335_ (.D(_03221_),
    .Q(\cpuregs[13][12] ),
    .CLK(clknet_leaf_158_clk));
 sky130_fd_sc_hd__dfxtp_2 _42336_ (.D(_03222_),
    .Q(\cpuregs[13][13] ),
    .CLK(clknet_leaf_159_clk));
 sky130_fd_sc_hd__dfxtp_2 _42337_ (.D(_03223_),
    .Q(\cpuregs[13][14] ),
    .CLK(clknet_leaf_263_clk));
 sky130_fd_sc_hd__dfxtp_2 _42338_ (.D(_03224_),
    .Q(\cpuregs[13][15] ),
    .CLK(clknet_leaf_257_clk));
 sky130_fd_sc_hd__dfxtp_2 _42339_ (.D(_03225_),
    .Q(\cpuregs[13][16] ),
    .CLK(clknet_leaf_264_clk));
 sky130_fd_sc_hd__dfxtp_2 _42340_ (.D(_03226_),
    .Q(\cpuregs[13][17] ),
    .CLK(clknet_leaf_257_clk));
 sky130_fd_sc_hd__dfxtp_2 _42341_ (.D(_03227_),
    .Q(\cpuregs[13][18] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__dfxtp_2 _42342_ (.D(_03228_),
    .Q(\cpuregs[13][19] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__dfxtp_2 _42343_ (.D(_03229_),
    .Q(\cpuregs[13][20] ),
    .CLK(clknet_leaf_167_clk));
 sky130_fd_sc_hd__dfxtp_2 _42344_ (.D(_03230_),
    .Q(\cpuregs[13][21] ),
    .CLK(clknet_leaf_175_clk));
 sky130_fd_sc_hd__dfxtp_2 _42345_ (.D(_03231_),
    .Q(\cpuregs[13][22] ),
    .CLK(clknet_leaf_182_clk));
 sky130_fd_sc_hd__dfxtp_2 _42346_ (.D(_03232_),
    .Q(\cpuregs[13][23] ),
    .CLK(clknet_leaf_174_clk));
 sky130_fd_sc_hd__dfxtp_2 _42347_ (.D(_03233_),
    .Q(\cpuregs[13][24] ),
    .CLK(clknet_leaf_183_clk));
 sky130_fd_sc_hd__dfxtp_2 _42348_ (.D(_03234_),
    .Q(\cpuregs[13][25] ),
    .CLK(clknet_leaf_167_clk));
 sky130_fd_sc_hd__dfxtp_2 _42349_ (.D(_03235_),
    .Q(\cpuregs[13][26] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__dfxtp_2 _42350_ (.D(_03236_),
    .Q(\cpuregs[13][27] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__dfxtp_2 _42351_ (.D(_03237_),
    .Q(\cpuregs[13][28] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__dfxtp_2 _42352_ (.D(_03238_),
    .Q(\cpuregs[13][29] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__dfxtp_2 _42353_ (.D(_03239_),
    .Q(\cpuregs[13][30] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__dfxtp_2 _42354_ (.D(_03240_),
    .Q(\cpuregs[13][31] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__dfxtp_2 _42355_ (.D(_03241_),
    .Q(is_alu_reg_imm),
    .CLK(clknet_leaf_212_clk));
 sky130_fd_sc_hd__dfxtp_2 _42356_ (.D(_03242_),
    .Q(is_alu_reg_reg),
    .CLK(clknet_leaf_212_clk));
 sky130_fd_sc_hd__dfxtp_2 _42357_ (.D(_03243_),
    .Q(mem_wstrb[0]),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__dfxtp_2 _42358_ (.D(_03244_),
    .Q(mem_wstrb[1]),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__dfxtp_2 _42359_ (.D(_03245_),
    .Q(mem_wstrb[2]),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__dfxtp_2 _42360_ (.D(_03246_),
    .Q(mem_wstrb[3]),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__dfxtp_2 _42361_ (.D(_03247_),
    .Q(\pcpi_mul.rs2[0] ),
    .CLK(clknet_leaf_105_clk));
 sky130_fd_sc_hd__dfxtp_2 _42362_ (.D(_03248_),
    .Q(\pcpi_mul.rs2[1] ),
    .CLK(clknet_leaf_105_clk));
 sky130_fd_sc_hd__dfxtp_2 _42363_ (.D(_03249_),
    .Q(\pcpi_mul.rs2[2] ),
    .CLK(clknet_leaf_208_clk));
 sky130_fd_sc_hd__dfxtp_2 _42364_ (.D(_03250_),
    .Q(\pcpi_mul.rs2[3] ),
    .CLK(clknet_leaf_105_clk));
 sky130_fd_sc_hd__dfxtp_2 _42365_ (.D(_03251_),
    .Q(\pcpi_mul.rs2[4] ),
    .CLK(clknet_leaf_106_clk));
 sky130_fd_sc_hd__dfxtp_2 _42366_ (.D(_03252_),
    .Q(\pcpi_mul.rs2[5] ),
    .CLK(clknet_leaf_106_clk));
 sky130_fd_sc_hd__dfxtp_2 _42367_ (.D(_03253_),
    .Q(\pcpi_mul.rs2[6] ),
    .CLK(clknet_leaf_106_clk));
 sky130_fd_sc_hd__dfxtp_2 _42368_ (.D(_03254_),
    .Q(\pcpi_mul.rs2[7] ),
    .CLK(clknet_leaf_105_clk));
 sky130_fd_sc_hd__dfxtp_2 _42369_ (.D(_03255_),
    .Q(\pcpi_mul.rs2[8] ),
    .CLK(clknet_leaf_106_clk));
 sky130_fd_sc_hd__dfxtp_2 _42370_ (.D(_03256_),
    .Q(\pcpi_mul.rs2[9] ),
    .CLK(clknet_leaf_107_clk));
 sky130_fd_sc_hd__dfxtp_2 _42371_ (.D(_03257_),
    .Q(\pcpi_mul.rs2[10] ),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__dfxtp_2 _42372_ (.D(_03258_),
    .Q(\pcpi_mul.rs2[11] ),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__dfxtp_2 _42373_ (.D(_03259_),
    .Q(\pcpi_mul.rs2[12] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__dfxtp_2 _42374_ (.D(_03260_),
    .Q(\pcpi_mul.rs2[13] ),
    .CLK(clknet_5_22_0_clk));
 sky130_fd_sc_hd__dfxtp_2 _42375_ (.D(_03261_),
    .Q(\pcpi_mul.rs2[14] ),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__dfxtp_2 _42376_ (.D(_03262_),
    .Q(\pcpi_mul.rs2[15] ),
    .CLK(clknet_leaf_104_clk));
 sky130_fd_sc_hd__dfxtp_2 _42377_ (.D(_03263_),
    .Q(\pcpi_mul.rs2[16] ),
    .CLK(clknet_5_5_0_clk));
 sky130_fd_sc_hd__dfxtp_2 _42378_ (.D(_03264_),
    .Q(\pcpi_mul.rs2[17] ),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__dfxtp_2 _42379_ (.D(_03265_),
    .Q(\pcpi_mul.rs2[18] ),
    .CLK(clknet_leaf_103_clk));
 sky130_fd_sc_hd__dfxtp_2 _42380_ (.D(_03266_),
    .Q(\pcpi_mul.rs2[19] ),
    .CLK(clknet_leaf_103_clk));
 sky130_fd_sc_hd__dfxtp_2 _42381_ (.D(_03267_),
    .Q(\pcpi_mul.rs2[20] ),
    .CLK(clknet_5_13_0_clk));
 sky130_fd_sc_hd__dfxtp_2 _42382_ (.D(_03268_),
    .Q(\pcpi_mul.rs2[21] ),
    .CLK(clknet_leaf_103_clk));
 sky130_fd_sc_hd__dfxtp_2 _42383_ (.D(_03269_),
    .Q(\pcpi_mul.rs2[22] ),
    .CLK(clknet_leaf_107_clk));
 sky130_fd_sc_hd__dfxtp_2 _42384_ (.D(_03270_),
    .Q(\pcpi_mul.rs2[23] ),
    .CLK(clknet_leaf_107_clk));
 sky130_fd_sc_hd__dfxtp_2 _42385_ (.D(_03271_),
    .Q(\pcpi_mul.rs2[24] ),
    .CLK(clknet_leaf_106_clk));
 sky130_fd_sc_hd__dfxtp_2 _42386_ (.D(_03272_),
    .Q(\pcpi_mul.rs2[25] ),
    .CLK(clknet_leaf_107_clk));
 sky130_fd_sc_hd__dfxtp_2 _42387_ (.D(_03273_),
    .Q(\pcpi_mul.rs2[26] ),
    .CLK(clknet_leaf_104_clk));
 sky130_fd_sc_hd__dfxtp_2 _42388_ (.D(_03274_),
    .Q(\pcpi_mul.rs2[27] ),
    .CLK(clknet_opt_5_clk));
 sky130_fd_sc_hd__dfxtp_2 _42389_ (.D(_03275_),
    .Q(\pcpi_mul.rs2[28] ),
    .CLK(clknet_leaf_103_clk));
 sky130_fd_sc_hd__dfxtp_2 _42390_ (.D(_03276_),
    .Q(\pcpi_mul.rs2[29] ),
    .CLK(clknet_leaf_103_clk));
 sky130_fd_sc_hd__dfxtp_2 _42391_ (.D(_03277_),
    .Q(\pcpi_mul.rs2[30] ),
    .CLK(clknet_leaf_91_clk));
 sky130_fd_sc_hd__dfxtp_2 _42392_ (.D(_03278_),
    .Q(\pcpi_mul.rs2[31] ),
    .CLK(clknet_leaf_92_clk));
 sky130_fd_sc_hd__dfxtp_2 _42393_ (.D(_03279_),
    .Q(\cpuregs[17][0] ),
    .CLK(clknet_leaf_257_clk));
 sky130_fd_sc_hd__dfxtp_2 _42394_ (.D(_03280_),
    .Q(\cpuregs[17][1] ),
    .CLK(clknet_leaf_243_clk));
 sky130_fd_sc_hd__dfxtp_2 _42395_ (.D(_03281_),
    .Q(\cpuregs[17][2] ),
    .CLK(clknet_leaf_137_clk));
 sky130_fd_sc_hd__dfxtp_2 _42396_ (.D(_03282_),
    .Q(\cpuregs[17][3] ),
    .CLK(clknet_leaf_140_clk));
 sky130_fd_sc_hd__dfxtp_2 _42397_ (.D(_03283_),
    .Q(\cpuregs[17][4] ),
    .CLK(clknet_leaf_141_clk));
 sky130_fd_sc_hd__dfxtp_2 _42398_ (.D(_03284_),
    .Q(\cpuregs[17][5] ),
    .CLK(clknet_leaf_141_clk));
 sky130_fd_sc_hd__dfxtp_2 _42399_ (.D(_03285_),
    .Q(\cpuregs[17][6] ),
    .CLK(clknet_leaf_136_clk));
 sky130_fd_sc_hd__dfxtp_2 _42400_ (.D(_03286_),
    .Q(\cpuregs[17][7] ),
    .CLK(clknet_leaf_141_clk));
 sky130_fd_sc_hd__dfxtp_2 _42401_ (.D(_03287_),
    .Q(\cpuregs[17][8] ),
    .CLK(clknet_leaf_160_clk));
 sky130_fd_sc_hd__dfxtp_2 _42402_ (.D(_03288_),
    .Q(\cpuregs[17][9] ),
    .CLK(clknet_leaf_139_clk));
 sky130_fd_sc_hd__dfxtp_2 _42403_ (.D(_03289_),
    .Q(\cpuregs[17][10] ),
    .CLK(clknet_leaf_146_clk));
 sky130_fd_sc_hd__dfxtp_2 _42404_ (.D(_03290_),
    .Q(\cpuregs[17][11] ),
    .CLK(clknet_leaf_139_clk));
 sky130_fd_sc_hd__dfxtp_2 _42405_ (.D(_03291_),
    .Q(\cpuregs[17][12] ),
    .CLK(clknet_leaf_161_clk));
 sky130_fd_sc_hd__dfxtp_2 _42406_ (.D(_03292_),
    .Q(\cpuregs[17][13] ),
    .CLK(clknet_leaf_161_clk));
 sky130_fd_sc_hd__dfxtp_2 _42407_ (.D(_03293_),
    .Q(\cpuregs[17][14] ),
    .CLK(clknet_leaf_264_clk));
 sky130_fd_sc_hd__dfxtp_2 _42408_ (.D(_03294_),
    .Q(\cpuregs[17][15] ),
    .CLK(clknet_leaf_254_clk));
 sky130_fd_sc_hd__dfxtp_2 _42409_ (.D(_03295_),
    .Q(\cpuregs[17][16] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__dfxtp_2 _42410_ (.D(_03296_),
    .Q(\cpuregs[17][17] ),
    .CLK(clknet_leaf_254_clk));
 sky130_fd_sc_hd__dfxtp_2 _42411_ (.D(_03297_),
    .Q(\cpuregs[17][18] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__dfxtp_2 _42412_ (.D(_03298_),
    .Q(\cpuregs[17][19] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__dfxtp_2 _42413_ (.D(_03299_),
    .Q(\cpuregs[17][20] ),
    .CLK(clknet_leaf_167_clk));
 sky130_fd_sc_hd__dfxtp_2 _42414_ (.D(_03300_),
    .Q(\cpuregs[17][21] ),
    .CLK(clknet_leaf_175_clk));
 sky130_fd_sc_hd__dfxtp_2 _42415_ (.D(_03301_),
    .Q(\cpuregs[17][22] ),
    .CLK(clknet_leaf_183_clk));
 sky130_fd_sc_hd__dfxtp_2 _42416_ (.D(_03302_),
    .Q(\cpuregs[17][23] ),
    .CLK(clknet_leaf_167_clk));
 sky130_fd_sc_hd__dfxtp_2 _42417_ (.D(_03303_),
    .Q(\cpuregs[17][24] ),
    .CLK(clknet_leaf_175_clk));
 sky130_fd_sc_hd__dfxtp_2 _42418_ (.D(_03304_),
    .Q(\cpuregs[17][25] ),
    .CLK(clknet_leaf_168_clk));
 sky130_fd_sc_hd__dfxtp_2 _42419_ (.D(_03305_),
    .Q(\cpuregs[17][26] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__dfxtp_2 _42420_ (.D(_03306_),
    .Q(\cpuregs[17][27] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__dfxtp_2 _42421_ (.D(_03307_),
    .Q(\cpuregs[17][28] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__dfxtp_2 _42422_ (.D(_03308_),
    .Q(\cpuregs[17][29] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__dfxtp_2 _42423_ (.D(_03309_),
    .Q(\cpuregs[17][30] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__dfxtp_2 _42424_ (.D(_03310_),
    .Q(\cpuregs[17][31] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__dfxtp_2 _42425_ (.D(_03311_),
    .Q(\cpuregs[16][0] ),
    .CLK(clknet_leaf_257_clk));
 sky130_fd_sc_hd__dfxtp_2 _42426_ (.D(_03312_),
    .Q(\cpuregs[16][1] ),
    .CLK(clknet_leaf_244_clk));
 sky130_fd_sc_hd__dfxtp_2 _42427_ (.D(_03313_),
    .Q(\cpuregs[16][2] ),
    .CLK(clknet_leaf_137_clk));
 sky130_fd_sc_hd__dfxtp_2 _42428_ (.D(_03314_),
    .Q(\cpuregs[16][3] ),
    .CLK(clknet_leaf_140_clk));
 sky130_fd_sc_hd__dfxtp_2 _42429_ (.D(_03315_),
    .Q(\cpuregs[16][4] ),
    .CLK(clknet_leaf_141_clk));
 sky130_fd_sc_hd__dfxtp_2 _42430_ (.D(_03316_),
    .Q(\cpuregs[16][5] ),
    .CLK(clknet_leaf_141_clk));
 sky130_fd_sc_hd__dfxtp_2 _42431_ (.D(_03317_),
    .Q(\cpuregs[16][6] ),
    .CLK(clknet_leaf_136_clk));
 sky130_fd_sc_hd__dfxtp_2 _42432_ (.D(_03318_),
    .Q(\cpuregs[16][7] ),
    .CLK(clknet_leaf_141_clk));
 sky130_fd_sc_hd__dfxtp_2 _42433_ (.D(_03319_),
    .Q(\cpuregs[16][8] ),
    .CLK(clknet_leaf_160_clk));
 sky130_fd_sc_hd__dfxtp_2 _42434_ (.D(_03320_),
    .Q(\cpuregs[16][9] ),
    .CLK(clknet_leaf_139_clk));
 sky130_fd_sc_hd__dfxtp_2 _42435_ (.D(_03321_),
    .Q(\cpuregs[16][10] ),
    .CLK(clknet_leaf_146_clk));
 sky130_fd_sc_hd__dfxtp_2 _42436_ (.D(_03322_),
    .Q(\cpuregs[16][11] ),
    .CLK(clknet_leaf_139_clk));
 sky130_fd_sc_hd__dfxtp_2 _42437_ (.D(_03323_),
    .Q(\cpuregs[16][12] ),
    .CLK(clknet_leaf_161_clk));
 sky130_fd_sc_hd__dfxtp_2 _42438_ (.D(_03324_),
    .Q(\cpuregs[16][13] ),
    .CLK(clknet_leaf_161_clk));
 sky130_fd_sc_hd__dfxtp_2 _42439_ (.D(_03325_),
    .Q(\cpuregs[16][14] ),
    .CLK(clknet_leaf_254_clk));
 sky130_fd_sc_hd__dfxtp_2 _42440_ (.D(_03326_),
    .Q(\cpuregs[16][15] ),
    .CLK(clknet_leaf_253_clk));
 sky130_fd_sc_hd__dfxtp_2 _42441_ (.D(_03327_),
    .Q(\cpuregs[16][16] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__dfxtp_2 _42442_ (.D(_03328_),
    .Q(\cpuregs[16][17] ),
    .CLK(clknet_leaf_254_clk));
 sky130_fd_sc_hd__dfxtp_2 _42443_ (.D(_03329_),
    .Q(\cpuregs[16][18] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__dfxtp_2 _42444_ (.D(_03330_),
    .Q(\cpuregs[16][19] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__dfxtp_2 _42445_ (.D(_03331_),
    .Q(\cpuregs[16][20] ),
    .CLK(clknet_leaf_168_clk));
 sky130_fd_sc_hd__dfxtp_2 _42446_ (.D(_03332_),
    .Q(\cpuregs[16][21] ),
    .CLK(clknet_leaf_166_clk));
 sky130_fd_sc_hd__dfxtp_2 _42447_ (.D(_03333_),
    .Q(\cpuregs[16][22] ),
    .CLK(clknet_leaf_183_clk));
 sky130_fd_sc_hd__dfxtp_2 _42448_ (.D(_03334_),
    .Q(\cpuregs[16][23] ),
    .CLK(clknet_leaf_167_clk));
 sky130_fd_sc_hd__dfxtp_2 _42449_ (.D(_03335_),
    .Q(\cpuregs[16][24] ),
    .CLK(clknet_leaf_175_clk));
 sky130_fd_sc_hd__dfxtp_2 _42450_ (.D(_03336_),
    .Q(\cpuregs[16][25] ),
    .CLK(clknet_leaf_168_clk));
 sky130_fd_sc_hd__dfxtp_2 _42451_ (.D(_03337_),
    .Q(\cpuregs[16][26] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__dfxtp_2 _42452_ (.D(_03338_),
    .Q(\cpuregs[16][27] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__dfxtp_2 _42453_ (.D(_03339_),
    .Q(\cpuregs[16][28] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__dfxtp_2 _42454_ (.D(_03340_),
    .Q(\cpuregs[16][29] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__dfxtp_2 _42455_ (.D(_03341_),
    .Q(\cpuregs[16][30] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__dfxtp_2 _42456_ (.D(_03342_),
    .Q(\cpuregs[16][31] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__dfxtp_2 _42457_ (.D(_03343_),
    .Q(\cpuregs[12][0] ),
    .CLK(clknet_leaf_243_clk));
 sky130_fd_sc_hd__dfxtp_2 _42458_ (.D(_03344_),
    .Q(\cpuregs[12][1] ),
    .CLK(clknet_leaf_241_clk));
 sky130_fd_sc_hd__dfxtp_2 _42459_ (.D(_03345_),
    .Q(\cpuregs[12][2] ),
    .CLK(clknet_leaf_138_clk));
 sky130_fd_sc_hd__dfxtp_2 _42460_ (.D(_03346_),
    .Q(\cpuregs[12][3] ),
    .CLK(clknet_leaf_145_clk));
 sky130_fd_sc_hd__dfxtp_2 _42461_ (.D(_03347_),
    .Q(\cpuregs[12][4] ),
    .CLK(clknet_leaf_128_clk));
 sky130_fd_sc_hd__dfxtp_2 _42462_ (.D(_03348_),
    .Q(\cpuregs[12][5] ),
    .CLK(clknet_leaf_129_clk));
 sky130_fd_sc_hd__dfxtp_2 _42463_ (.D(_03349_),
    .Q(\cpuregs[12][6] ),
    .CLK(clknet_leaf_133_clk));
 sky130_fd_sc_hd__dfxtp_2 _42464_ (.D(_03350_),
    .Q(\cpuregs[12][7] ),
    .CLK(clknet_leaf_142_clk));
 sky130_fd_sc_hd__dfxtp_2 _42465_ (.D(_03351_),
    .Q(\cpuregs[12][8] ),
    .CLK(clknet_leaf_153_clk));
 sky130_fd_sc_hd__dfxtp_2 _42466_ (.D(_03352_),
    .Q(\cpuregs[12][9] ),
    .CLK(clknet_leaf_151_clk));
 sky130_fd_sc_hd__dfxtp_2 _42467_ (.D(_03353_),
    .Q(\cpuregs[12][10] ),
    .CLK(clknet_leaf_150_clk));
 sky130_fd_sc_hd__dfxtp_2 _42468_ (.D(_03354_),
    .Q(\cpuregs[12][11] ),
    .CLK(clknet_leaf_154_clk));
 sky130_fd_sc_hd__dfxtp_2 _42469_ (.D(_03355_),
    .Q(\cpuregs[12][12] ),
    .CLK(clknet_leaf_157_clk));
 sky130_fd_sc_hd__dfxtp_2 _42470_ (.D(_03356_),
    .Q(\cpuregs[12][13] ),
    .CLK(clknet_leaf_155_clk));
 sky130_fd_sc_hd__dfxtp_2 _42471_ (.D(_03357_),
    .Q(\cpuregs[12][14] ),
    .CLK(clknet_leaf_262_clk));
 sky130_fd_sc_hd__dfxtp_2 _42472_ (.D(_03358_),
    .Q(\cpuregs[12][15] ),
    .CLK(clknet_leaf_262_clk));
 sky130_fd_sc_hd__dfxtp_2 _42473_ (.D(_03359_),
    .Q(\cpuregs[12][16] ),
    .CLK(clknet_leaf_265_clk));
 sky130_fd_sc_hd__dfxtp_2 _42474_ (.D(_03360_),
    .Q(\cpuregs[12][17] ),
    .CLK(clknet_leaf_257_clk));
 sky130_fd_sc_hd__dfxtp_2 _42475_ (.D(_03361_),
    .Q(\cpuregs[12][18] ),
    .CLK(clknet_leaf_268_clk));
 sky130_fd_sc_hd__dfxtp_2 _42476_ (.D(_03362_),
    .Q(\cpuregs[12][19] ),
    .CLK(clknet_leaf_269_clk));
 sky130_fd_sc_hd__dfxtp_2 _42477_ (.D(_03363_),
    .Q(\cpuregs[12][20] ),
    .CLK(clknet_leaf_171_clk));
 sky130_fd_sc_hd__dfxtp_2 _42478_ (.D(_03364_),
    .Q(\cpuregs[12][21] ),
    .CLK(clknet_leaf_177_clk));
 sky130_fd_sc_hd__dfxtp_2 _42479_ (.D(_03365_),
    .Q(\cpuregs[12][22] ),
    .CLK(clknet_leaf_176_clk));
 sky130_fd_sc_hd__dfxtp_2 _42480_ (.D(_03366_),
    .Q(\cpuregs[12][23] ),
    .CLK(clknet_leaf_174_clk));
 sky130_fd_sc_hd__dfxtp_2 _42481_ (.D(_03367_),
    .Q(\cpuregs[12][24] ),
    .CLK(clknet_leaf_179_clk));
 sky130_fd_sc_hd__dfxtp_2 _42482_ (.D(_03368_),
    .Q(\cpuregs[12][25] ),
    .CLK(clknet_leaf_169_clk));
 sky130_fd_sc_hd__dfxtp_2 _42483_ (.D(_03369_),
    .Q(\cpuregs[12][26] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__dfxtp_2 _42484_ (.D(_03370_),
    .Q(\cpuregs[12][27] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__dfxtp_2 _42485_ (.D(_03371_),
    .Q(\cpuregs[12][28] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__dfxtp_2 _42486_ (.D(_03372_),
    .Q(\cpuregs[12][29] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__dfxtp_2 _42487_ (.D(_03373_),
    .Q(\cpuregs[12][30] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__dfxtp_2 _42488_ (.D(_03374_),
    .Q(\cpuregs[12][31] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__dfxtp_2 _42489_ (.D(_03375_),
    .Q(\cpuregs[1][0] ),
    .CLK(clknet_leaf_257_clk));
 sky130_fd_sc_hd__dfxtp_2 _42490_ (.D(_03376_),
    .Q(\cpuregs[1][1] ),
    .CLK(clknet_leaf_243_clk));
 sky130_fd_sc_hd__dfxtp_2 _42491_ (.D(_03377_),
    .Q(\cpuregs[1][2] ),
    .CLK(clknet_leaf_138_clk));
 sky130_fd_sc_hd__dfxtp_2 _42492_ (.D(_03378_),
    .Q(\cpuregs[1][3] ),
    .CLK(clknet_leaf_145_clk));
 sky130_fd_sc_hd__dfxtp_2 _42493_ (.D(_03379_),
    .Q(\cpuregs[1][4] ),
    .CLK(clknet_leaf_130_clk));
 sky130_fd_sc_hd__dfxtp_2 _42494_ (.D(_03380_),
    .Q(\cpuregs[1][5] ),
    .CLK(clknet_leaf_130_clk));
 sky130_fd_sc_hd__dfxtp_2 _42495_ (.D(_03381_),
    .Q(\cpuregs[1][6] ),
    .CLK(clknet_leaf_132_clk));
 sky130_fd_sc_hd__dfxtp_2 _42496_ (.D(_03382_),
    .Q(\cpuregs[1][7] ),
    .CLK(clknet_leaf_142_clk));
 sky130_fd_sc_hd__dfxtp_2 _42497_ (.D(_03383_),
    .Q(\cpuregs[1][8] ),
    .CLK(clknet_leaf_153_clk));
 sky130_fd_sc_hd__dfxtp_2 _42498_ (.D(_03384_),
    .Q(\cpuregs[1][9] ),
    .CLK(clknet_leaf_147_clk));
 sky130_fd_sc_hd__dfxtp_2 _42499_ (.D(_03385_),
    .Q(\cpuregs[1][10] ),
    .CLK(clknet_leaf_147_clk));
 sky130_fd_sc_hd__dfxtp_2 _42500_ (.D(_03386_),
    .Q(\cpuregs[1][11] ),
    .CLK(clknet_leaf_151_clk));
 sky130_fd_sc_hd__dfxtp_2 _42501_ (.D(_03387_),
    .Q(\cpuregs[1][12] ),
    .CLK(clknet_leaf_157_clk));
 sky130_fd_sc_hd__dfxtp_2 _42502_ (.D(_03388_),
    .Q(\cpuregs[1][13] ),
    .CLK(clknet_leaf_159_clk));
 sky130_fd_sc_hd__dfxtp_2 _42503_ (.D(_03389_),
    .Q(\cpuregs[1][14] ),
    .CLK(clknet_leaf_266_clk));
 sky130_fd_sc_hd__dfxtp_2 _42504_ (.D(_03390_),
    .Q(\cpuregs[1][15] ),
    .CLK(clknet_leaf_262_clk));
 sky130_fd_sc_hd__dfxtp_2 _42505_ (.D(_03391_),
    .Q(\cpuregs[1][16] ),
    .CLK(clknet_leaf_265_clk));
 sky130_fd_sc_hd__dfxtp_2 _42506_ (.D(_03392_),
    .Q(\cpuregs[1][17] ),
    .CLK(clknet_leaf_262_clk));
 sky130_fd_sc_hd__dfxtp_2 _42507_ (.D(_03393_),
    .Q(\cpuregs[1][18] ),
    .CLK(clknet_leaf_269_clk));
 sky130_fd_sc_hd__dfxtp_2 _42508_ (.D(_03394_),
    .Q(\cpuregs[1][19] ),
    .CLK(clknet_leaf_269_clk));
 sky130_fd_sc_hd__dfxtp_2 _42509_ (.D(_03395_),
    .Q(\cpuregs[1][20] ),
    .CLK(clknet_leaf_156_clk));
 sky130_fd_sc_hd__dfxtp_2 _42510_ (.D(_03396_),
    .Q(\cpuregs[1][21] ),
    .CLK(clknet_leaf_173_clk));
 sky130_fd_sc_hd__dfxtp_2 _42511_ (.D(_03397_),
    .Q(\cpuregs[1][22] ),
    .CLK(clknet_leaf_181_clk));
 sky130_fd_sc_hd__dfxtp_2 _42512_ (.D(_03398_),
    .Q(\cpuregs[1][23] ),
    .CLK(clknet_leaf_174_clk));
 sky130_fd_sc_hd__dfxtp_2 _42513_ (.D(_03399_),
    .Q(\cpuregs[1][24] ),
    .CLK(clknet_leaf_179_clk));
 sky130_fd_sc_hd__dfxtp_2 _42514_ (.D(_03400_),
    .Q(\cpuregs[1][25] ),
    .CLK(clknet_leaf_157_clk));
 sky130_fd_sc_hd__dfxtp_2 _42515_ (.D(_03401_),
    .Q(\cpuregs[1][26] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__dfxtp_2 _42516_ (.D(_03402_),
    .Q(\cpuregs[1][27] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfxtp_2 _42517_ (.D(_03403_),
    .Q(\cpuregs[1][28] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__dfxtp_2 _42518_ (.D(_03404_),
    .Q(\cpuregs[1][29] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__dfxtp_2 _42519_ (.D(_03405_),
    .Q(\cpuregs[1][30] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__dfxtp_2 _42520_ (.D(_03406_),
    .Q(\cpuregs[1][31] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfxtp_2 _42521_ (.D(_03407_),
    .Q(\cpuregs[3][0] ),
    .CLK(clknet_leaf_258_clk));
 sky130_fd_sc_hd__dfxtp_2 _42522_ (.D(_03408_),
    .Q(\cpuregs[3][1] ),
    .CLK(clknet_leaf_243_clk));
 sky130_fd_sc_hd__dfxtp_2 _42523_ (.D(_03409_),
    .Q(\cpuregs[3][2] ),
    .CLK(clknet_leaf_138_clk));
 sky130_fd_sc_hd__dfxtp_2 _42524_ (.D(_03410_),
    .Q(\cpuregs[3][3] ),
    .CLK(clknet_leaf_145_clk));
 sky130_fd_sc_hd__dfxtp_2 _42525_ (.D(_03411_),
    .Q(\cpuregs[3][4] ),
    .CLK(clknet_leaf_130_clk));
 sky130_fd_sc_hd__dfxtp_2 _42526_ (.D(_03412_),
    .Q(\cpuregs[3][5] ),
    .CLK(clknet_leaf_130_clk));
 sky130_fd_sc_hd__dfxtp_2 _42527_ (.D(_03413_),
    .Q(\cpuregs[3][6] ),
    .CLK(clknet_leaf_131_clk));
 sky130_fd_sc_hd__dfxtp_2 _42528_ (.D(_03414_),
    .Q(\cpuregs[3][7] ),
    .CLK(clknet_leaf_127_clk));
 sky130_fd_sc_hd__dfxtp_2 _42529_ (.D(_03415_),
    .Q(\cpuregs[3][8] ),
    .CLK(clknet_leaf_153_clk));
 sky130_fd_sc_hd__dfxtp_2 _42530_ (.D(_03416_),
    .Q(\cpuregs[3][9] ),
    .CLK(clknet_leaf_148_clk));
 sky130_fd_sc_hd__dfxtp_2 _42531_ (.D(_03417_),
    .Q(\cpuregs[3][10] ),
    .CLK(clknet_leaf_148_clk));
 sky130_fd_sc_hd__dfxtp_2 _42532_ (.D(_03418_),
    .Q(\cpuregs[3][11] ),
    .CLK(clknet_leaf_151_clk));
 sky130_fd_sc_hd__dfxtp_2 _42533_ (.D(_03419_),
    .Q(\cpuregs[3][12] ),
    .CLK(clknet_leaf_157_clk));
 sky130_fd_sc_hd__dfxtp_2 _42534_ (.D(_03420_),
    .Q(\cpuregs[3][13] ),
    .CLK(clknet_leaf_159_clk));
 sky130_fd_sc_hd__dfxtp_2 _42535_ (.D(_03421_),
    .Q(\cpuregs[3][14] ),
    .CLK(clknet_leaf_261_clk));
 sky130_fd_sc_hd__dfxtp_2 _42536_ (.D(_03422_),
    .Q(\cpuregs[3][15] ),
    .CLK(clknet_leaf_260_clk));
 sky130_fd_sc_hd__dfxtp_2 _42537_ (.D(_03423_),
    .Q(\cpuregs[3][16] ),
    .CLK(clknet_leaf_266_clk));
 sky130_fd_sc_hd__dfxtp_2 _42538_ (.D(_03424_),
    .Q(\cpuregs[3][17] ),
    .CLK(clknet_leaf_259_clk));
 sky130_fd_sc_hd__dfxtp_2 _42539_ (.D(_03425_),
    .Q(\cpuregs[3][18] ),
    .CLK(clknet_leaf_268_clk));
 sky130_fd_sc_hd__dfxtp_2 _42540_ (.D(_03426_),
    .Q(\cpuregs[3][19] ),
    .CLK(clknet_leaf_269_clk));
 sky130_fd_sc_hd__dfxtp_2 _42541_ (.D(_03427_),
    .Q(\cpuregs[3][20] ),
    .CLK(clknet_leaf_156_clk));
 sky130_fd_sc_hd__dfxtp_2 _42542_ (.D(_03428_),
    .Q(\cpuregs[3][21] ),
    .CLK(clknet_leaf_173_clk));
 sky130_fd_sc_hd__dfxtp_2 _42543_ (.D(_03429_),
    .Q(\cpuregs[3][22] ),
    .CLK(clknet_leaf_181_clk));
 sky130_fd_sc_hd__dfxtp_2 _42544_ (.D(_03430_),
    .Q(\cpuregs[3][23] ),
    .CLK(clknet_leaf_172_clk));
 sky130_fd_sc_hd__dfxtp_2 _42545_ (.D(_03431_),
    .Q(\cpuregs[3][24] ),
    .CLK(clknet_leaf_179_clk));
 sky130_fd_sc_hd__dfxtp_2 _42546_ (.D(_03432_),
    .Q(\cpuregs[3][25] ),
    .CLK(clknet_leaf_156_clk));
 sky130_fd_sc_hd__dfxtp_2 _42547_ (.D(_03433_),
    .Q(\cpuregs[3][26] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__dfxtp_2 _42548_ (.D(_03434_),
    .Q(\cpuregs[3][27] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfxtp_2 _42549_ (.D(_03435_),
    .Q(\cpuregs[3][28] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__dfxtp_2 _42550_ (.D(_03436_),
    .Q(\cpuregs[3][29] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__dfxtp_2 _42551_ (.D(_03437_),
    .Q(\cpuregs[3][30] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__dfxtp_2 _42552_ (.D(_03438_),
    .Q(\cpuregs[3][31] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfxtp_2 _42553_ (.D(_03439_),
    .Q(\cpuregs[11][0] ),
    .CLK(clknet_leaf_242_clk));
 sky130_fd_sc_hd__dfxtp_2 _42554_ (.D(_03440_),
    .Q(\cpuregs[11][1] ),
    .CLK(clknet_leaf_241_clk));
 sky130_fd_sc_hd__dfxtp_2 _42555_ (.D(_03441_),
    .Q(\cpuregs[11][2] ),
    .CLK(clknet_leaf_141_clk));
 sky130_fd_sc_hd__dfxtp_2 _42556_ (.D(_03442_),
    .Q(\cpuregs[11][3] ),
    .CLK(clknet_leaf_143_clk));
 sky130_fd_sc_hd__dfxtp_2 _42557_ (.D(_03443_),
    .Q(\cpuregs[11][4] ),
    .CLK(clknet_leaf_126_clk));
 sky130_fd_sc_hd__dfxtp_2 _42558_ (.D(_03444_),
    .Q(\cpuregs[11][5] ),
    .CLK(clknet_leaf_130_clk));
 sky130_fd_sc_hd__dfxtp_2 _42559_ (.D(_03445_),
    .Q(\cpuregs[11][6] ),
    .CLK(clknet_leaf_131_clk));
 sky130_fd_sc_hd__dfxtp_2 _42560_ (.D(_03446_),
    .Q(\cpuregs[11][7] ),
    .CLK(clknet_leaf_142_clk));
 sky130_fd_sc_hd__dfxtp_2 _42561_ (.D(_03447_),
    .Q(\cpuregs[11][8] ),
    .CLK(clknet_leaf_160_clk));
 sky130_fd_sc_hd__dfxtp_2 _42562_ (.D(_03448_),
    .Q(\cpuregs[11][9] ),
    .CLK(clknet_leaf_147_clk));
 sky130_fd_sc_hd__dfxtp_2 _42563_ (.D(_03449_),
    .Q(\cpuregs[11][10] ),
    .CLK(clknet_leaf_147_clk));
 sky130_fd_sc_hd__dfxtp_2 _42564_ (.D(_03450_),
    .Q(\cpuregs[11][11] ),
    .CLK(clknet_leaf_152_clk));
 sky130_fd_sc_hd__dfxtp_2 _42565_ (.D(_03451_),
    .Q(\cpuregs[11][12] ),
    .CLK(clknet_leaf_158_clk));
 sky130_fd_sc_hd__dfxtp_2 _42566_ (.D(_03452_),
    .Q(\cpuregs[11][13] ),
    .CLK(clknet_leaf_159_clk));
 sky130_fd_sc_hd__dfxtp_2 _42567_ (.D(_03453_),
    .Q(\cpuregs[11][14] ),
    .CLK(clknet_leaf_263_clk));
 sky130_fd_sc_hd__dfxtp_2 _42568_ (.D(_03454_),
    .Q(\cpuregs[11][15] ),
    .CLK(clknet_leaf_255_clk));
 sky130_fd_sc_hd__dfxtp_2 _42569_ (.D(_03455_),
    .Q(\cpuregs[11][16] ),
    .CLK(clknet_leaf_264_clk));
 sky130_fd_sc_hd__dfxtp_2 _42570_ (.D(_03456_),
    .Q(\cpuregs[11][17] ),
    .CLK(clknet_leaf_255_clk));
 sky130_fd_sc_hd__dfxtp_2 _42571_ (.D(_03457_),
    .Q(\cpuregs[11][18] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__dfxtp_2 _42572_ (.D(_03458_),
    .Q(\cpuregs[11][19] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__dfxtp_2 _42573_ (.D(_03459_),
    .Q(\cpuregs[11][20] ),
    .CLK(clknet_leaf_156_clk));
 sky130_fd_sc_hd__dfxtp_2 _42574_ (.D(_03460_),
    .Q(\cpuregs[11][21] ),
    .CLK(clknet_leaf_174_clk));
 sky130_fd_sc_hd__dfxtp_2 _42575_ (.D(_03461_),
    .Q(\cpuregs[11][22] ),
    .CLK(clknet_leaf_177_clk));
 sky130_fd_sc_hd__dfxtp_2 _42576_ (.D(_03462_),
    .Q(\cpuregs[11][23] ),
    .CLK(clknet_leaf_174_clk));
 sky130_fd_sc_hd__dfxtp_2 _42577_ (.D(_03463_),
    .Q(\cpuregs[11][24] ),
    .CLK(clknet_leaf_177_clk));
 sky130_fd_sc_hd__dfxtp_2 _42578_ (.D(_03464_),
    .Q(\cpuregs[11][25] ),
    .CLK(clknet_leaf_169_clk));
 sky130_fd_sc_hd__dfxtp_2 _42579_ (.D(_03465_),
    .Q(\cpuregs[11][26] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__dfxtp_2 _42580_ (.D(_03466_),
    .Q(\cpuregs[11][27] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__dfxtp_2 _42581_ (.D(_03467_),
    .Q(\cpuregs[11][28] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__dfxtp_2 _42582_ (.D(_03468_),
    .Q(\cpuregs[11][29] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__dfxtp_2 _42583_ (.D(_03469_),
    .Q(\cpuregs[11][30] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__dfxtp_2 _42584_ (.D(_03470_),
    .Q(\cpuregs[11][31] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__dfxtp_2 _42585_ (.D(_03471_),
    .Q(\cpuregs[15][0] ),
    .CLK(clknet_leaf_243_clk));
 sky130_fd_sc_hd__dfxtp_2 _42586_ (.D(_03472_),
    .Q(\cpuregs[15][1] ),
    .CLK(clknet_leaf_240_clk));
 sky130_fd_sc_hd__dfxtp_2 _42587_ (.D(_03473_),
    .Q(\cpuregs[15][2] ),
    .CLK(clknet_leaf_139_clk));
 sky130_fd_sc_hd__dfxtp_2 _42588_ (.D(_03474_),
    .Q(\cpuregs[15][3] ),
    .CLK(clknet_leaf_145_clk));
 sky130_fd_sc_hd__dfxtp_2 _42589_ (.D(_03475_),
    .Q(\cpuregs[15][4] ),
    .CLK(clknet_leaf_127_clk));
 sky130_fd_sc_hd__dfxtp_2 _42590_ (.D(_03476_),
    .Q(\cpuregs[15][5] ),
    .CLK(clknet_leaf_128_clk));
 sky130_fd_sc_hd__dfxtp_2 _42591_ (.D(_03477_),
    .Q(\cpuregs[15][6] ),
    .CLK(clknet_leaf_133_clk));
 sky130_fd_sc_hd__dfxtp_2 _42592_ (.D(_03478_),
    .Q(\cpuregs[15][7] ),
    .CLK(clknet_leaf_142_clk));
 sky130_fd_sc_hd__dfxtp_2 _42593_ (.D(_03479_),
    .Q(\cpuregs[15][8] ),
    .CLK(clknet_leaf_152_clk));
 sky130_fd_sc_hd__dfxtp_2 _42594_ (.D(_03480_),
    .Q(\cpuregs[15][9] ),
    .CLK(clknet_leaf_151_clk));
 sky130_fd_sc_hd__dfxtp_2 _42595_ (.D(_03481_),
    .Q(\cpuregs[15][10] ),
    .CLK(clknet_leaf_150_clk));
 sky130_fd_sc_hd__dfxtp_2 _42596_ (.D(_03482_),
    .Q(\cpuregs[15][11] ),
    .CLK(clknet_leaf_152_clk));
 sky130_fd_sc_hd__dfxtp_2 _42597_ (.D(_03483_),
    .Q(\cpuregs[15][12] ),
    .CLK(clknet_leaf_157_clk));
 sky130_fd_sc_hd__dfxtp_2 _42598_ (.D(_03484_),
    .Q(\cpuregs[15][13] ),
    .CLK(clknet_leaf_153_clk));
 sky130_fd_sc_hd__dfxtp_2 _42599_ (.D(_03485_),
    .Q(\cpuregs[15][14] ),
    .CLK(clknet_leaf_262_clk));
 sky130_fd_sc_hd__dfxtp_2 _42600_ (.D(_03486_),
    .Q(\cpuregs[15][15] ),
    .CLK(clknet_leaf_260_clk));
 sky130_fd_sc_hd__dfxtp_2 _42601_ (.D(_03487_),
    .Q(\cpuregs[15][16] ),
    .CLK(clknet_leaf_265_clk));
 sky130_fd_sc_hd__dfxtp_2 _42602_ (.D(_03488_),
    .Q(\cpuregs[15][17] ),
    .CLK(clknet_leaf_257_clk));
 sky130_fd_sc_hd__dfxtp_2 _42603_ (.D(_03489_),
    .Q(\cpuregs[15][18] ),
    .CLK(clknet_leaf_265_clk));
 sky130_fd_sc_hd__dfxtp_2 _42604_ (.D(_03490_),
    .Q(\cpuregs[15][19] ),
    .CLK(clknet_leaf_265_clk));
 sky130_fd_sc_hd__dfxtp_2 _42605_ (.D(_03491_),
    .Q(\cpuregs[15][20] ),
    .CLK(clknet_leaf_171_clk));
 sky130_fd_sc_hd__dfxtp_2 _42606_ (.D(_03492_),
    .Q(\cpuregs[15][21] ),
    .CLK(clknet_leaf_177_clk));
 sky130_fd_sc_hd__dfxtp_2 _42607_ (.D(_03493_),
    .Q(\cpuregs[15][22] ),
    .CLK(clknet_leaf_176_clk));
 sky130_fd_sc_hd__dfxtp_2 _42608_ (.D(_03494_),
    .Q(\cpuregs[15][23] ),
    .CLK(clknet_leaf_171_clk));
 sky130_fd_sc_hd__dfxtp_2 _42609_ (.D(_03495_),
    .Q(\cpuregs[15][24] ),
    .CLK(clknet_leaf_176_clk));
 sky130_fd_sc_hd__dfxtp_2 _42610_ (.D(_03496_),
    .Q(\cpuregs[15][25] ),
    .CLK(clknet_leaf_169_clk));
 sky130_fd_sc_hd__dfxtp_2 _42611_ (.D(_03497_),
    .Q(\cpuregs[15][26] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__dfxtp_2 _42612_ (.D(_03498_),
    .Q(\cpuregs[15][27] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__dfxtp_2 _42613_ (.D(_03499_),
    .Q(\cpuregs[15][28] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__dfxtp_2 _42614_ (.D(_03500_),
    .Q(\cpuregs[15][29] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__dfxtp_2 _42615_ (.D(_03501_),
    .Q(\cpuregs[15][30] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__dfxtp_2 _42616_ (.D(_03502_),
    .Q(\cpuregs[15][31] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__dfxtp_2 _42617_ (.D(_03503_),
    .Q(\latched_rd[4] ),
    .CLK(clknet_leaf_221_clk));
 sky130_fd_sc_hd__dfxtp_2 _42618_ (.D(_03504_),
    .Q(\cpuregs[7][0] ),
    .CLK(clknet_leaf_242_clk));
 sky130_fd_sc_hd__dfxtp_2 _42619_ (.D(_03505_),
    .Q(\cpuregs[7][1] ),
    .CLK(clknet_leaf_241_clk));
 sky130_fd_sc_hd__dfxtp_2 _42620_ (.D(_03506_),
    .Q(\cpuregs[7][2] ),
    .CLK(clknet_leaf_139_clk));
 sky130_fd_sc_hd__dfxtp_2 _42621_ (.D(_03507_),
    .Q(\cpuregs[7][3] ),
    .CLK(clknet_leaf_144_clk));
 sky130_fd_sc_hd__dfxtp_2 _42622_ (.D(_03508_),
    .Q(\cpuregs[7][4] ),
    .CLK(clknet_leaf_127_clk));
 sky130_fd_sc_hd__dfxtp_2 _42623_ (.D(_03509_),
    .Q(\cpuregs[7][5] ),
    .CLK(clknet_leaf_129_clk));
 sky130_fd_sc_hd__dfxtp_2 _42624_ (.D(_03510_),
    .Q(\cpuregs[7][6] ),
    .CLK(clknet_leaf_133_clk));
 sky130_fd_sc_hd__dfxtp_2 _42625_ (.D(_03511_),
    .Q(\cpuregs[7][7] ),
    .CLK(clknet_leaf_143_clk));
 sky130_fd_sc_hd__dfxtp_2 _42626_ (.D(_03512_),
    .Q(\cpuregs[7][8] ),
    .CLK(clknet_leaf_155_clk));
 sky130_fd_sc_hd__dfxtp_2 _42627_ (.D(_03513_),
    .Q(\cpuregs[7][9] ),
    .CLK(clknet_leaf_150_clk));
 sky130_fd_sc_hd__dfxtp_2 _42628_ (.D(_03514_),
    .Q(\cpuregs[7][10] ),
    .CLK(clknet_leaf_150_clk));
 sky130_fd_sc_hd__dfxtp_2 _42629_ (.D(_03515_),
    .Q(\cpuregs[7][11] ),
    .CLK(clknet_leaf_150_clk));
 sky130_fd_sc_hd__dfxtp_2 _42630_ (.D(_03516_),
    .Q(\cpuregs[7][12] ),
    .CLK(clknet_leaf_155_clk));
 sky130_fd_sc_hd__dfxtp_2 _42631_ (.D(_03517_),
    .Q(\cpuregs[7][13] ),
    .CLK(clknet_leaf_155_clk));
 sky130_fd_sc_hd__dfxtp_2 _42632_ (.D(_03518_),
    .Q(\cpuregs[7][14] ),
    .CLK(clknet_leaf_261_clk));
 sky130_fd_sc_hd__dfxtp_2 _42633_ (.D(_03519_),
    .Q(\cpuregs[7][15] ),
    .CLK(clknet_leaf_260_clk));
 sky130_fd_sc_hd__dfxtp_2 _42634_ (.D(_03520_),
    .Q(\cpuregs[7][16] ),
    .CLK(clknet_leaf_266_clk));
 sky130_fd_sc_hd__dfxtp_2 _42635_ (.D(_03521_),
    .Q(\cpuregs[7][17] ),
    .CLK(clknet_leaf_259_clk));
 sky130_fd_sc_hd__dfxtp_2 _42636_ (.D(_03522_),
    .Q(\cpuregs[7][18] ),
    .CLK(clknet_leaf_267_clk));
 sky130_fd_sc_hd__dfxtp_2 _42637_ (.D(_03523_),
    .Q(\cpuregs[7][19] ),
    .CLK(clknet_leaf_267_clk));
 sky130_fd_sc_hd__dfxtp_2 _42638_ (.D(_03524_),
    .Q(\cpuregs[7][20] ),
    .CLK(clknet_leaf_170_clk));
 sky130_fd_sc_hd__dfxtp_2 _42639_ (.D(_03525_),
    .Q(\cpuregs[7][21] ),
    .CLK(clknet_leaf_173_clk));
 sky130_fd_sc_hd__dfxtp_2 _42640_ (.D(_03526_),
    .Q(\cpuregs[7][22] ),
    .CLK(clknet_leaf_178_clk));
 sky130_fd_sc_hd__dfxtp_2 _42641_ (.D(_03527_),
    .Q(\cpuregs[7][23] ),
    .CLK(clknet_leaf_172_clk));
 sky130_fd_sc_hd__dfxtp_2 _42642_ (.D(_03528_),
    .Q(\cpuregs[7][24] ),
    .CLK(clknet_leaf_178_clk));
 sky130_fd_sc_hd__dfxtp_2 _42643_ (.D(_03529_),
    .Q(\cpuregs[7][25] ),
    .CLK(clknet_leaf_170_clk));
 sky130_fd_sc_hd__dfxtp_2 _42644_ (.D(_03530_),
    .Q(\cpuregs[7][26] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__dfxtp_2 _42645_ (.D(_03531_),
    .Q(\cpuregs[7][27] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__dfxtp_2 _42646_ (.D(_03532_),
    .Q(\cpuregs[7][28] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__dfxtp_2 _42647_ (.D(_03533_),
    .Q(\cpuregs[7][29] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__dfxtp_2 _42648_ (.D(_03534_),
    .Q(\cpuregs[7][30] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__dfxtp_2 _42649_ (.D(_03535_),
    .Q(\cpuregs[7][31] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__dfxtp_2 _42650_ (.D(_03536_),
    .Q(mem_wdata[0]),
    .CLK(clknet_leaf_207_clk));
 sky130_fd_sc_hd__dfxtp_2 _42651_ (.D(_03537_),
    .Q(mem_wdata[1]),
    .CLK(clknet_leaf_207_clk));
 sky130_fd_sc_hd__dfxtp_2 _42652_ (.D(_03538_),
    .Q(mem_wdata[2]),
    .CLK(clknet_leaf_123_clk));
 sky130_fd_sc_hd__dfxtp_2 _42653_ (.D(_03539_),
    .Q(mem_wdata[3]),
    .CLK(clknet_leaf_208_clk));
 sky130_fd_sc_hd__dfxtp_2 _42654_ (.D(_03540_),
    .Q(mem_wdata[4]),
    .CLK(clknet_leaf_131_clk));
 sky130_fd_sc_hd__dfxtp_2 _42655_ (.D(_03541_),
    .Q(mem_wdata[5]),
    .CLK(clknet_leaf_208_clk));
 sky130_fd_sc_hd__dfxtp_2 _42656_ (.D(_03542_),
    .Q(mem_wdata[6]),
    .CLK(clknet_leaf_131_clk));
 sky130_fd_sc_hd__dfxtp_2 _42657_ (.D(_03543_),
    .Q(mem_wdata[7]),
    .CLK(clknet_leaf_123_clk));
 sky130_fd_sc_hd__dfxtp_2 _42658_ (.D(_03544_),
    .Q(mem_wdata[8]),
    .CLK(clknet_leaf_180_clk));
 sky130_fd_sc_hd__dfxtp_2 _42659_ (.D(_03545_),
    .Q(mem_wdata[9]),
    .CLK(clknet_leaf_179_clk));
 sky130_fd_sc_hd__dfxtp_2 _42660_ (.D(_03546_),
    .Q(mem_wdata[10]),
    .CLK(clknet_leaf_95_clk));
 sky130_fd_sc_hd__dfxtp_2 _42661_ (.D(_03547_),
    .Q(mem_wdata[11]),
    .CLK(clknet_leaf_95_clk));
 sky130_fd_sc_hd__dfxtp_2 _42662_ (.D(_03548_),
    .Q(mem_wdata[12]),
    .CLK(clknet_opt_1_clk));
 sky130_fd_sc_hd__dfxtp_2 _42663_ (.D(_03549_),
    .Q(mem_wdata[13]),
    .CLK(clknet_leaf_180_clk));
 sky130_fd_sc_hd__dfxtp_2 _42664_ (.D(_03550_),
    .Q(mem_wdata[14]),
    .CLK(clknet_leaf_95_clk));
 sky130_fd_sc_hd__dfxtp_2 _42665_ (.D(_03551_),
    .Q(mem_wdata[15]),
    .CLK(clknet_leaf_121_clk));
 sky130_fd_sc_hd__dfxtp_2 _42666_ (.D(_03552_),
    .Q(mem_wdata[16]),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__dfxtp_2 _42667_ (.D(_03553_),
    .Q(mem_wdata[17]),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__dfxtp_2 _42668_ (.D(_03554_),
    .Q(mem_wdata[18]),
    .CLK(clknet_leaf_205_clk));
 sky130_fd_sc_hd__dfxtp_2 _42669_ (.D(_03555_),
    .Q(mem_wdata[19]),
    .CLK(clknet_leaf_121_clk));
 sky130_fd_sc_hd__dfxtp_2 _42670_ (.D(_03556_),
    .Q(mem_wdata[20]),
    .CLK(clknet_opt_15_clk));
 sky130_fd_sc_hd__dfxtp_2 _42671_ (.D(_03557_),
    .Q(mem_wdata[21]),
    .CLK(clknet_leaf_109_clk));
 sky130_fd_sc_hd__dfxtp_2 _42672_ (.D(_03558_),
    .Q(mem_wdata[22]),
    .CLK(clknet_leaf_95_clk));
 sky130_fd_sc_hd__dfxtp_2 _42673_ (.D(_03559_),
    .Q(mem_wdata[23]),
    .CLK(clknet_leaf_95_clk));
 sky130_fd_sc_hd__dfxtp_2 _42674_ (.D(_03560_),
    .Q(mem_wdata[24]),
    .CLK(clknet_leaf_94_clk));
 sky130_fd_sc_hd__dfxtp_2 _42675_ (.D(_03561_),
    .Q(mem_wdata[25]),
    .CLK(clknet_leaf_95_clk));
 sky130_fd_sc_hd__dfxtp_2 _42676_ (.D(_03562_),
    .Q(mem_wdata[26]),
    .CLK(clknet_opt_14_clk));
 sky130_fd_sc_hd__dfxtp_2 _42677_ (.D(_03563_),
    .Q(mem_wdata[27]),
    .CLK(clknet_leaf_177_clk));
 sky130_fd_sc_hd__dfxtp_2 _42678_ (.D(_03564_),
    .Q(mem_wdata[28]),
    .CLK(clknet_opt_4_clk));
 sky130_fd_sc_hd__dfxtp_2 _42679_ (.D(_03565_),
    .Q(mem_wdata[29]),
    .CLK(clknet_leaf_109_clk));
 sky130_fd_sc_hd__dfxtp_2 _42680_ (.D(_03566_),
    .Q(mem_wdata[30]),
    .CLK(clknet_leaf_94_clk));
 sky130_fd_sc_hd__dfxtp_2 _42681_ (.D(_03567_),
    .Q(mem_wdata[31]),
    .CLK(clknet_opt_16_clk));
 sky130_fd_sc_hd__dfxtp_2 _42682_ (.D(_03568_),
    .Q(\cpuregs[19][0] ),
    .CLK(clknet_leaf_257_clk));
 sky130_fd_sc_hd__dfxtp_2 _42683_ (.D(_03569_),
    .Q(\cpuregs[19][1] ),
    .CLK(clknet_leaf_246_clk));
 sky130_fd_sc_hd__dfxtp_2 _42684_ (.D(_03570_),
    .Q(\cpuregs[19][2] ),
    .CLK(clknet_leaf_141_clk));
 sky130_fd_sc_hd__dfxtp_2 _42685_ (.D(_03571_),
    .Q(\cpuregs[19][3] ),
    .CLK(clknet_leaf_140_clk));
 sky130_fd_sc_hd__dfxtp_2 _42686_ (.D(_03572_),
    .Q(\cpuregs[19][4] ),
    .CLK(clknet_leaf_128_clk));
 sky130_fd_sc_hd__dfxtp_2 _42687_ (.D(_03573_),
    .Q(\cpuregs[19][5] ),
    .CLK(clknet_leaf_129_clk));
 sky130_fd_sc_hd__dfxtp_2 _42688_ (.D(_03574_),
    .Q(\cpuregs[19][6] ),
    .CLK(clknet_leaf_137_clk));
 sky130_fd_sc_hd__dfxtp_2 _42689_ (.D(_03575_),
    .Q(\cpuregs[19][7] ),
    .CLK(clknet_leaf_140_clk));
 sky130_fd_sc_hd__dfxtp_2 _42690_ (.D(_03576_),
    .Q(\cpuregs[19][8] ),
    .CLK(clknet_leaf_160_clk));
 sky130_fd_sc_hd__dfxtp_2 _42691_ (.D(_03577_),
    .Q(\cpuregs[19][9] ),
    .CLK(clknet_leaf_146_clk));
 sky130_fd_sc_hd__dfxtp_2 _42692_ (.D(_03578_),
    .Q(\cpuregs[19][10] ),
    .CLK(clknet_leaf_146_clk));
 sky130_fd_sc_hd__dfxtp_2 _42693_ (.D(_03579_),
    .Q(\cpuregs[19][11] ),
    .CLK(clknet_leaf_152_clk));
 sky130_fd_sc_hd__dfxtp_2 _42694_ (.D(_03580_),
    .Q(\cpuregs[19][12] ),
    .CLK(clknet_leaf_158_clk));
 sky130_fd_sc_hd__dfxtp_2 _42695_ (.D(_03581_),
    .Q(\cpuregs[19][13] ),
    .CLK(clknet_leaf_160_clk));
 sky130_fd_sc_hd__dfxtp_2 _42696_ (.D(_03582_),
    .Q(\cpuregs[19][14] ),
    .CLK(clknet_leaf_263_clk));
 sky130_fd_sc_hd__dfxtp_2 _42697_ (.D(_03583_),
    .Q(\cpuregs[19][15] ),
    .CLK(clknet_leaf_263_clk));
 sky130_fd_sc_hd__dfxtp_2 _42698_ (.D(_03584_),
    .Q(\cpuregs[19][16] ),
    .CLK(clknet_leaf_264_clk));
 sky130_fd_sc_hd__dfxtp_2 _42699_ (.D(_03585_),
    .Q(\cpuregs[19][17] ),
    .CLK(clknet_leaf_255_clk));
 sky130_fd_sc_hd__dfxtp_2 _42700_ (.D(_03586_),
    .Q(\cpuregs[19][18] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__dfxtp_2 _42701_ (.D(_03587_),
    .Q(\cpuregs[19][19] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__dfxtp_2 _42702_ (.D(_03588_),
    .Q(\cpuregs[19][20] ),
    .CLK(clknet_leaf_168_clk));
 sky130_fd_sc_hd__dfxtp_2 _42703_ (.D(_03589_),
    .Q(\cpuregs[19][21] ),
    .CLK(clknet_leaf_175_clk));
 sky130_fd_sc_hd__dfxtp_2 _42704_ (.D(_03590_),
    .Q(\cpuregs[19][22] ),
    .CLK(clknet_leaf_176_clk));
 sky130_fd_sc_hd__dfxtp_2 _42705_ (.D(_03591_),
    .Q(\cpuregs[19][23] ),
    .CLK(clknet_leaf_167_clk));
 sky130_fd_sc_hd__dfxtp_2 _42706_ (.D(_03592_),
    .Q(\cpuregs[19][24] ),
    .CLK(clknet_leaf_175_clk));
 sky130_fd_sc_hd__dfxtp_2 _42707_ (.D(_03593_),
    .Q(\cpuregs[19][25] ),
    .CLK(clknet_leaf_168_clk));
 sky130_fd_sc_hd__dfxtp_2 _42708_ (.D(_03594_),
    .Q(\cpuregs[19][26] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__dfxtp_2 _42709_ (.D(_03595_),
    .Q(\cpuregs[19][27] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__dfxtp_2 _42710_ (.D(_03596_),
    .Q(\cpuregs[19][28] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__dfxtp_2 _42711_ (.D(_03597_),
    .Q(\cpuregs[19][29] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__dfxtp_2 _42712_ (.D(_03598_),
    .Q(\cpuregs[19][30] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__dfxtp_2 _42713_ (.D(_03599_),
    .Q(\cpuregs[19][31] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__dfxtp_2 _42714_ (.D(_03600_),
    .Q(\cpuregs[4][0] ),
    .CLK(clknet_leaf_258_clk));
 sky130_fd_sc_hd__dfxtp_2 _42715_ (.D(_03601_),
    .Q(\cpuregs[4][1] ),
    .CLK(clknet_leaf_242_clk));
 sky130_fd_sc_hd__dfxtp_2 _42716_ (.D(_03602_),
    .Q(\cpuregs[4][2] ),
    .CLK(clknet_leaf_140_clk));
 sky130_fd_sc_hd__dfxtp_2 _42717_ (.D(_03603_),
    .Q(\cpuregs[4][3] ),
    .CLK(clknet_leaf_144_clk));
 sky130_fd_sc_hd__dfxtp_2 _42718_ (.D(_03604_),
    .Q(\cpuregs[4][4] ),
    .CLK(clknet_leaf_127_clk));
 sky130_fd_sc_hd__dfxtp_2 _42719_ (.D(_03605_),
    .Q(\cpuregs[4][5] ),
    .CLK(clknet_leaf_129_clk));
 sky130_fd_sc_hd__dfxtp_2 _42720_ (.D(_03606_),
    .Q(\cpuregs[4][6] ),
    .CLK(clknet_leaf_132_clk));
 sky130_fd_sc_hd__dfxtp_2 _42721_ (.D(_03607_),
    .Q(\cpuregs[4][7] ),
    .CLK(clknet_leaf_143_clk));
 sky130_fd_sc_hd__dfxtp_2 _42722_ (.D(_03608_),
    .Q(\cpuregs[4][8] ),
    .CLK(clknet_leaf_155_clk));
 sky130_fd_sc_hd__dfxtp_2 _42723_ (.D(_03609_),
    .Q(\cpuregs[4][9] ),
    .CLK(clknet_leaf_150_clk));
 sky130_fd_sc_hd__dfxtp_2 _42724_ (.D(_03610_),
    .Q(\cpuregs[4][10] ),
    .CLK(clknet_leaf_150_clk));
 sky130_fd_sc_hd__dfxtp_2 _42725_ (.D(_03611_),
    .Q(\cpuregs[4][11] ),
    .CLK(clknet_leaf_154_clk));
 sky130_fd_sc_hd__dfxtp_2 _42726_ (.D(_03612_),
    .Q(\cpuregs[4][12] ),
    .CLK(clknet_leaf_155_clk));
 sky130_fd_sc_hd__dfxtp_2 _42727_ (.D(_03613_),
    .Q(\cpuregs[4][13] ),
    .CLK(clknet_leaf_155_clk));
 sky130_fd_sc_hd__dfxtp_2 _42728_ (.D(_03614_),
    .Q(\cpuregs[4][14] ),
    .CLK(clknet_leaf_261_clk));
 sky130_fd_sc_hd__dfxtp_2 _42729_ (.D(_03615_),
    .Q(\cpuregs[4][15] ),
    .CLK(clknet_leaf_261_clk));
 sky130_fd_sc_hd__dfxtp_2 _42730_ (.D(_03616_),
    .Q(\cpuregs[4][16] ),
    .CLK(clknet_leaf_266_clk));
 sky130_fd_sc_hd__dfxtp_2 _42731_ (.D(_03617_),
    .Q(\cpuregs[4][17] ),
    .CLK(clknet_leaf_259_clk));
 sky130_fd_sc_hd__dfxtp_2 _42732_ (.D(_03618_),
    .Q(\cpuregs[4][18] ),
    .CLK(clknet_leaf_268_clk));
 sky130_fd_sc_hd__dfxtp_2 _42733_ (.D(_03619_),
    .Q(\cpuregs[4][19] ),
    .CLK(clknet_leaf_268_clk));
 sky130_fd_sc_hd__dfxtp_2 _42734_ (.D(_03620_),
    .Q(\cpuregs[4][20] ),
    .CLK(clknet_leaf_171_clk));
 sky130_fd_sc_hd__dfxtp_2 _42735_ (.D(_03621_),
    .Q(\cpuregs[4][21] ),
    .CLK(clknet_leaf_177_clk));
 sky130_fd_sc_hd__dfxtp_2 _42736_ (.D(_03622_),
    .Q(\cpuregs[4][22] ),
    .CLK(clknet_leaf_178_clk));
 sky130_fd_sc_hd__dfxtp_2 _42737_ (.D(_03623_),
    .Q(\cpuregs[4][23] ),
    .CLK(clknet_leaf_172_clk));
 sky130_fd_sc_hd__dfxtp_2 _42738_ (.D(_03624_),
    .Q(\cpuregs[4][24] ),
    .CLK(clknet_leaf_178_clk));
 sky130_fd_sc_hd__dfxtp_2 _42739_ (.D(_03625_),
    .Q(\cpuregs[4][25] ),
    .CLK(clknet_leaf_170_clk));
 sky130_fd_sc_hd__dfxtp_2 _42740_ (.D(_03626_),
    .Q(\cpuregs[4][26] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__dfxtp_2 _42741_ (.D(_03627_),
    .Q(\cpuregs[4][27] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__dfxtp_2 _42742_ (.D(_03628_),
    .Q(\cpuregs[4][28] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__dfxtp_2 _42743_ (.D(_03629_),
    .Q(\cpuregs[4][29] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__dfxtp_2 _42744_ (.D(_03630_),
    .Q(\cpuregs[4][30] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__dfxtp_2 _42745_ (.D(_03631_),
    .Q(\cpuregs[4][31] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__dfxtp_2 _42746_ (.D(_03632_),
    .Q(mem_la_wdata[0]),
    .CLK(clknet_leaf_203_clk));
 sky130_fd_sc_hd__dfxtp_2 _42747_ (.D(_03633_),
    .Q(mem_la_wdata[1]),
    .CLK(clknet_leaf_204_clk));
 sky130_fd_sc_hd__dfxtp_2 _42748_ (.D(_03634_),
    .Q(mem_la_wdata[2]),
    .CLK(clknet_leaf_204_clk));
 sky130_fd_sc_hd__dfxtp_2 _42749_ (.D(_03635_),
    .Q(mem_la_wdata[3]),
    .CLK(clknet_leaf_204_clk));
 sky130_fd_sc_hd__dfxtp_2 _42750_ (.D(_03636_),
    .Q(mem_la_wdata[4]),
    .CLK(clknet_leaf_204_clk));
 sky130_fd_sc_hd__dfxtp_2 _42751_ (.D(_03637_),
    .Q(mem_la_wdata[5]),
    .CLK(clknet_leaf_113_clk));
 sky130_fd_sc_hd__dfxtp_2 _42752_ (.D(_03638_),
    .Q(mem_la_wdata[6]),
    .CLK(clknet_leaf_203_clk));
 sky130_fd_sc_hd__dfxtp_2 _42753_ (.D(_03639_),
    .Q(mem_la_wdata[7]),
    .CLK(clknet_leaf_203_clk));
 sky130_fd_sc_hd__dfxtp_2 _42754_ (.D(_03640_),
    .Q(pcpi_rs2[8]),
    .CLK(clknet_leaf_197_clk));
 sky130_fd_sc_hd__dfxtp_2 _42755_ (.D(_03641_),
    .Q(pcpi_rs2[9]),
    .CLK(clknet_leaf_198_clk));
 sky130_fd_sc_hd__dfxtp_2 _42756_ (.D(_03642_),
    .Q(pcpi_rs2[10]),
    .CLK(clknet_leaf_198_clk));
 sky130_fd_sc_hd__dfxtp_2 _42757_ (.D(_03643_),
    .Q(pcpi_rs2[11]),
    .CLK(clknet_leaf_194_clk));
 sky130_fd_sc_hd__dfxtp_2 _42758_ (.D(_03644_),
    .Q(pcpi_rs2[12]),
    .CLK(clknet_leaf_188_clk));
 sky130_fd_sc_hd__dfxtp_2 _42759_ (.D(_03645_),
    .Q(pcpi_rs2[13]),
    .CLK(clknet_leaf_189_clk));
 sky130_fd_sc_hd__dfxtp_2 _42760_ (.D(_03646_),
    .Q(pcpi_rs2[14]),
    .CLK(clknet_leaf_188_clk));
 sky130_fd_sc_hd__dfxtp_2 _42761_ (.D(_03647_),
    .Q(pcpi_rs2[15]),
    .CLK(clknet_leaf_189_clk));
 sky130_fd_sc_hd__dfxtp_2 _42762_ (.D(_03648_),
    .Q(pcpi_rs2[16]),
    .CLK(clknet_leaf_185_clk));
 sky130_fd_sc_hd__dfxtp_2 _42763_ (.D(_03649_),
    .Q(pcpi_rs2[17]),
    .CLK(clknet_leaf_185_clk));
 sky130_fd_sc_hd__dfxtp_2 _42764_ (.D(_03650_),
    .Q(pcpi_rs2[18]),
    .CLK(clknet_leaf_190_clk));
 sky130_fd_sc_hd__dfxtp_2 _42765_ (.D(_03651_),
    .Q(pcpi_rs2[19]),
    .CLK(clknet_leaf_184_clk));
 sky130_fd_sc_hd__dfxtp_2 _42766_ (.D(_03652_),
    .Q(pcpi_rs2[20]),
    .CLK(clknet_leaf_190_clk));
 sky130_fd_sc_hd__dfxtp_2 _42767_ (.D(_03653_),
    .Q(pcpi_rs2[21]),
    .CLK(clknet_leaf_190_clk));
 sky130_fd_sc_hd__dfxtp_2 _42768_ (.D(_03654_),
    .Q(pcpi_rs2[22]),
    .CLK(clknet_leaf_189_clk));
 sky130_fd_sc_hd__dfxtp_2 _42769_ (.D(_03655_),
    .Q(pcpi_rs2[23]),
    .CLK(clknet_leaf_191_clk));
 sky130_fd_sc_hd__dfxtp_2 _42770_ (.D(_03656_),
    .Q(pcpi_rs2[24]),
    .CLK(clknet_leaf_189_clk));
 sky130_fd_sc_hd__dfxtp_2 _42771_ (.D(_03657_),
    .Q(pcpi_rs2[25]),
    .CLK(clknet_leaf_192_clk));
 sky130_fd_sc_hd__dfxtp_2 _42772_ (.D(_03658_),
    .Q(pcpi_rs2[26]),
    .CLK(clknet_leaf_188_clk));
 sky130_fd_sc_hd__dfxtp_2 _42773_ (.D(_03659_),
    .Q(pcpi_rs2[27]),
    .CLK(clknet_leaf_194_clk));
 sky130_fd_sc_hd__dfxtp_2 _42774_ (.D(_03660_),
    .Q(pcpi_rs2[28]),
    .CLK(clknet_leaf_199_clk));
 sky130_fd_sc_hd__dfxtp_2 _42775_ (.D(_03661_),
    .Q(pcpi_rs2[29]),
    .CLK(clknet_leaf_198_clk));
 sky130_fd_sc_hd__dfxtp_2 _42776_ (.D(_03662_),
    .Q(pcpi_rs2[30]),
    .CLK(clknet_leaf_195_clk));
 sky130_fd_sc_hd__dfxtp_2 _42777_ (.D(_03663_),
    .Q(pcpi_rs2[31]),
    .CLK(clknet_leaf_197_clk));
 sky130_fd_sc_hd__dfxtp_2 _42778_ (.D(_03664_),
    .Q(\cpuregs[9][0] ),
    .CLK(clknet_leaf_242_clk));
 sky130_fd_sc_hd__dfxtp_2 _42779_ (.D(_03665_),
    .Q(\cpuregs[9][1] ),
    .CLK(clknet_leaf_241_clk));
 sky130_fd_sc_hd__dfxtp_2 _42780_ (.D(_03666_),
    .Q(\cpuregs[9][2] ),
    .CLK(clknet_leaf_141_clk));
 sky130_fd_sc_hd__dfxtp_2 _42781_ (.D(_03667_),
    .Q(\cpuregs[9][3] ),
    .CLK(clknet_leaf_140_clk));
 sky130_fd_sc_hd__dfxtp_2 _42782_ (.D(_03668_),
    .Q(\cpuregs[9][4] ),
    .CLK(clknet_leaf_128_clk));
 sky130_fd_sc_hd__dfxtp_2 _42783_ (.D(_03669_),
    .Q(\cpuregs[9][5] ),
    .CLK(clknet_leaf_130_clk));
 sky130_fd_sc_hd__dfxtp_2 _42784_ (.D(_03670_),
    .Q(\cpuregs[9][6] ),
    .CLK(clknet_leaf_132_clk));
 sky130_fd_sc_hd__dfxtp_2 _42785_ (.D(_03671_),
    .Q(\cpuregs[9][7] ),
    .CLK(clknet_leaf_142_clk));
 sky130_fd_sc_hd__dfxtp_2 _42786_ (.D(_03672_),
    .Q(\cpuregs[9][8] ),
    .CLK(clknet_leaf_160_clk));
 sky130_fd_sc_hd__dfxtp_2 _42787_ (.D(_03673_),
    .Q(\cpuregs[9][9] ),
    .CLK(clknet_leaf_146_clk));
 sky130_fd_sc_hd__dfxtp_2 _42788_ (.D(_03674_),
    .Q(\cpuregs[9][10] ),
    .CLK(clknet_leaf_146_clk));
 sky130_fd_sc_hd__dfxtp_2 _42789_ (.D(_03675_),
    .Q(\cpuregs[9][11] ),
    .CLK(clknet_leaf_152_clk));
 sky130_fd_sc_hd__dfxtp_2 _42790_ (.D(_03676_),
    .Q(\cpuregs[9][12] ),
    .CLK(clknet_leaf_158_clk));
 sky130_fd_sc_hd__dfxtp_2 _42791_ (.D(_03677_),
    .Q(\cpuregs[9][13] ),
    .CLK(clknet_leaf_159_clk));
 sky130_fd_sc_hd__dfxtp_2 _42792_ (.D(_03678_),
    .Q(\cpuregs[9][14] ),
    .CLK(clknet_leaf_263_clk));
 sky130_fd_sc_hd__dfxtp_2 _42793_ (.D(_03679_),
    .Q(\cpuregs[9][15] ),
    .CLK(clknet_leaf_263_clk));
 sky130_fd_sc_hd__dfxtp_2 _42794_ (.D(_03680_),
    .Q(\cpuregs[9][16] ),
    .CLK(clknet_leaf_265_clk));
 sky130_fd_sc_hd__dfxtp_2 _42795_ (.D(_03681_),
    .Q(\cpuregs[9][17] ),
    .CLK(clknet_leaf_255_clk));
 sky130_fd_sc_hd__dfxtp_2 _42796_ (.D(_03682_),
    .Q(\cpuregs[9][18] ),
    .CLK(clknet_leaf_265_clk));
 sky130_fd_sc_hd__dfxtp_2 _42797_ (.D(_03683_),
    .Q(\cpuregs[9][19] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__dfxtp_2 _42798_ (.D(_03684_),
    .Q(\cpuregs[9][20] ),
    .CLK(clknet_leaf_170_clk));
 sky130_fd_sc_hd__dfxtp_2 _42799_ (.D(_03685_),
    .Q(\cpuregs[9][21] ),
    .CLK(clknet_leaf_174_clk));
 sky130_fd_sc_hd__dfxtp_2 _42800_ (.D(_03686_),
    .Q(\cpuregs[9][22] ),
    .CLK(clknet_leaf_176_clk));
 sky130_fd_sc_hd__dfxtp_2 _42801_ (.D(_03687_),
    .Q(\cpuregs[9][23] ),
    .CLK(clknet_leaf_174_clk));
 sky130_fd_sc_hd__dfxtp_2 _42802_ (.D(_03688_),
    .Q(\cpuregs[9][24] ),
    .CLK(clknet_leaf_178_clk));
 sky130_fd_sc_hd__dfxtp_2 _42803_ (.D(_03689_),
    .Q(\cpuregs[9][25] ),
    .CLK(clknet_leaf_169_clk));
 sky130_fd_sc_hd__dfxtp_2 _42804_ (.D(_03690_),
    .Q(\cpuregs[9][26] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__dfxtp_2 _42805_ (.D(_03691_),
    .Q(\cpuregs[9][27] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__dfxtp_2 _42806_ (.D(_03692_),
    .Q(\cpuregs[9][28] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__dfxtp_2 _42807_ (.D(_03693_),
    .Q(\cpuregs[9][29] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__dfxtp_2 _42808_ (.D(_03694_),
    .Q(\cpuregs[9][30] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__dfxtp_2 _42809_ (.D(_03695_),
    .Q(\cpuregs[9][31] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__dfxtp_2 _42810_ (.D(_03696_),
    .Q(\cpuregs[6][0] ),
    .CLK(clknet_leaf_242_clk));
 sky130_fd_sc_hd__dfxtp_2 _42811_ (.D(_03697_),
    .Q(\cpuregs[6][1] ),
    .CLK(clknet_leaf_240_clk));
 sky130_fd_sc_hd__dfxtp_2 _42812_ (.D(_03698_),
    .Q(\cpuregs[6][2] ),
    .CLK(clknet_leaf_140_clk));
 sky130_fd_sc_hd__dfxtp_2 _42813_ (.D(_03699_),
    .Q(\cpuregs[6][3] ),
    .CLK(clknet_leaf_144_clk));
 sky130_fd_sc_hd__dfxtp_2 _42814_ (.D(_03700_),
    .Q(\cpuregs[6][4] ),
    .CLK(clknet_leaf_127_clk));
 sky130_fd_sc_hd__dfxtp_2 _42815_ (.D(_03701_),
    .Q(\cpuregs[6][5] ),
    .CLK(clknet_leaf_129_clk));
 sky130_fd_sc_hd__dfxtp_2 _42816_ (.D(_03702_),
    .Q(\cpuregs[6][6] ),
    .CLK(clknet_leaf_133_clk));
 sky130_fd_sc_hd__dfxtp_2 _42817_ (.D(_03703_),
    .Q(\cpuregs[6][7] ),
    .CLK(clknet_leaf_142_clk));
 sky130_fd_sc_hd__dfxtp_2 _42818_ (.D(_03704_),
    .Q(\cpuregs[6][8] ),
    .CLK(clknet_leaf_154_clk));
 sky130_fd_sc_hd__dfxtp_2 _42819_ (.D(_03705_),
    .Q(\cpuregs[6][9] ),
    .CLK(clknet_leaf_149_clk));
 sky130_fd_sc_hd__dfxtp_2 _42820_ (.D(_03706_),
    .Q(\cpuregs[6][10] ),
    .CLK(clknet_leaf_149_clk));
 sky130_fd_sc_hd__dfxtp_2 _42821_ (.D(_03707_),
    .Q(\cpuregs[6][11] ),
    .CLK(clknet_leaf_154_clk));
 sky130_fd_sc_hd__dfxtp_2 _42822_ (.D(_03708_),
    .Q(\cpuregs[6][12] ),
    .CLK(clknet_leaf_155_clk));
 sky130_fd_sc_hd__dfxtp_2 _42823_ (.D(_03709_),
    .Q(\cpuregs[6][13] ),
    .CLK(clknet_leaf_155_clk));
 sky130_fd_sc_hd__dfxtp_2 _42824_ (.D(_03710_),
    .Q(\cpuregs[6][14] ),
    .CLK(clknet_leaf_261_clk));
 sky130_fd_sc_hd__dfxtp_2 _42825_ (.D(_03711_),
    .Q(\cpuregs[6][15] ),
    .CLK(clknet_leaf_260_clk));
 sky130_fd_sc_hd__dfxtp_2 _42826_ (.D(_03712_),
    .Q(\cpuregs[6][16] ),
    .CLK(clknet_leaf_266_clk));
 sky130_fd_sc_hd__dfxtp_2 _42827_ (.D(_03713_),
    .Q(\cpuregs[6][17] ),
    .CLK(clknet_leaf_259_clk));
 sky130_fd_sc_hd__dfxtp_2 _42828_ (.D(_03714_),
    .Q(\cpuregs[6][18] ),
    .CLK(clknet_leaf_267_clk));
 sky130_fd_sc_hd__dfxtp_2 _42829_ (.D(_03715_),
    .Q(\cpuregs[6][19] ),
    .CLK(clknet_leaf_266_clk));
 sky130_fd_sc_hd__dfxtp_2 _42830_ (.D(_03716_),
    .Q(\cpuregs[6][20] ),
    .CLK(clknet_leaf_170_clk));
 sky130_fd_sc_hd__dfxtp_2 _42831_ (.D(_03717_),
    .Q(\cpuregs[6][21] ),
    .CLK(clknet_leaf_173_clk));
 sky130_fd_sc_hd__dfxtp_2 _42832_ (.D(_03718_),
    .Q(\cpuregs[6][22] ),
    .CLK(clknet_leaf_178_clk));
 sky130_fd_sc_hd__dfxtp_2 _42833_ (.D(_03719_),
    .Q(\cpuregs[6][23] ),
    .CLK(clknet_leaf_171_clk));
 sky130_fd_sc_hd__dfxtp_2 _42834_ (.D(_03720_),
    .Q(\cpuregs[6][24] ),
    .CLK(clknet_leaf_178_clk));
 sky130_fd_sc_hd__dfxtp_2 _42835_ (.D(_03721_),
    .Q(\cpuregs[6][25] ),
    .CLK(clknet_leaf_170_clk));
 sky130_fd_sc_hd__dfxtp_2 _42836_ (.D(_03722_),
    .Q(\cpuregs[6][26] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__dfxtp_2 _42837_ (.D(_03723_),
    .Q(\cpuregs[6][27] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__dfxtp_2 _42838_ (.D(_03724_),
    .Q(\cpuregs[6][28] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__dfxtp_2 _42839_ (.D(_03725_),
    .Q(\cpuregs[6][29] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__dfxtp_2 _42840_ (.D(_03726_),
    .Q(\cpuregs[6][30] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__dfxtp_2 _42841_ (.D(_03727_),
    .Q(\cpuregs[6][31] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__dfxtp_2 _42842_ (.D(_03728_),
    .Q(\pcpi_mul.active[0] ),
    .CLK(clknet_5_6_0_clk));
 sky130_fd_sc_hd__dfxtp_2 _42843_ (.D(_03729_),
    .Q(\pcpi_mul.active[1] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__dfxtp_2 _42844_ (.D(_03730_),
    .Q(trap),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__dfxtp_2 _42845_ (.D(_03731_),
    .Q(\count_cycle[0] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__dfxtp_2 _42846_ (.D(_03732_),
    .Q(\count_cycle[1] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__dfxtp_2 _42847_ (.D(_03733_),
    .Q(\count_cycle[2] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfxtp_2 _42848_ (.D(_03734_),
    .Q(\count_cycle[3] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfxtp_2 _42849_ (.D(_03735_),
    .Q(\count_cycle[4] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfxtp_2 _42850_ (.D(_03736_),
    .Q(\count_cycle[5] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__dfxtp_2 _42851_ (.D(_03737_),
    .Q(\count_cycle[6] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__dfxtp_2 _42852_ (.D(_03738_),
    .Q(\count_cycle[7] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__dfxtp_2 _42853_ (.D(_03739_),
    .Q(\count_cycle[8] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__dfxtp_2 _42854_ (.D(_03740_),
    .Q(\count_cycle[9] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__dfxtp_2 _42855_ (.D(_03741_),
    .Q(\count_cycle[10] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__dfxtp_2 _42856_ (.D(_03742_),
    .Q(\count_cycle[11] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__dfxtp_2 _42857_ (.D(_03743_),
    .Q(\count_cycle[12] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__dfxtp_2 _42858_ (.D(_03744_),
    .Q(\count_cycle[13] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__dfxtp_2 _42859_ (.D(_03745_),
    .Q(\count_cycle[14] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__dfxtp_2 _42860_ (.D(_03746_),
    .Q(\count_cycle[15] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__dfxtp_2 _42861_ (.D(_03747_),
    .Q(\count_cycle[16] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__dfxtp_2 _42862_ (.D(_03748_),
    .Q(\count_cycle[17] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__dfxtp_2 _42863_ (.D(_03749_),
    .Q(\count_cycle[18] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__dfxtp_2 _42864_ (.D(_03750_),
    .Q(\count_cycle[19] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__dfxtp_2 _42865_ (.D(_03751_),
    .Q(\count_cycle[20] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfxtp_2 _42866_ (.D(_03752_),
    .Q(\count_cycle[21] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfxtp_2 _42867_ (.D(_03753_),
    .Q(\count_cycle[22] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__dfxtp_2 _42868_ (.D(_03754_),
    .Q(\count_cycle[23] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__dfxtp_2 _42869_ (.D(_03755_),
    .Q(\count_cycle[24] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__dfxtp_2 _42870_ (.D(_03756_),
    .Q(\count_cycle[25] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__dfxtp_2 _42871_ (.D(_03757_),
    .Q(\count_cycle[26] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__dfxtp_2 _42872_ (.D(_03758_),
    .Q(\count_cycle[27] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__dfxtp_2 _42873_ (.D(_03759_),
    .Q(\count_cycle[28] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__dfxtp_2 _42874_ (.D(_03760_),
    .Q(\count_cycle[29] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__dfxtp_2 _42875_ (.D(_03761_),
    .Q(\count_cycle[30] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__dfxtp_2 _42876_ (.D(_03762_),
    .Q(\count_cycle[31] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__dfxtp_2 _42877_ (.D(_03763_),
    .Q(\count_cycle[32] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__dfxtp_2 _42878_ (.D(_03764_),
    .Q(\count_cycle[33] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__dfxtp_2 _42879_ (.D(_03765_),
    .Q(\count_cycle[34] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfxtp_2 _42880_ (.D(_03766_),
    .Q(\count_cycle[35] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfxtp_2 _42881_ (.D(_03767_),
    .Q(\count_cycle[36] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__dfxtp_2 _42882_ (.D(_03768_),
    .Q(\count_cycle[37] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__dfxtp_2 _42883_ (.D(_03769_),
    .Q(\count_cycle[38] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__dfxtp_2 _42884_ (.D(_03770_),
    .Q(\count_cycle[39] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__dfxtp_2 _42885_ (.D(_03771_),
    .Q(\count_cycle[40] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__dfxtp_2 _42886_ (.D(_03772_),
    .Q(\count_cycle[41] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__dfxtp_2 _42887_ (.D(_03773_),
    .Q(\count_cycle[42] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__dfxtp_2 _42888_ (.D(_03774_),
    .Q(\count_cycle[43] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__dfxtp_2 _42889_ (.D(_03775_),
    .Q(\count_cycle[44] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__dfxtp_2 _42890_ (.D(_03776_),
    .Q(\count_cycle[45] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__dfxtp_2 _42891_ (.D(_03777_),
    .Q(\count_cycle[46] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__dfxtp_2 _42892_ (.D(_03778_),
    .Q(\count_cycle[47] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__dfxtp_2 _42893_ (.D(_03779_),
    .Q(\count_cycle[48] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__dfxtp_2 _42894_ (.D(_03780_),
    .Q(\count_cycle[49] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__dfxtp_2 _42895_ (.D(_03781_),
    .Q(\count_cycle[50] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__dfxtp_2 _42896_ (.D(_03782_),
    .Q(\count_cycle[51] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__dfxtp_2 _42897_ (.D(_03783_),
    .Q(\count_cycle[52] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__dfxtp_2 _42898_ (.D(_03784_),
    .Q(\count_cycle[53] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__dfxtp_2 _42899_ (.D(_03785_),
    .Q(\count_cycle[54] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfxtp_2 _42900_ (.D(_03786_),
    .Q(\count_cycle[55] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfxtp_2 _42901_ (.D(_03787_),
    .Q(\count_cycle[56] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfxtp_2 _42902_ (.D(_03788_),
    .Q(\count_cycle[57] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfxtp_2 _42903_ (.D(_03789_),
    .Q(\count_cycle[58] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfxtp_2 _42904_ (.D(_03790_),
    .Q(\count_cycle[59] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfxtp_2 _42905_ (.D(_03791_),
    .Q(\count_cycle[60] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__dfxtp_2 _42906_ (.D(_03792_),
    .Q(\count_cycle[61] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfxtp_2 _42907_ (.D(_03793_),
    .Q(\count_cycle[62] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__dfxtp_2 _42908_ (.D(_03794_),
    .Q(\count_cycle[63] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfxtp_2 _42909_ (.D(_03795_),
    .Q(\timer[0] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__dfxtp_2 _42910_ (.D(_03796_),
    .Q(\timer[1] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__dfxtp_2 _42911_ (.D(_03797_),
    .Q(\timer[2] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__dfxtp_2 _42912_ (.D(_03798_),
    .Q(\timer[3] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__dfxtp_2 _42913_ (.D(_03799_),
    .Q(\timer[4] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__dfxtp_2 _42914_ (.D(_03800_),
    .Q(\timer[5] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__dfxtp_2 _42915_ (.D(_03801_),
    .Q(\timer[6] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__dfxtp_2 _42916_ (.D(_03802_),
    .Q(\timer[7] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__dfxtp_2 _42917_ (.D(_03803_),
    .Q(\timer[8] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__dfxtp_2 _42918_ (.D(_03804_),
    .Q(\timer[9] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__dfxtp_2 _42919_ (.D(_03805_),
    .Q(\timer[10] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__dfxtp_2 _42920_ (.D(_03806_),
    .Q(\timer[11] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__dfxtp_2 _42921_ (.D(_03807_),
    .Q(\timer[12] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__dfxtp_2 _42922_ (.D(_03808_),
    .Q(\timer[13] ),
    .CLK(clknet_5_25_0_clk));
 sky130_fd_sc_hd__dfxtp_2 _42923_ (.D(_03809_),
    .Q(\timer[14] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__dfxtp_2 _42924_ (.D(_03810_),
    .Q(\timer[15] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__dfxtp_2 _42925_ (.D(_03811_),
    .Q(\timer[16] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__dfxtp_2 _42926_ (.D(_03812_),
    .Q(\timer[17] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__dfxtp_2 _42927_ (.D(_03813_),
    .Q(\timer[18] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__dfxtp_2 _42928_ (.D(_03814_),
    .Q(\timer[19] ),
    .CLK(clknet_leaf_253_clk));
 sky130_fd_sc_hd__dfxtp_2 _42929_ (.D(_03815_),
    .Q(\timer[20] ),
    .CLK(clknet_leaf_253_clk));
 sky130_fd_sc_hd__dfxtp_2 _42930_ (.D(_03816_),
    .Q(\timer[21] ),
    .CLK(clknet_leaf_254_clk));
 sky130_fd_sc_hd__dfxtp_2 _42931_ (.D(_03817_),
    .Q(\timer[22] ),
    .CLK(clknet_leaf_255_clk));
 sky130_fd_sc_hd__dfxtp_2 _42932_ (.D(_03818_),
    .Q(\timer[23] ),
    .CLK(clknet_leaf_253_clk));
 sky130_fd_sc_hd__dfxtp_2 _42933_ (.D(_03819_),
    .Q(\timer[24] ),
    .CLK(clknet_leaf_253_clk));
 sky130_fd_sc_hd__dfxtp_2 _42934_ (.D(_03820_),
    .Q(\timer[25] ),
    .CLK(clknet_leaf_253_clk));
 sky130_fd_sc_hd__dfxtp_2 _42935_ (.D(_03821_),
    .Q(\timer[26] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__dfxtp_2 _42936_ (.D(_03822_),
    .Q(\timer[27] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__dfxtp_2 _42937_ (.D(_03823_),
    .Q(\timer[28] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__dfxtp_2 _42938_ (.D(_03824_),
    .Q(\timer[29] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__dfxtp_2 _42939_ (.D(_03825_),
    .Q(\timer[30] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__dfxtp_2 _42940_ (.D(_03826_),
    .Q(\timer[31] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__dfxtp_2 _42941_ (.D(_03827_),
    .Q(pcpi_timeout),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__dfxtp_2 _42942_ (.D(_03828_),
    .Q(decoder_pseudo_trigger),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__dfxtp_2 _42943_ (.D(_03829_),
    .Q(is_compare),
    .CLK(clknet_5_15_0_clk));
 sky130_fd_sc_hd__dfxtp_2 _42944_ (.D(_03830_),
    .Q(do_waitirq),
    .CLK(clknet_leaf_221_clk));
 sky130_fd_sc_hd__dfxtp_2 _42945_ (.D(_03831_),
    .Q(mem_valid),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__dfxtp_2 _42946_ (.D(_03832_),
    .Q(pcpi_valid),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfxtp_2 _42947_ (.D(_03833_),
    .Q(eoi[0]),
    .CLK(clknet_leaf_223_clk));
 sky130_fd_sc_hd__dfxtp_2 _42948_ (.D(_03834_),
    .Q(eoi[1]),
    .CLK(clknet_leaf_250_clk));
 sky130_fd_sc_hd__dfxtp_2 _42949_ (.D(_03835_),
    .Q(eoi[2]),
    .CLK(clknet_leaf_225_clk));
 sky130_fd_sc_hd__dfxtp_2 _42950_ (.D(_03836_),
    .Q(eoi[3]),
    .CLK(clknet_leaf_248_clk));
 sky130_fd_sc_hd__dfxtp_2 _42951_ (.D(_03837_),
    .Q(eoi[4]),
    .CLK(clknet_leaf_250_clk));
 sky130_fd_sc_hd__dfxtp_2 _42952_ (.D(_03838_),
    .Q(eoi[5]),
    .CLK(clknet_leaf_223_clk));
 sky130_fd_sc_hd__dfxtp_2 _42953_ (.D(_03839_),
    .Q(eoi[6]),
    .CLK(clknet_leaf_223_clk));
 sky130_fd_sc_hd__dfxtp_2 _42954_ (.D(_03840_),
    .Q(eoi[7]),
    .CLK(clknet_leaf_250_clk));
 sky130_fd_sc_hd__dfxtp_2 _42955_ (.D(_03841_),
    .Q(eoi[8]),
    .CLK(clknet_leaf_250_clk));
 sky130_fd_sc_hd__dfxtp_2 _42956_ (.D(_03842_),
    .Q(eoi[9]),
    .CLK(clknet_leaf_250_clk));
 sky130_fd_sc_hd__dfxtp_2 _42957_ (.D(_03843_),
    .Q(eoi[10]),
    .CLK(clknet_leaf_248_clk));
 sky130_fd_sc_hd__dfxtp_2 _42958_ (.D(_03844_),
    .Q(eoi[11]),
    .CLK(clknet_leaf_249_clk));
 sky130_fd_sc_hd__dfxtp_2 _42959_ (.D(_03845_),
    .Q(eoi[12]),
    .CLK(clknet_leaf_248_clk));
 sky130_fd_sc_hd__dfxtp_2 _42960_ (.D(_03846_),
    .Q(eoi[13]),
    .CLK(clknet_leaf_247_clk));
 sky130_fd_sc_hd__dfxtp_2 _42961_ (.D(_03847_),
    .Q(eoi[14]),
    .CLK(clknet_leaf_249_clk));
 sky130_fd_sc_hd__dfxtp_2 _42962_ (.D(_03848_),
    .Q(eoi[15]),
    .CLK(clknet_leaf_249_clk));
 sky130_fd_sc_hd__dfxtp_2 _42963_ (.D(_03849_),
    .Q(eoi[16]),
    .CLK(clknet_leaf_247_clk));
 sky130_fd_sc_hd__dfxtp_2 _42964_ (.D(_03850_),
    .Q(eoi[17]),
    .CLK(clknet_leaf_246_clk));
 sky130_fd_sc_hd__dfxtp_2 _42965_ (.D(_03851_),
    .Q(eoi[18]),
    .CLK(clknet_leaf_247_clk));
 sky130_fd_sc_hd__dfxtp_2 _42966_ (.D(_03852_),
    .Q(eoi[19]),
    .CLK(clknet_leaf_247_clk));
 sky130_fd_sc_hd__dfxtp_2 _42967_ (.D(_03853_),
    .Q(eoi[20]),
    .CLK(clknet_leaf_246_clk));
 sky130_fd_sc_hd__dfxtp_2 _42968_ (.D(_03854_),
    .Q(eoi[21]),
    .CLK(clknet_leaf_246_clk));
 sky130_fd_sc_hd__dfxtp_2 _42969_ (.D(_03855_),
    .Q(eoi[22]),
    .CLK(clknet_leaf_245_clk));
 sky130_fd_sc_hd__dfxtp_2 _42970_ (.D(_03856_),
    .Q(eoi[23]),
    .CLK(clknet_leaf_246_clk));
 sky130_fd_sc_hd__dfxtp_2 _42971_ (.D(_03857_),
    .Q(eoi[24]),
    .CLK(clknet_leaf_249_clk));
 sky130_fd_sc_hd__dfxtp_2 _42972_ (.D(_03858_),
    .Q(eoi[25]),
    .CLK(clknet_leaf_245_clk));
 sky130_fd_sc_hd__dfxtp_2 _42973_ (.D(_03859_),
    .Q(eoi[26]),
    .CLK(clknet_leaf_250_clk));
 sky130_fd_sc_hd__dfxtp_2 _42974_ (.D(_03860_),
    .Q(eoi[27]),
    .CLK(clknet_leaf_223_clk));
 sky130_fd_sc_hd__dfxtp_2 _42975_ (.D(_03861_),
    .Q(eoi[28]),
    .CLK(clknet_leaf_251_clk));
 sky130_fd_sc_hd__dfxtp_2 _42976_ (.D(_03862_),
    .Q(eoi[29]),
    .CLK(clknet_leaf_251_clk));
 sky130_fd_sc_hd__dfxtp_2 _42977_ (.D(_03863_),
    .Q(eoi[30]),
    .CLK(clknet_leaf_251_clk));
 sky130_fd_sc_hd__dfxtp_2 _42978_ (.D(_03864_),
    .Q(eoi[31]),
    .CLK(clknet_leaf_223_clk));
 sky130_fd_sc_hd__dfxtp_2 _42979_ (.D(_03865_),
    .Q(\count_instr[0] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__dfxtp_2 _42980_ (.D(_03866_),
    .Q(\count_instr[1] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfxtp_2 _42981_ (.D(_03867_),
    .Q(\count_instr[2] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__dfxtp_2 _42982_ (.D(_03868_),
    .Q(\count_instr[3] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfxtp_2 _42983_ (.D(_03869_),
    .Q(\count_instr[4] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfxtp_2 _42984_ (.D(_03870_),
    .Q(\count_instr[5] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfxtp_2 _42985_ (.D(_03871_),
    .Q(\count_instr[6] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__dfxtp_2 _42986_ (.D(_03872_),
    .Q(\count_instr[7] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__dfxtp_2 _42987_ (.D(_03873_),
    .Q(\count_instr[8] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__dfxtp_2 _42988_ (.D(_03874_),
    .Q(\count_instr[9] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__dfxtp_2 _42989_ (.D(_03875_),
    .Q(\count_instr[10] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__dfxtp_2 _42990_ (.D(_03876_),
    .Q(\count_instr[11] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__dfxtp_2 _42991_ (.D(_03877_),
    .Q(\count_instr[12] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfxtp_2 _42992_ (.D(_03878_),
    .Q(\count_instr[13] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__dfxtp_2 _42993_ (.D(_03879_),
    .Q(\count_instr[14] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__dfxtp_2 _42994_ (.D(_03880_),
    .Q(\count_instr[15] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__dfxtp_2 _42995_ (.D(_03881_),
    .Q(\count_instr[16] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__dfxtp_2 _42996_ (.D(_03882_),
    .Q(\count_instr[17] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__dfxtp_2 _42997_ (.D(_03883_),
    .Q(\count_instr[18] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__dfxtp_2 _42998_ (.D(_03884_),
    .Q(\count_instr[19] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfxtp_2 _42999_ (.D(_03885_),
    .Q(\count_instr[20] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfxtp_2 _43000_ (.D(_03886_),
    .Q(\count_instr[21] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfxtp_2 _43001_ (.D(_03887_),
    .Q(\count_instr[22] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfxtp_2 _43002_ (.D(_03888_),
    .Q(\count_instr[23] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__dfxtp_2 _43003_ (.D(_03889_),
    .Q(\count_instr[24] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfxtp_2 _43004_ (.D(_03890_),
    .Q(\count_instr[25] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfxtp_2 _43005_ (.D(_03891_),
    .Q(\count_instr[26] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__dfxtp_2 _43006_ (.D(_03892_),
    .Q(\count_instr[27] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__dfxtp_2 _43007_ (.D(_03893_),
    .Q(\count_instr[28] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__dfxtp_2 _43008_ (.D(_03894_),
    .Q(\count_instr[29] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfxtp_2 _43009_ (.D(_03895_),
    .Q(\count_instr[30] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfxtp_2 _43010_ (.D(_03896_),
    .Q(\count_instr[31] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__dfxtp_2 _43011_ (.D(_03897_),
    .Q(\count_instr[32] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__dfxtp_2 _43012_ (.D(_03898_),
    .Q(\count_instr[33] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfxtp_2 _43013_ (.D(_03899_),
    .Q(\count_instr[34] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfxtp_2 _43014_ (.D(_03900_),
    .Q(\count_instr[35] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfxtp_2 _43015_ (.D(_03901_),
    .Q(\count_instr[36] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfxtp_2 _43016_ (.D(_03902_),
    .Q(\count_instr[37] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__dfxtp_2 _43017_ (.D(_03903_),
    .Q(\count_instr[38] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__dfxtp_2 _43018_ (.D(_03904_),
    .Q(\count_instr[39] ),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__dfxtp_2 _43019_ (.D(_03905_),
    .Q(\count_instr[40] ),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__dfxtp_2 _43020_ (.D(_03906_),
    .Q(\count_instr[41] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__dfxtp_2 _43021_ (.D(_03907_),
    .Q(\count_instr[42] ),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__dfxtp_2 _43022_ (.D(_03908_),
    .Q(\count_instr[43] ),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__dfxtp_2 _43023_ (.D(_03909_),
    .Q(\count_instr[44] ),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__dfxtp_2 _43024_ (.D(_03910_),
    .Q(\count_instr[45] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__dfxtp_2 _43025_ (.D(_03911_),
    .Q(\count_instr[46] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__dfxtp_2 _43026_ (.D(_03912_),
    .Q(\count_instr[47] ),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__dfxtp_2 _43027_ (.D(_03913_),
    .Q(\count_instr[48] ),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__dfxtp_2 _43028_ (.D(_03914_),
    .Q(\count_instr[49] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__dfxtp_2 _43029_ (.D(_03915_),
    .Q(\count_instr[50] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__dfxtp_2 _43030_ (.D(_03916_),
    .Q(\count_instr[51] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__dfxtp_2 _43031_ (.D(_03917_),
    .Q(\count_instr[52] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__dfxtp_2 _43032_ (.D(_03918_),
    .Q(\count_instr[53] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__dfxtp_2 _43033_ (.D(_03919_),
    .Q(\count_instr[54] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__dfxtp_2 _43034_ (.D(_03920_),
    .Q(\count_instr[55] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__dfxtp_2 _43035_ (.D(_03921_),
    .Q(\count_instr[56] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__dfxtp_2 _43036_ (.D(_03922_),
    .Q(\count_instr[57] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__dfxtp_2 _43037_ (.D(_03923_),
    .Q(\count_instr[58] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfxtp_2 _43038_ (.D(_03924_),
    .Q(\count_instr[59] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfxtp_2 _43039_ (.D(_03925_),
    .Q(\count_instr[60] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__dfxtp_2 _43040_ (.D(_03926_),
    .Q(\count_instr[61] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfxtp_2 _43041_ (.D(_03927_),
    .Q(\count_instr[62] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfxtp_2 _43042_ (.D(_03928_),
    .Q(\count_instr[63] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfxtp_2 _43043_ (.D(_03929_),
    .Q(\reg_pc[1] ),
    .CLK(clknet_leaf_227_clk));
 sky130_fd_sc_hd__dfxtp_2 _43044_ (.D(_03930_),
    .Q(\reg_pc[2] ),
    .CLK(clknet_leaf_227_clk));
 sky130_fd_sc_hd__dfxtp_2 _43045_ (.D(_03931_),
    .Q(\reg_pc[3] ),
    .CLK(clknet_leaf_200_clk));
 sky130_fd_sc_hd__dfxtp_2 _43046_ (.D(_03932_),
    .Q(\reg_pc[4] ),
    .CLK(clknet_leaf_200_clk));
 sky130_fd_sc_hd__dfxtp_2 _43047_ (.D(_03933_),
    .Q(\reg_pc[5] ),
    .CLK(clknet_leaf_187_clk));
 sky130_fd_sc_hd__dfxtp_2 _43048_ (.D(_03934_),
    .Q(\reg_pc[6] ),
    .CLK(clknet_leaf_187_clk));
 sky130_fd_sc_hd__dfxtp_2 _43049_ (.D(_03935_),
    .Q(\reg_pc[7] ),
    .CLK(clknet_leaf_187_clk));
 sky130_fd_sc_hd__dfxtp_2 _43050_ (.D(_03936_),
    .Q(\reg_pc[8] ),
    .CLK(clknet_leaf_186_clk));
 sky130_fd_sc_hd__dfxtp_2 _43051_ (.D(_03937_),
    .Q(\reg_pc[9] ),
    .CLK(clknet_leaf_186_clk));
 sky130_fd_sc_hd__dfxtp_2 _43052_ (.D(_03938_),
    .Q(\reg_pc[10] ),
    .CLK(clknet_leaf_186_clk));
 sky130_fd_sc_hd__dfxtp_2 _43053_ (.D(_03939_),
    .Q(\reg_pc[11] ),
    .CLK(clknet_leaf_185_clk));
 sky130_fd_sc_hd__dfxtp_2 _43054_ (.D(_03940_),
    .Q(\reg_pc[12] ),
    .CLK(clknet_leaf_182_clk));
 sky130_fd_sc_hd__dfxtp_2 _43055_ (.D(_03941_),
    .Q(\reg_pc[13] ),
    .CLK(clknet_leaf_182_clk));
 sky130_fd_sc_hd__dfxtp_2 _43056_ (.D(_03942_),
    .Q(\reg_pc[14] ),
    .CLK(clknet_leaf_181_clk));
 sky130_fd_sc_hd__dfxtp_2 _43057_ (.D(_03943_),
    .Q(\reg_pc[15] ),
    .CLK(clknet_leaf_181_clk));
 sky130_fd_sc_hd__dfxtp_2 _43058_ (.D(_03944_),
    .Q(\reg_pc[16] ),
    .CLK(clknet_leaf_181_clk));
 sky130_fd_sc_hd__dfxtp_2 _43059_ (.D(_03945_),
    .Q(\reg_pc[17] ),
    .CLK(clknet_leaf_181_clk));
 sky130_fd_sc_hd__dfxtp_2 _43060_ (.D(_03946_),
    .Q(\reg_pc[18] ),
    .CLK(clknet_leaf_181_clk));
 sky130_fd_sc_hd__dfxtp_2 _43061_ (.D(_03947_),
    .Q(\reg_pc[19] ),
    .CLK(clknet_leaf_181_clk));
 sky130_fd_sc_hd__dfxtp_2 _43062_ (.D(_03948_),
    .Q(\reg_pc[20] ),
    .CLK(clknet_leaf_179_clk));
 sky130_fd_sc_hd__dfxtp_2 _43063_ (.D(_03949_),
    .Q(\reg_pc[21] ),
    .CLK(clknet_leaf_179_clk));
 sky130_fd_sc_hd__dfxtp_2 _43064_ (.D(_03950_),
    .Q(\reg_pc[22] ),
    .CLK(clknet_leaf_179_clk));
 sky130_fd_sc_hd__dfxtp_2 _43065_ (.D(_03951_),
    .Q(\reg_pc[23] ),
    .CLK(clknet_leaf_180_clk));
 sky130_fd_sc_hd__dfxtp_2 _43066_ (.D(_03952_),
    .Q(\reg_pc[24] ),
    .CLK(clknet_leaf_181_clk));
 sky130_fd_sc_hd__dfxtp_2 _43067_ (.D(_03953_),
    .Q(\reg_pc[25] ),
    .CLK(clknet_leaf_181_clk));
 sky130_fd_sc_hd__dfxtp_2 _43068_ (.D(_03954_),
    .Q(\reg_pc[26] ),
    .CLK(clknet_leaf_237_clk));
 sky130_fd_sc_hd__dfxtp_2 _43069_ (.D(_03955_),
    .Q(\reg_pc[27] ),
    .CLK(clknet_leaf_237_clk));
 sky130_fd_sc_hd__dfxtp_2 _43070_ (.D(_03956_),
    .Q(\reg_pc[28] ),
    .CLK(clknet_leaf_238_clk));
 sky130_fd_sc_hd__dfxtp_2 _43071_ (.D(_03957_),
    .Q(\reg_pc[29] ),
    .CLK(clknet_leaf_238_clk));
 sky130_fd_sc_hd__dfxtp_2 _43072_ (.D(_03958_),
    .Q(\reg_pc[30] ),
    .CLK(clknet_leaf_227_clk));
 sky130_fd_sc_hd__dfxtp_2 _43073_ (.D(_03959_),
    .Q(\reg_pc[31] ),
    .CLK(clknet_leaf_226_clk));
 sky130_fd_sc_hd__dfxtp_2 _43074_ (.D(_03960_),
    .Q(\reg_next_pc[1] ),
    .CLK(clknet_leaf_227_clk));
 sky130_fd_sc_hd__dfxtp_2 _43075_ (.D(_03961_),
    .Q(\reg_next_pc[2] ),
    .CLK(clknet_leaf_228_clk));
 sky130_fd_sc_hd__dfxtp_2 _43076_ (.D(_03962_),
    .Q(\reg_next_pc[3] ),
    .CLK(clknet_leaf_229_clk));
 sky130_fd_sc_hd__dfxtp_2 _43077_ (.D(_03963_),
    .Q(\reg_next_pc[4] ),
    .CLK(clknet_leaf_229_clk));
 sky130_fd_sc_hd__dfxtp_2 _43078_ (.D(_03964_),
    .Q(\reg_next_pc[5] ),
    .CLK(clknet_leaf_228_clk));
 sky130_fd_sc_hd__dfxtp_2 _43079_ (.D(_03965_),
    .Q(\reg_next_pc[6] ),
    .CLK(clknet_leaf_229_clk));
 sky130_fd_sc_hd__dfxtp_2 _43080_ (.D(_03966_),
    .Q(\reg_next_pc[7] ),
    .CLK(clknet_leaf_229_clk));
 sky130_fd_sc_hd__dfxtp_2 _43081_ (.D(_03967_),
    .Q(\reg_next_pc[8] ),
    .CLK(clknet_leaf_230_clk));
 sky130_fd_sc_hd__dfxtp_2 _43082_ (.D(_03968_),
    .Q(\reg_next_pc[9] ),
    .CLK(clknet_leaf_230_clk));
 sky130_fd_sc_hd__dfxtp_2 _43083_ (.D(_03969_),
    .Q(\reg_next_pc[10] ),
    .CLK(clknet_leaf_231_clk));
 sky130_fd_sc_hd__dfxtp_2 _43084_ (.D(_03970_),
    .Q(\reg_next_pc[11] ),
    .CLK(clknet_leaf_231_clk));
 sky130_fd_sc_hd__dfxtp_2 _43085_ (.D(_03971_),
    .Q(\reg_next_pc[12] ),
    .CLK(clknet_leaf_230_clk));
 sky130_fd_sc_hd__dfxtp_2 _43086_ (.D(_03972_),
    .Q(\reg_next_pc[13] ),
    .CLK(clknet_leaf_230_clk));
 sky130_fd_sc_hd__dfxtp_2 _43087_ (.D(_03973_),
    .Q(\reg_next_pc[14] ),
    .CLK(clknet_leaf_233_clk));
 sky130_fd_sc_hd__dfxtp_2 _43088_ (.D(_03974_),
    .Q(\reg_next_pc[15] ),
    .CLK(clknet_leaf_233_clk));
 sky130_fd_sc_hd__dfxtp_2 _43089_ (.D(_03975_),
    .Q(\reg_next_pc[16] ),
    .CLK(clknet_leaf_237_clk));
 sky130_fd_sc_hd__dfxtp_2 _43090_ (.D(_03976_),
    .Q(\reg_next_pc[17] ),
    .CLK(clknet_leaf_237_clk));
 sky130_fd_sc_hd__dfxtp_2 _43091_ (.D(_03977_),
    .Q(\reg_next_pc[18] ),
    .CLK(clknet_leaf_236_clk));
 sky130_fd_sc_hd__dfxtp_2 _43092_ (.D(_03978_),
    .Q(\reg_next_pc[19] ),
    .CLK(clknet_leaf_237_clk));
 sky130_fd_sc_hd__dfxtp_2 _43093_ (.D(_03979_),
    .Q(\reg_next_pc[20] ),
    .CLK(clknet_leaf_235_clk));
 sky130_fd_sc_hd__dfxtp_2 _43094_ (.D(_03980_),
    .Q(\reg_next_pc[21] ),
    .CLK(clknet_leaf_235_clk));
 sky130_fd_sc_hd__dfxtp_2 _43095_ (.D(_03981_),
    .Q(\reg_next_pc[22] ),
    .CLK(clknet_leaf_235_clk));
 sky130_fd_sc_hd__dfxtp_2 _43096_ (.D(_03982_),
    .Q(\reg_next_pc[23] ),
    .CLK(clknet_leaf_180_clk));
 sky130_fd_sc_hd__dfxtp_2 _43097_ (.D(_03983_),
    .Q(\reg_next_pc[24] ),
    .CLK(clknet_leaf_235_clk));
 sky130_fd_sc_hd__dfxtp_2 _43098_ (.D(_03984_),
    .Q(\reg_next_pc[25] ),
    .CLK(clknet_leaf_237_clk));
 sky130_fd_sc_hd__dfxtp_2 _43099_ (.D(_03985_),
    .Q(\reg_next_pc[26] ),
    .CLK(clknet_leaf_237_clk));
 sky130_fd_sc_hd__dfxtp_2 _43100_ (.D(_03986_),
    .Q(\reg_next_pc[27] ),
    .CLK(clknet_leaf_239_clk));
 sky130_fd_sc_hd__dfxtp_2 _43101_ (.D(_03987_),
    .Q(\reg_next_pc[28] ),
    .CLK(clknet_leaf_238_clk));
 sky130_fd_sc_hd__dfxtp_2 _43102_ (.D(_03988_),
    .Q(\reg_next_pc[29] ),
    .CLK(clknet_leaf_238_clk));
 sky130_fd_sc_hd__dfxtp_2 _43103_ (.D(_03989_),
    .Q(\reg_next_pc[30] ),
    .CLK(clknet_leaf_238_clk));
 sky130_fd_sc_hd__dfxtp_2 _43104_ (.D(_03990_),
    .Q(\reg_next_pc[31] ),
    .CLK(clknet_leaf_247_clk));
 sky130_fd_sc_hd__dfxtp_2 _43105_ (.D(_03991_),
    .Q(mem_do_rdata),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__dfxtp_2 _43106_ (.D(_03992_),
    .Q(mem_do_wdata),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfxtp_2 _43107_ (.D(_03993_),
    .Q(\pcpi_timeout_counter[0] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__dfxtp_2 _43108_ (.D(_03994_),
    .Q(\pcpi_timeout_counter[1] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__dfxtp_2 _43109_ (.D(_03995_),
    .Q(\pcpi_timeout_counter[2] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__dfxtp_2 _43110_ (.D(_03996_),
    .Q(\pcpi_timeout_counter[3] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__dfxtp_2 _43111_ (.D(_03997_),
    .Q(instr_beq),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__dfxtp_2 _43112_ (.D(_03998_),
    .Q(instr_bne),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__dfxtp_2 _43113_ (.D(_03999_),
    .Q(instr_blt),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__dfxtp_2 _43114_ (.D(_04000_),
    .Q(instr_bge),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__dfxtp_2 _43115_ (.D(_04001_),
    .Q(instr_bltu),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__dfxtp_2 _43116_ (.D(_04002_),
    .Q(instr_bgeu),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__dfxtp_2 _43117_ (.D(_04003_),
    .Q(instr_addi),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__dfxtp_2 _43118_ (.D(_04004_),
    .Q(instr_slti),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__dfxtp_2 _43119_ (.D(_04005_),
    .Q(instr_sltiu),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__dfxtp_2 _43120_ (.D(_04006_),
    .Q(instr_xori),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__dfxtp_2 _43121_ (.D(_04007_),
    .Q(instr_ori),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__dfxtp_2 _43122_ (.D(_04008_),
    .Q(instr_andi),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__dfxtp_2 _43123_ (.D(_04009_),
    .Q(instr_add),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__dfxtp_2 _43124_ (.D(_04010_),
    .Q(instr_sub),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__dfxtp_2 _43125_ (.D(_04011_),
    .Q(instr_sll),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__dfxtp_2 _43126_ (.D(_04012_),
    .Q(instr_slt),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__dfxtp_2 _43127_ (.D(_04013_),
    .Q(instr_sltu),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__dfxtp_2 _43128_ (.D(_04014_),
    .Q(instr_xor),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__dfxtp_2 _43129_ (.D(_04015_),
    .Q(instr_srl),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__dfxtp_2 _43130_ (.D(_04016_),
    .Q(instr_sra),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__dfxtp_2 _43131_ (.D(_04017_),
    .Q(instr_or),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__dfxtp_2 _43132_ (.D(_04018_),
    .Q(instr_and),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__dfxtp_2 _43133_ (.D(_04019_),
    .Q(\decoded_rs1[0] ),
    .CLK(clknet_leaf_215_clk));
 sky130_fd_sc_hd__dfxtp_2 _43134_ (.D(_04020_),
    .Q(\decoded_rs1[1] ),
    .CLK(clknet_leaf_216_clk));
 sky130_fd_sc_hd__dfxtp_2 _43135_ (.D(_04021_),
    .Q(\decoded_rs1[2] ),
    .CLK(clknet_leaf_216_clk));
 sky130_fd_sc_hd__dfxtp_2 _43136_ (.D(_04022_),
    .Q(\decoded_rs1[3] ),
    .CLK(clknet_leaf_217_clk));
 sky130_fd_sc_hd__dfxtp_2 _43137_ (.D(_04023_),
    .Q(is_beq_bne_blt_bge_bltu_bgeu),
    .CLK(clknet_leaf_220_clk));
 sky130_fd_sc_hd__dfxtp_2 _43138_ (.D(_04024_),
    .Q(mem_instr),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__dfxtp_2 _43139_ (.D(_04025_),
    .Q(\irq_mask[0] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__dfxtp_2 _43140_ (.D(_04026_),
    .Q(\irq_mask[1] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__dfxtp_2 _43141_ (.D(_04027_),
    .Q(\irq_mask[2] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__dfxtp_2 _43142_ (.D(_04028_),
    .Q(\irq_mask[3] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__dfxtp_2 _43143_ (.D(_04029_),
    .Q(\irq_mask[4] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__dfxtp_2 _43144_ (.D(_04030_),
    .Q(\irq_mask[5] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__dfxtp_2 _43145_ (.D(_04031_),
    .Q(\irq_mask[6] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__dfxtp_2 _43146_ (.D(_04032_),
    .Q(\irq_mask[7] ),
    .CLK(clknet_leaf_251_clk));
 sky130_fd_sc_hd__dfxtp_2 _43147_ (.D(_04033_),
    .Q(\irq_mask[8] ),
    .CLK(clknet_leaf_252_clk));
 sky130_fd_sc_hd__dfxtp_2 _43148_ (.D(_04034_),
    .Q(\irq_mask[9] ),
    .CLK(clknet_leaf_252_clk));
 sky130_fd_sc_hd__dfxtp_2 _43149_ (.D(_04035_),
    .Q(\irq_mask[10] ),
    .CLK(clknet_leaf_252_clk));
 sky130_fd_sc_hd__dfxtp_2 _43150_ (.D(_04036_),
    .Q(\irq_mask[11] ),
    .CLK(clknet_leaf_252_clk));
 sky130_fd_sc_hd__dfxtp_2 _43151_ (.D(_04037_),
    .Q(\irq_mask[12] ),
    .CLK(clknet_leaf_252_clk));
 sky130_fd_sc_hd__dfxtp_2 _43152_ (.D(_04038_),
    .Q(\irq_mask[13] ),
    .CLK(clknet_leaf_252_clk));
 sky130_fd_sc_hd__dfxtp_2 _43153_ (.D(_04039_),
    .Q(\irq_mask[14] ),
    .CLK(clknet_leaf_252_clk));
 sky130_fd_sc_hd__dfxtp_2 _43154_ (.D(_04040_),
    .Q(\irq_mask[15] ),
    .CLK(clknet_leaf_249_clk));
 sky130_fd_sc_hd__dfxtp_2 _43155_ (.D(_04041_),
    .Q(\irq_mask[16] ),
    .CLK(clknet_leaf_256_clk));
 sky130_fd_sc_hd__dfxtp_2 _43156_ (.D(_04042_),
    .Q(\irq_mask[17] ),
    .CLK(clknet_leaf_245_clk));
 sky130_fd_sc_hd__dfxtp_2 _43157_ (.D(_04043_),
    .Q(\irq_mask[18] ),
    .CLK(clknet_leaf_252_clk));
 sky130_fd_sc_hd__dfxtp_2 _43158_ (.D(_04044_),
    .Q(\irq_mask[19] ),
    .CLK(clknet_leaf_256_clk));
 sky130_fd_sc_hd__dfxtp_2 _43159_ (.D(_04045_),
    .Q(\irq_mask[20] ),
    .CLK(clknet_leaf_244_clk));
 sky130_fd_sc_hd__dfxtp_2 _43160_ (.D(_04046_),
    .Q(\irq_mask[21] ),
    .CLK(clknet_leaf_245_clk));
 sky130_fd_sc_hd__dfxtp_2 _43161_ (.D(_04047_),
    .Q(\irq_mask[22] ),
    .CLK(clknet_leaf_244_clk));
 sky130_fd_sc_hd__dfxtp_2 _43162_ (.D(_04048_),
    .Q(\irq_mask[23] ),
    .CLK(clknet_leaf_244_clk));
 sky130_fd_sc_hd__dfxtp_2 _43163_ (.D(_04049_),
    .Q(\irq_mask[24] ),
    .CLK(clknet_leaf_256_clk));
 sky130_fd_sc_hd__dfxtp_2 _43164_ (.D(_04050_),
    .Q(\irq_mask[25] ),
    .CLK(clknet_leaf_256_clk));
 sky130_fd_sc_hd__dfxtp_2 _43165_ (.D(_04051_),
    .Q(\irq_mask[26] ),
    .CLK(clknet_leaf_251_clk));
 sky130_fd_sc_hd__dfxtp_2 _43166_ (.D(_04052_),
    .Q(\irq_mask[27] ),
    .CLK(clknet_leaf_251_clk));
 sky130_fd_sc_hd__dfxtp_2 _43167_ (.D(_04053_),
    .Q(\irq_mask[28] ),
    .CLK(clknet_leaf_251_clk));
 sky130_fd_sc_hd__dfxtp_2 _43168_ (.D(_04054_),
    .Q(\irq_mask[29] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__dfxtp_2 _43169_ (.D(_04055_),
    .Q(\irq_mask[30] ),
    .CLK(clknet_leaf_251_clk));
 sky130_fd_sc_hd__dfxtp_2 _43170_ (.D(_04056_),
    .Q(\irq_mask[31] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__dfxtp_2 _43171_ (.D(_04057_),
    .Q(mem_do_prefetch),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfxtp_2 _43172_ (.D(_04058_),
    .Q(mem_do_rinst),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__dfxtp_2 _43173_ (.D(_04059_),
    .Q(\irq_state[0] ),
    .CLK(clknet_leaf_221_clk));
 sky130_fd_sc_hd__dfxtp_2 _43174_ (.D(_04060_),
    .Q(\irq_state[1] ),
    .CLK(clknet_leaf_222_clk));
 sky130_fd_sc_hd__dfxtp_2 _43175_ (.D(_04061_),
    .Q(latched_store),
    .CLK(clknet_leaf_221_clk));
 sky130_fd_sc_hd__dfxtp_2 _43176_ (.D(_04062_),
    .Q(latched_stalu),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__dfxtp_2 _43177_ (.D(_04063_),
    .Q(\pcpi_mul.rs2[32] ),
    .CLK(clknet_leaf_107_clk));
 sky130_fd_sc_hd__dfxtp_2 _43178_ (.D(_04064_),
    .Q(\pcpi_mul.rs1[32] ),
    .CLK(clknet_5_7_0_clk));
 sky130_fd_sc_hd__dfxtp_2 _43179_ (.D(_04065_),
    .Q(irq_delay),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__dfxtp_2 _43180_ (.D(_04066_),
    .Q(\decoded_rs1[4] ),
    .CLK(clknet_leaf_217_clk));
 sky130_fd_sc_hd__dfxtp_2 _43181_ (.D(_04067_),
    .Q(\mem_state[0] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__dfxtp_2 _43182_ (.D(_04068_),
    .Q(\mem_state[1] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__dfxtp_2 _43183_ (.D(_04069_),
    .Q(latched_branch),
    .CLK(clknet_leaf_222_clk));
 sky130_fd_sc_hd__dfxtp_2 _43184_ (.D(_04070_),
    .Q(latched_is_lh),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__dfxtp_2 _43185_ (.D(_04071_),
    .Q(latched_is_lb),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__dfxtp_2 _43186_ (.D(_04072_),
    .Q(irq_active),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_262 ();
 sky130_fd_sc_hd__decap_3 PHY_263 ();
 sky130_fd_sc_hd__decap_3 PHY_264 ();
 sky130_fd_sc_hd__decap_3 PHY_265 ();
 sky130_fd_sc_hd__decap_3 PHY_266 ();
 sky130_fd_sc_hd__decap_3 PHY_267 ();
 sky130_fd_sc_hd__decap_3 PHY_268 ();
 sky130_fd_sc_hd__decap_3 PHY_269 ();
 sky130_fd_sc_hd__decap_3 PHY_270 ();
 sky130_fd_sc_hd__decap_3 PHY_271 ();
 sky130_fd_sc_hd__decap_3 PHY_272 ();
 sky130_fd_sc_hd__decap_3 PHY_273 ();
 sky130_fd_sc_hd__decap_3 PHY_274 ();
 sky130_fd_sc_hd__decap_3 PHY_275 ();
 sky130_fd_sc_hd__decap_3 PHY_276 ();
 sky130_fd_sc_hd__decap_3 PHY_277 ();
 sky130_fd_sc_hd__decap_3 PHY_278 ();
 sky130_fd_sc_hd__decap_3 PHY_279 ();
 sky130_fd_sc_hd__decap_3 PHY_280 ();
 sky130_fd_sc_hd__decap_3 PHY_281 ();
 sky130_fd_sc_hd__decap_3 PHY_282 ();
 sky130_fd_sc_hd__decap_3 PHY_283 ();
 sky130_fd_sc_hd__decap_3 PHY_284 ();
 sky130_fd_sc_hd__decap_3 PHY_285 ();
 sky130_fd_sc_hd__decap_3 PHY_286 ();
 sky130_fd_sc_hd__decap_3 PHY_287 ();
 sky130_fd_sc_hd__decap_3 PHY_288 ();
 sky130_fd_sc_hd__decap_3 PHY_289 ();
 sky130_fd_sc_hd__decap_3 PHY_290 ();
 sky130_fd_sc_hd__decap_3 PHY_291 ();
 sky130_fd_sc_hd__decap_3 PHY_292 ();
 sky130_fd_sc_hd__decap_3 PHY_293 ();
 sky130_fd_sc_hd__decap_3 PHY_294 ();
 sky130_fd_sc_hd__decap_3 PHY_295 ();
 sky130_fd_sc_hd__decap_3 PHY_296 ();
 sky130_fd_sc_hd__decap_3 PHY_297 ();
 sky130_fd_sc_hd__decap_3 PHY_298 ();
 sky130_fd_sc_hd__decap_3 PHY_299 ();
 sky130_fd_sc_hd__decap_3 PHY_300 ();
 sky130_fd_sc_hd__decap_3 PHY_301 ();
 sky130_fd_sc_hd__decap_3 PHY_302 ();
 sky130_fd_sc_hd__decap_3 PHY_303 ();
 sky130_fd_sc_hd__decap_3 PHY_304 ();
 sky130_fd_sc_hd__decap_3 PHY_305 ();
 sky130_fd_sc_hd__decap_3 PHY_306 ();
 sky130_fd_sc_hd__decap_3 PHY_307 ();
 sky130_fd_sc_hd__decap_3 PHY_308 ();
 sky130_fd_sc_hd__decap_3 PHY_309 ();
 sky130_fd_sc_hd__decap_3 PHY_310 ();
 sky130_fd_sc_hd__decap_3 PHY_311 ();
 sky130_fd_sc_hd__decap_3 PHY_312 ();
 sky130_fd_sc_hd__decap_3 PHY_313 ();
 sky130_fd_sc_hd__decap_3 PHY_314 ();
 sky130_fd_sc_hd__decap_3 PHY_315 ();
 sky130_fd_sc_hd__decap_3 PHY_316 ();
 sky130_fd_sc_hd__decap_3 PHY_317 ();
 sky130_fd_sc_hd__decap_3 PHY_318 ();
 sky130_fd_sc_hd__decap_3 PHY_319 ();
 sky130_fd_sc_hd__decap_3 PHY_320 ();
 sky130_fd_sc_hd__decap_3 PHY_321 ();
 sky130_fd_sc_hd__decap_3 PHY_322 ();
 sky130_fd_sc_hd__decap_3 PHY_323 ();
 sky130_fd_sc_hd__decap_3 PHY_324 ();
 sky130_fd_sc_hd__decap_3 PHY_325 ();
 sky130_fd_sc_hd__decap_3 PHY_326 ();
 sky130_fd_sc_hd__decap_3 PHY_327 ();
 sky130_fd_sc_hd__decap_3 PHY_328 ();
 sky130_fd_sc_hd__decap_3 PHY_329 ();
 sky130_fd_sc_hd__decap_3 PHY_330 ();
 sky130_fd_sc_hd__decap_3 PHY_331 ();
 sky130_fd_sc_hd__decap_3 PHY_332 ();
 sky130_fd_sc_hd__decap_3 PHY_333 ();
 sky130_fd_sc_hd__decap_3 PHY_334 ();
 sky130_fd_sc_hd__decap_3 PHY_335 ();
 sky130_fd_sc_hd__decap_3 PHY_336 ();
 sky130_fd_sc_hd__decap_3 PHY_337 ();
 sky130_fd_sc_hd__decap_3 PHY_338 ();
 sky130_fd_sc_hd__decap_3 PHY_339 ();
 sky130_fd_sc_hd__decap_3 PHY_340 ();
 sky130_fd_sc_hd__decap_3 PHY_341 ();
 sky130_fd_sc_hd__decap_3 PHY_342 ();
 sky130_fd_sc_hd__decap_3 PHY_343 ();
 sky130_fd_sc_hd__decap_3 PHY_344 ();
 sky130_fd_sc_hd__decap_3 PHY_345 ();
 sky130_fd_sc_hd__decap_3 PHY_346 ();
 sky130_fd_sc_hd__decap_3 PHY_347 ();
 sky130_fd_sc_hd__decap_3 PHY_348 ();
 sky130_fd_sc_hd__decap_3 PHY_349 ();
 sky130_fd_sc_hd__decap_3 PHY_350 ();
 sky130_fd_sc_hd__decap_3 PHY_351 ();
 sky130_fd_sc_hd__decap_3 PHY_352 ();
 sky130_fd_sc_hd__decap_3 PHY_353 ();
 sky130_fd_sc_hd__decap_3 PHY_354 ();
 sky130_fd_sc_hd__decap_3 PHY_355 ();
 sky130_fd_sc_hd__decap_3 PHY_356 ();
 sky130_fd_sc_hd__decap_3 PHY_357 ();
 sky130_fd_sc_hd__decap_3 PHY_358 ();
 sky130_fd_sc_hd__decap_3 PHY_359 ();
 sky130_fd_sc_hd__decap_3 PHY_360 ();
 sky130_fd_sc_hd__decap_3 PHY_361 ();
 sky130_fd_sc_hd__decap_3 PHY_362 ();
 sky130_fd_sc_hd__decap_3 PHY_363 ();
 sky130_fd_sc_hd__decap_3 PHY_364 ();
 sky130_fd_sc_hd__decap_3 PHY_365 ();
 sky130_fd_sc_hd__decap_3 PHY_366 ();
 sky130_fd_sc_hd__decap_3 PHY_367 ();
 sky130_fd_sc_hd__decap_3 PHY_368 ();
 sky130_fd_sc_hd__decap_3 PHY_369 ();
 sky130_fd_sc_hd__decap_3 PHY_370 ();
 sky130_fd_sc_hd__decap_3 PHY_371 ();
 sky130_fd_sc_hd__decap_3 PHY_372 ();
 sky130_fd_sc_hd__decap_3 PHY_373 ();
 sky130_fd_sc_hd__decap_3 PHY_374 ();
 sky130_fd_sc_hd__decap_3 PHY_375 ();
 sky130_fd_sc_hd__decap_3 PHY_376 ();
 sky130_fd_sc_hd__decap_3 PHY_377 ();
 sky130_fd_sc_hd__decap_3 PHY_378 ();
 sky130_fd_sc_hd__decap_3 PHY_379 ();
 sky130_fd_sc_hd__decap_3 PHY_380 ();
 sky130_fd_sc_hd__decap_3 PHY_381 ();
 sky130_fd_sc_hd__decap_3 PHY_382 ();
 sky130_fd_sc_hd__decap_3 PHY_383 ();
 sky130_fd_sc_hd__decap_3 PHY_384 ();
 sky130_fd_sc_hd__decap_3 PHY_385 ();
 sky130_fd_sc_hd__decap_3 PHY_386 ();
 sky130_fd_sc_hd__decap_3 PHY_387 ();
 sky130_fd_sc_hd__decap_3 PHY_388 ();
 sky130_fd_sc_hd__decap_3 PHY_389 ();
 sky130_fd_sc_hd__decap_3 PHY_390 ();
 sky130_fd_sc_hd__decap_3 PHY_391 ();
 sky130_fd_sc_hd__decap_3 PHY_392 ();
 sky130_fd_sc_hd__decap_3 PHY_393 ();
 sky130_fd_sc_hd__decap_3 PHY_394 ();
 sky130_fd_sc_hd__decap_3 PHY_395 ();
 sky130_fd_sc_hd__decap_3 PHY_396 ();
 sky130_fd_sc_hd__decap_3 PHY_397 ();
 sky130_fd_sc_hd__decap_3 PHY_398 ();
 sky130_fd_sc_hd__decap_3 PHY_399 ();
 sky130_fd_sc_hd__decap_3 PHY_400 ();
 sky130_fd_sc_hd__decap_3 PHY_401 ();
 sky130_fd_sc_hd__decap_3 PHY_402 ();
 sky130_fd_sc_hd__decap_3 PHY_403 ();
 sky130_fd_sc_hd__decap_3 PHY_404 ();
 sky130_fd_sc_hd__decap_3 PHY_405 ();
 sky130_fd_sc_hd__decap_3 PHY_406 ();
 sky130_fd_sc_hd__decap_3 PHY_407 ();
 sky130_fd_sc_hd__decap_3 PHY_408 ();
 sky130_fd_sc_hd__decap_3 PHY_409 ();
 sky130_fd_sc_hd__decap_3 PHY_410 ();
 sky130_fd_sc_hd__decap_3 PHY_411 ();
 sky130_fd_sc_hd__decap_3 PHY_412 ();
 sky130_fd_sc_hd__decap_3 PHY_413 ();
 sky130_fd_sc_hd__decap_3 PHY_414 ();
 sky130_fd_sc_hd__decap_3 PHY_415 ();
 sky130_fd_sc_hd__decap_3 PHY_416 ();
 sky130_fd_sc_hd__decap_3 PHY_417 ();
 sky130_fd_sc_hd__decap_3 PHY_418 ();
 sky130_fd_sc_hd__decap_3 PHY_419 ();
 sky130_fd_sc_hd__decap_3 PHY_420 ();
 sky130_fd_sc_hd__decap_3 PHY_421 ();
 sky130_fd_sc_hd__decap_3 PHY_422 ();
 sky130_fd_sc_hd__decap_3 PHY_423 ();
 sky130_fd_sc_hd__decap_3 PHY_424 ();
 sky130_fd_sc_hd__decap_3 PHY_425 ();
 sky130_fd_sc_hd__decap_3 PHY_426 ();
 sky130_fd_sc_hd__decap_3 PHY_427 ();
 sky130_fd_sc_hd__decap_3 PHY_428 ();
 sky130_fd_sc_hd__decap_3 PHY_429 ();
 sky130_fd_sc_hd__decap_3 PHY_430 ();
 sky130_fd_sc_hd__decap_3 PHY_431 ();
 sky130_fd_sc_hd__decap_3 PHY_432 ();
 sky130_fd_sc_hd__decap_3 PHY_433 ();
 sky130_fd_sc_hd__decap_3 PHY_434 ();
 sky130_fd_sc_hd__decap_3 PHY_435 ();
 sky130_fd_sc_hd__decap_3 PHY_436 ();
 sky130_fd_sc_hd__decap_3 PHY_437 ();
 sky130_fd_sc_hd__decap_3 PHY_438 ();
 sky130_fd_sc_hd__decap_3 PHY_439 ();
 sky130_fd_sc_hd__decap_3 PHY_440 ();
 sky130_fd_sc_hd__decap_3 PHY_441 ();
 sky130_fd_sc_hd__decap_3 PHY_442 ();
 sky130_fd_sc_hd__decap_3 PHY_443 ();
 sky130_fd_sc_hd__decap_3 PHY_444 ();
 sky130_fd_sc_hd__decap_3 PHY_445 ();
 sky130_fd_sc_hd__decap_3 PHY_446 ();
 sky130_fd_sc_hd__decap_3 PHY_447 ();
 sky130_fd_sc_hd__decap_3 PHY_448 ();
 sky130_fd_sc_hd__decap_3 PHY_449 ();
 sky130_fd_sc_hd__decap_3 PHY_450 ();
 sky130_fd_sc_hd__decap_3 PHY_451 ();
 sky130_fd_sc_hd__decap_3 PHY_452 ();
 sky130_fd_sc_hd__decap_3 PHY_453 ();
 sky130_fd_sc_hd__decap_3 PHY_454 ();
 sky130_fd_sc_hd__decap_3 PHY_455 ();
 sky130_fd_sc_hd__decap_3 PHY_456 ();
 sky130_fd_sc_hd__decap_3 PHY_457 ();
 sky130_fd_sc_hd__decap_3 PHY_458 ();
 sky130_fd_sc_hd__decap_3 PHY_459 ();
 sky130_fd_sc_hd__decap_3 PHY_460 ();
 sky130_fd_sc_hd__decap_3 PHY_461 ();
 sky130_fd_sc_hd__decap_3 PHY_462 ();
 sky130_fd_sc_hd__decap_3 PHY_463 ();
 sky130_fd_sc_hd__decap_3 PHY_464 ();
 sky130_fd_sc_hd__decap_3 PHY_465 ();
 sky130_fd_sc_hd__decap_3 PHY_466 ();
 sky130_fd_sc_hd__decap_3 PHY_467 ();
 sky130_fd_sc_hd__decap_3 PHY_468 ();
 sky130_fd_sc_hd__decap_3 PHY_469 ();
 sky130_fd_sc_hd__decap_3 PHY_470 ();
 sky130_fd_sc_hd__decap_3 PHY_471 ();
 sky130_fd_sc_hd__decap_3 PHY_472 ();
 sky130_fd_sc_hd__decap_3 PHY_473 ();
 sky130_fd_sc_hd__decap_3 PHY_474 ();
 sky130_fd_sc_hd__decap_3 PHY_475 ();
 sky130_fd_sc_hd__decap_3 PHY_476 ();
 sky130_fd_sc_hd__decap_3 PHY_477 ();
 sky130_fd_sc_hd__decap_3 PHY_478 ();
 sky130_fd_sc_hd__decap_3 PHY_479 ();
 sky130_fd_sc_hd__decap_3 PHY_480 ();
 sky130_fd_sc_hd__decap_3 PHY_481 ();
 sky130_fd_sc_hd__decap_3 PHY_482 ();
 sky130_fd_sc_hd__decap_3 PHY_483 ();
 sky130_fd_sc_hd__decap_3 PHY_484 ();
 sky130_fd_sc_hd__decap_3 PHY_485 ();
 sky130_fd_sc_hd__decap_3 PHY_486 ();
 sky130_fd_sc_hd__decap_3 PHY_487 ();
 sky130_fd_sc_hd__decap_3 PHY_488 ();
 sky130_fd_sc_hd__decap_3 PHY_489 ();
 sky130_fd_sc_hd__decap_3 PHY_490 ();
 sky130_fd_sc_hd__decap_3 PHY_491 ();
 sky130_fd_sc_hd__decap_3 PHY_492 ();
 sky130_fd_sc_hd__decap_3 PHY_493 ();
 sky130_fd_sc_hd__decap_3 PHY_494 ();
 sky130_fd_sc_hd__decap_3 PHY_495 ();
 sky130_fd_sc_hd__decap_3 PHY_496 ();
 sky130_fd_sc_hd__decap_3 PHY_497 ();
 sky130_fd_sc_hd__decap_3 PHY_498 ();
 sky130_fd_sc_hd__decap_3 PHY_499 ();
 sky130_fd_sc_hd__decap_3 PHY_500 ();
 sky130_fd_sc_hd__decap_3 PHY_501 ();
 sky130_fd_sc_hd__decap_3 PHY_502 ();
 sky130_fd_sc_hd__decap_3 PHY_503 ();
 sky130_fd_sc_hd__decap_3 PHY_504 ();
 sky130_fd_sc_hd__decap_3 PHY_505 ();
 sky130_fd_sc_hd__decap_3 PHY_506 ();
 sky130_fd_sc_hd__decap_3 PHY_507 ();
 sky130_fd_sc_hd__decap_3 PHY_508 ();
 sky130_fd_sc_hd__decap_3 PHY_509 ();
 sky130_fd_sc_hd__decap_3 PHY_510 ();
 sky130_fd_sc_hd__decap_3 PHY_511 ();
 sky130_fd_sc_hd__decap_3 PHY_512 ();
 sky130_fd_sc_hd__decap_3 PHY_513 ();
 sky130_fd_sc_hd__decap_3 PHY_514 ();
 sky130_fd_sc_hd__decap_3 PHY_515 ();
 sky130_fd_sc_hd__decap_3 PHY_516 ();
 sky130_fd_sc_hd__decap_3 PHY_517 ();
 sky130_fd_sc_hd__decap_3 PHY_518 ();
 sky130_fd_sc_hd__decap_3 PHY_519 ();
 sky130_fd_sc_hd__decap_3 PHY_520 ();
 sky130_fd_sc_hd__decap_3 PHY_521 ();
 sky130_fd_sc_hd__decap_3 PHY_522 ();
 sky130_fd_sc_hd__decap_3 PHY_523 ();
 sky130_fd_sc_hd__decap_3 PHY_524 ();
 sky130_fd_sc_hd__decap_3 PHY_525 ();
 sky130_fd_sc_hd__decap_3 PHY_526 ();
 sky130_fd_sc_hd__decap_3 PHY_527 ();
 sky130_fd_sc_hd__decap_3 PHY_528 ();
 sky130_fd_sc_hd__decap_3 PHY_529 ();
 sky130_fd_sc_hd__decap_3 PHY_530 ();
 sky130_fd_sc_hd__decap_3 PHY_531 ();
 sky130_fd_sc_hd__decap_3 PHY_532 ();
 sky130_fd_sc_hd__decap_3 PHY_533 ();
 sky130_fd_sc_hd__decap_3 PHY_534 ();
 sky130_fd_sc_hd__decap_3 PHY_535 ();
 sky130_fd_sc_hd__decap_3 PHY_536 ();
 sky130_fd_sc_hd__decap_3 PHY_537 ();
 sky130_fd_sc_hd__decap_3 PHY_538 ();
 sky130_fd_sc_hd__decap_3 PHY_539 ();
 sky130_fd_sc_hd__decap_3 PHY_540 ();
 sky130_fd_sc_hd__decap_3 PHY_541 ();
 sky130_fd_sc_hd__decap_3 PHY_542 ();
 sky130_fd_sc_hd__decap_3 PHY_543 ();
 sky130_fd_sc_hd__decap_3 PHY_544 ();
 sky130_fd_sc_hd__decap_3 PHY_545 ();
 sky130_fd_sc_hd__decap_3 PHY_546 ();
 sky130_fd_sc_hd__decap_3 PHY_547 ();
 sky130_fd_sc_hd__decap_3 PHY_548 ();
 sky130_fd_sc_hd__decap_3 PHY_549 ();
 sky130_fd_sc_hd__decap_3 PHY_550 ();
 sky130_fd_sc_hd__decap_3 PHY_551 ();
 sky130_fd_sc_hd__decap_3 PHY_552 ();
 sky130_fd_sc_hd__decap_3 PHY_553 ();
 sky130_fd_sc_hd__decap_3 PHY_554 ();
 sky130_fd_sc_hd__decap_3 PHY_555 ();
 sky130_fd_sc_hd__decap_3 PHY_556 ();
 sky130_fd_sc_hd__decap_3 PHY_557 ();
 sky130_fd_sc_hd__decap_3 PHY_558 ();
 sky130_fd_sc_hd__decap_3 PHY_559 ();
 sky130_fd_sc_hd__decap_3 PHY_560 ();
 sky130_fd_sc_hd__decap_3 PHY_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8766 ();
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_clk (.A(clknet_5_24_0_clk),
    .X(clknet_leaf_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_clk (.A(clknet_5_24_0_clk),
    .X(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_clk (.A(clknet_5_24_0_clk),
    .X(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_clk (.A(clknet_5_25_0_clk),
    .X(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_clk (.A(clknet_5_25_0_clk),
    .X(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_clk (.A(clknet_5_25_0_clk),
    .X(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_clk (.A(clknet_5_25_0_clk),
    .X(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_clk (.A(clknet_5_16_0_clk),
    .X(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_clk (.A(clknet_5_25_0_clk),
    .X(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_clk (.A(clknet_5_25_0_clk),
    .X(clknet_leaf_9_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_clk (.A(clknet_5_25_0_clk),
    .X(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_clk (.A(clknet_5_25_0_clk),
    .X(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_clk (.A(clknet_5_25_0_clk),
    .X(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_clk (.A(clknet_5_25_0_clk),
    .X(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_clk (.A(clknet_5_29_0_clk),
    .X(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_clk (.A(clknet_opt_31_clk),
    .X(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_clk (.A(clknet_5_16_0_clk),
    .X(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_clk (.A(clknet_5_16_0_clk),
    .X(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_clk (.A(clknet_5_16_0_clk),
    .X(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_clk (.A(clknet_5_16_0_clk),
    .X(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_clk (.A(clknet_5_16_0_clk),
    .X(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_clk (.A(clknet_5_16_0_clk),
    .X(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_clk (.A(clknet_5_16_0_clk),
    .X(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_clk (.A(clknet_5_16_0_clk),
    .X(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_clk (.A(clknet_5_16_0_clk),
    .X(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_clk (.A(clknet_5_16_0_clk),
    .X(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_clk (.A(clknet_5_16_0_clk),
    .X(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_clk (.A(clknet_5_17_0_clk),
    .X(clknet_leaf_28_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_clk (.A(clknet_5_17_0_clk),
    .X(clknet_leaf_29_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_clk (.A(clknet_5_17_0_clk),
    .X(clknet_leaf_30_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_clk (.A(clknet_5_17_0_clk),
    .X(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_clk (.A(clknet_5_17_0_clk),
    .X(clknet_leaf_32_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_clk (.A(clknet_5_17_0_clk),
    .X(clknet_leaf_33_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_clk (.A(clknet_5_17_0_clk),
    .X(clknet_leaf_34_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_clk (.A(clknet_5_17_0_clk),
    .X(clknet_leaf_35_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_clk (.A(clknet_5_17_0_clk),
    .X(clknet_leaf_36_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_clk (.A(clknet_5_18_0_clk),
    .X(clknet_leaf_37_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_clk (.A(clknet_5_18_0_clk),
    .X(clknet_leaf_38_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_clk (.A(clknet_5_18_0_clk),
    .X(clknet_leaf_39_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_clk (.A(clknet_opt_17_clk),
    .X(clknet_leaf_40_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_41_clk (.A(clknet_opt_18_clk),
    .X(clknet_leaf_41_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_42_clk (.A(clknet_opt_19_clk),
    .X(clknet_leaf_42_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_43_clk (.A(clknet_5_18_0_clk),
    .X(clknet_leaf_43_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_44_clk (.A(clknet_5_18_0_clk),
    .X(clknet_leaf_44_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_45_clk (.A(clknet_5_18_0_clk),
    .X(clknet_leaf_45_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_46_clk (.A(clknet_5_18_0_clk),
    .X(clknet_leaf_46_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_47_clk (.A(clknet_5_18_0_clk),
    .X(clknet_leaf_47_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_48_clk (.A(clknet_opt_32_clk),
    .X(clknet_leaf_48_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_49_clk (.A(clknet_5_30_0_clk),
    .X(clknet_leaf_49_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_50_clk (.A(clknet_5_30_0_clk),
    .X(clknet_leaf_50_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_51_clk (.A(clknet_5_31_0_clk),
    .X(clknet_leaf_51_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_52_clk (.A(clknet_5_31_0_clk),
    .X(clknet_leaf_52_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_53_clk (.A(clknet_5_31_0_clk),
    .X(clknet_leaf_53_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_54_clk (.A(clknet_5_19_0_clk),
    .X(clknet_leaf_54_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_55_clk (.A(clknet_5_18_0_clk),
    .X(clknet_leaf_55_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_56_clk (.A(clknet_opt_24_clk),
    .X(clknet_leaf_56_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_57_clk (.A(clknet_5_19_0_clk),
    .X(clknet_leaf_57_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_58_clk (.A(clknet_5_19_0_clk),
    .X(clknet_leaf_58_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_59_clk (.A(clknet_5_19_0_clk),
    .X(clknet_leaf_59_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_60_clk (.A(clknet_5_19_0_clk),
    .X(clknet_leaf_60_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_61_clk (.A(clknet_opt_25_clk),
    .X(clknet_leaf_61_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_67_clk (.A(clknet_5_17_0_clk),
    .X(clknet_leaf_67_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_68_clk (.A(clknet_opt_20_clk),
    .X(clknet_leaf_68_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_69_clk (.A(clknet_5_20_0_clk),
    .X(clknet_leaf_69_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_70_clk (.A(clknet_5_21_0_clk),
    .X(clknet_leaf_70_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_71_clk (.A(clknet_5_21_0_clk),
    .X(clknet_leaf_71_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_74_clk (.A(clknet_opt_22_clk),
    .X(clknet_leaf_74_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_75_clk (.A(clknet_opt_23_clk),
    .X(clknet_leaf_75_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_76_clk (.A(clknet_5_21_0_clk),
    .X(clknet_leaf_76_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_79_clk (.A(clknet_opt_29_clk),
    .X(clknet_leaf_79_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_82_clk (.A(clknet_5_22_0_clk),
    .X(clknet_leaf_82_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_83_clk (.A(clknet_5_22_0_clk),
    .X(clknet_leaf_83_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_84_clk (.A(clknet_5_5_0_clk),
    .X(clknet_leaf_84_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_87_clk (.A(clknet_5_5_0_clk),
    .X(clknet_leaf_87_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_89_clk (.A(clknet_opt_9_clk),
    .X(clknet_leaf_89_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_90_clk (.A(clknet_opt_10_clk),
    .X(clknet_leaf_90_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_91_clk (.A(clknet_opt_11_clk),
    .X(clknet_leaf_91_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_92_clk (.A(clknet_opt_3_clk),
    .X(clknet_leaf_92_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_94_clk (.A(clknet_opt_12_clk),
    .X(clknet_leaf_94_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_95_clk (.A(clknet_opt_13_clk),
    .X(clknet_leaf_95_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_103_clk (.A(clknet_opt_6_clk),
    .X(clknet_leaf_103_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_104_clk (.A(clknet_5_7_0_clk),
    .X(clknet_leaf_104_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_105_clk (.A(clknet_5_5_0_clk),
    .X(clknet_leaf_105_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_106_clk (.A(clknet_5_4_0_clk),
    .X(clknet_leaf_106_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_107_clk (.A(clknet_5_7_0_clk),
    .X(clknet_leaf_107_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_109_clk (.A(clknet_5_15_0_clk),
    .X(clknet_leaf_109_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_111_clk (.A(clknet_5_15_0_clk),
    .X(clknet_leaf_111_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_112_clk (.A(clknet_5_15_0_clk),
    .X(clknet_leaf_112_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_113_clk (.A(clknet_5_15_0_clk),
    .X(clknet_leaf_113_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_115_clk (.A(clknet_5_14_0_clk),
    .X(clknet_leaf_115_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_116_clk (.A(clknet_5_14_0_clk),
    .X(clknet_leaf_116_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_117_clk (.A(clknet_5_14_0_clk),
    .X(clknet_leaf_117_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_118_clk (.A(clknet_5_14_0_clk),
    .X(clknet_leaf_118_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_120_clk (.A(clknet_5_14_0_clk),
    .X(clknet_leaf_120_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_121_clk (.A(clknet_5_15_0_clk),
    .X(clknet_leaf_121_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_122_clk (.A(clknet_5_15_0_clk),
    .X(clknet_leaf_122_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_123_clk (.A(clknet_5_12_0_clk),
    .X(clknet_leaf_123_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_124_clk (.A(clknet_opt_7_clk),
    .X(clknet_leaf_124_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_125_clk (.A(clknet_opt_8_clk),
    .X(clknet_leaf_125_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_126_clk (.A(clknet_5_11_0_clk),
    .X(clknet_leaf_126_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_127_clk (.A(clknet_5_11_0_clk),
    .X(clknet_leaf_127_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_128_clk (.A(clknet_5_11_0_clk),
    .X(clknet_leaf_128_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_129_clk (.A(clknet_5_11_0_clk),
    .X(clknet_leaf_129_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_130_clk (.A(clknet_5_11_0_clk),
    .X(clknet_leaf_130_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_131_clk (.A(clknet_5_11_0_clk),
    .X(clknet_leaf_131_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_132_clk (.A(clknet_5_11_0_clk),
    .X(clknet_leaf_132_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_133_clk (.A(clknet_5_11_0_clk),
    .X(clknet_leaf_133_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_135_clk (.A(clknet_5_9_0_clk),
    .X(clknet_leaf_135_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_136_clk (.A(clknet_5_11_0_clk),
    .X(clknet_leaf_136_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_137_clk (.A(clknet_5_11_0_clk),
    .X(clknet_leaf_137_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_138_clk (.A(clknet_5_9_0_clk),
    .X(clknet_leaf_138_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_139_clk (.A(clknet_5_9_0_clk),
    .X(clknet_leaf_139_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_140_clk (.A(clknet_5_10_0_clk),
    .X(clknet_leaf_140_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_141_clk (.A(clknet_5_10_0_clk),
    .X(clknet_leaf_141_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_142_clk (.A(clknet_5_10_0_clk),
    .X(clknet_leaf_142_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_143_clk (.A(clknet_5_10_0_clk),
    .X(clknet_leaf_143_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_144_clk (.A(clknet_5_10_0_clk),
    .X(clknet_leaf_144_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_145_clk (.A(clknet_5_10_0_clk),
    .X(clknet_leaf_145_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_146_clk (.A(clknet_5_8_0_clk),
    .X(clknet_leaf_146_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_147_clk (.A(clknet_5_10_0_clk),
    .X(clknet_leaf_147_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_148_clk (.A(clknet_5_10_0_clk),
    .X(clknet_leaf_148_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_149_clk (.A(clknet_5_8_0_clk),
    .X(clknet_leaf_149_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_150_clk (.A(clknet_5_8_0_clk),
    .X(clknet_leaf_150_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_151_clk (.A(clknet_5_8_0_clk),
    .X(clknet_leaf_151_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_152_clk (.A(clknet_5_8_0_clk),
    .X(clknet_leaf_152_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_153_clk (.A(clknet_5_8_0_clk),
    .X(clknet_leaf_153_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_154_clk (.A(clknet_5_8_0_clk),
    .X(clknet_leaf_154_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_155_clk (.A(clknet_5_8_0_clk),
    .X(clknet_leaf_155_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_156_clk (.A(clknet_5_8_0_clk),
    .X(clknet_leaf_156_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_157_clk (.A(clknet_5_8_0_clk),
    .X(clknet_leaf_157_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_158_clk (.A(clknet_5_9_0_clk),
    .X(clknet_leaf_158_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_159_clk (.A(clknet_5_8_0_clk),
    .X(clknet_leaf_159_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_160_clk (.A(clknet_5_8_0_clk),
    .X(clknet_leaf_160_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_161_clk (.A(clknet_5_9_0_clk),
    .X(clknet_leaf_161_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_162_clk (.A(clknet_5_9_0_clk),
    .X(clknet_leaf_162_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_163_clk (.A(clknet_5_9_0_clk),
    .X(clknet_leaf_163_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_164_clk (.A(clknet_5_9_0_clk),
    .X(clknet_leaf_164_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_165_clk (.A(clknet_5_9_0_clk),
    .X(clknet_leaf_165_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_166_clk (.A(clknet_5_3_0_clk),
    .X(clknet_leaf_166_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_167_clk (.A(clknet_5_3_0_clk),
    .X(clknet_leaf_167_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_168_clk (.A(clknet_5_9_0_clk),
    .X(clknet_leaf_168_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_169_clk (.A(clknet_5_8_0_clk),
    .X(clknet_leaf_169_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_170_clk (.A(clknet_5_8_0_clk),
    .X(clknet_leaf_170_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_171_clk (.A(clknet_5_2_0_clk),
    .X(clknet_leaf_171_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_172_clk (.A(clknet_5_2_0_clk),
    .X(clknet_leaf_172_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_173_clk (.A(clknet_5_2_0_clk),
    .X(clknet_leaf_173_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_174_clk (.A(clknet_5_2_0_clk),
    .X(clknet_leaf_174_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_175_clk (.A(clknet_5_3_0_clk),
    .X(clknet_leaf_175_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_176_clk (.A(clknet_5_2_0_clk),
    .X(clknet_leaf_176_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_177_clk (.A(clknet_5_2_0_clk),
    .X(clknet_leaf_177_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_178_clk (.A(clknet_5_2_0_clk),
    .X(clknet_leaf_178_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_179_clk (.A(clknet_5_0_0_clk),
    .X(clknet_leaf_179_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_180_clk (.A(clknet_5_0_0_clk),
    .X(clknet_leaf_180_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_181_clk (.A(clknet_5_0_0_clk),
    .X(clknet_leaf_181_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_182_clk (.A(clknet_5_1_0_clk),
    .X(clknet_leaf_182_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_183_clk (.A(clknet_5_1_0_clk),
    .X(clknet_leaf_183_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_184_clk (.A(clknet_5_3_0_clk),
    .X(clknet_leaf_184_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_185_clk (.A(clknet_5_1_0_clk),
    .X(clknet_leaf_185_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_186_clk (.A(clknet_5_1_0_clk),
    .X(clknet_leaf_186_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_187_clk (.A(clknet_5_4_0_clk),
    .X(clknet_leaf_187_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_188_clk (.A(clknet_5_3_0_clk),
    .X(clknet_leaf_188_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_189_clk (.A(clknet_5_3_0_clk),
    .X(clknet_leaf_189_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_190_clk (.A(clknet_5_3_0_clk),
    .X(clknet_leaf_190_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_191_clk (.A(clknet_5_3_0_clk),
    .X(clknet_leaf_191_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_192_clk (.A(clknet_5_3_0_clk),
    .X(clknet_leaf_192_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_194_clk (.A(clknet_5_6_0_clk),
    .X(clknet_leaf_194_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_195_clk (.A(clknet_5_14_0_clk),
    .X(clknet_leaf_195_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_196_clk (.A(clknet_5_15_0_clk),
    .X(clknet_leaf_196_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_197_clk (.A(clknet_5_6_0_clk),
    .X(clknet_leaf_197_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_198_clk (.A(clknet_5_6_0_clk),
    .X(clknet_leaf_198_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_199_clk (.A(clknet_5_6_0_clk),
    .X(clknet_leaf_199_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_200_clk (.A(clknet_5_4_0_clk),
    .X(clknet_leaf_200_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_201_clk (.A(clknet_5_4_0_clk),
    .X(clknet_leaf_201_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_202_clk (.A(clknet_5_4_0_clk),
    .X(clknet_leaf_202_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_203_clk (.A(clknet_5_6_0_clk),
    .X(clknet_leaf_203_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_204_clk (.A(clknet_5_6_0_clk),
    .X(clknet_leaf_204_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_205_clk (.A(clknet_5_4_0_clk),
    .X(clknet_leaf_205_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_206_clk (.A(clknet_5_4_0_clk),
    .X(clknet_leaf_206_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_207_clk (.A(clknet_5_4_0_clk),
    .X(clknet_leaf_207_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_208_clk (.A(clknet_5_5_0_clk),
    .X(clknet_leaf_208_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_209_clk (.A(clknet_5_19_0_clk),
    .X(clknet_leaf_209_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_210_clk (.A(clknet_5_31_0_clk),
    .X(clknet_leaf_210_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_211_clk (.A(clknet_5_19_0_clk),
    .X(clknet_leaf_211_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_212_clk (.A(clknet_5_31_0_clk),
    .X(clknet_leaf_212_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_213_clk (.A(clknet_5_31_0_clk),
    .X(clknet_leaf_213_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_214_clk (.A(clknet_5_4_0_clk),
    .X(clknet_leaf_214_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_215_clk (.A(clknet_5_30_0_clk),
    .X(clknet_leaf_215_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_216_clk (.A(clknet_5_30_0_clk),
    .X(clknet_leaf_216_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_217_clk (.A(clknet_5_30_0_clk),
    .X(clknet_leaf_217_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_219_clk (.A(clknet_5_30_0_clk),
    .X(clknet_leaf_219_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_220_clk (.A(clknet_5_30_0_clk),
    .X(clknet_leaf_220_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_221_clk (.A(clknet_5_30_0_clk),
    .X(clknet_leaf_221_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_222_clk (.A(clknet_5_29_0_clk),
    .X(clknet_leaf_222_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_223_clk (.A(clknet_5_29_0_clk),
    .X(clknet_leaf_223_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_224_clk (.A(clknet_5_29_0_clk),
    .X(clknet_leaf_224_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_225_clk (.A(clknet_5_29_0_clk),
    .X(clknet_leaf_225_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_226_clk (.A(clknet_5_28_0_clk),
    .X(clknet_leaf_226_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_227_clk (.A(clknet_5_29_0_clk),
    .X(clknet_leaf_227_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_228_clk (.A(clknet_5_29_0_clk),
    .X(clknet_leaf_228_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_229_clk (.A(clknet_5_1_0_clk),
    .X(clknet_leaf_229_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_230_clk (.A(clknet_5_1_0_clk),
    .X(clknet_leaf_230_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_231_clk (.A(clknet_5_28_0_clk),
    .X(clknet_leaf_231_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_233_clk (.A(clknet_5_28_0_clk),
    .X(clknet_leaf_233_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_234_clk (.A(clknet_5_0_0_clk),
    .X(clknet_leaf_234_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_235_clk (.A(clknet_5_0_0_clk),
    .X(clknet_leaf_235_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_236_clk (.A(clknet_5_28_0_clk),
    .X(clknet_leaf_236_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_237_clk (.A(clknet_5_28_0_clk),
    .X(clknet_leaf_237_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_238_clk (.A(clknet_5_28_0_clk),
    .X(clknet_leaf_238_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_239_clk (.A(clknet_5_26_0_clk),
    .X(clknet_leaf_239_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_240_clk (.A(clknet_5_26_0_clk),
    .X(clknet_leaf_240_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_241_clk (.A(clknet_5_26_0_clk),
    .X(clknet_leaf_241_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_242_clk (.A(clknet_5_26_0_clk),
    .X(clknet_leaf_242_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_243_clk (.A(clknet_5_26_0_clk),
    .X(clknet_leaf_243_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_244_clk (.A(clknet_5_26_0_clk),
    .X(clknet_leaf_244_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_245_clk (.A(clknet_5_27_0_clk),
    .X(clknet_leaf_245_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_246_clk (.A(clknet_5_27_0_clk),
    .X(clknet_leaf_246_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_247_clk (.A(clknet_5_29_0_clk),
    .X(clknet_leaf_247_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_248_clk (.A(clknet_5_29_0_clk),
    .X(clknet_leaf_248_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_249_clk (.A(clknet_5_27_0_clk),
    .X(clknet_leaf_249_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_250_clk (.A(clknet_5_27_0_clk),
    .X(clknet_leaf_250_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_251_clk (.A(clknet_5_27_0_clk),
    .X(clknet_leaf_251_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_252_clk (.A(clknet_5_27_0_clk),
    .X(clknet_leaf_252_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_253_clk (.A(clknet_5_25_0_clk),
    .X(clknet_leaf_253_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_254_clk (.A(clknet_5_24_0_clk),
    .X(clknet_leaf_254_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_255_clk (.A(clknet_5_27_0_clk),
    .X(clknet_leaf_255_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_256_clk (.A(clknet_5_27_0_clk),
    .X(clknet_leaf_256_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_257_clk (.A(clknet_5_26_0_clk),
    .X(clknet_leaf_257_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_258_clk (.A(clknet_5_26_0_clk),
    .X(clknet_leaf_258_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_259_clk (.A(clknet_5_26_0_clk),
    .X(clknet_leaf_259_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_260_clk (.A(clknet_5_26_0_clk),
    .X(clknet_leaf_260_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_261_clk (.A(clknet_5_24_0_clk),
    .X(clknet_leaf_261_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_262_clk (.A(clknet_5_24_0_clk),
    .X(clknet_leaf_262_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_263_clk (.A(clknet_5_24_0_clk),
    .X(clknet_leaf_263_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_264_clk (.A(clknet_5_24_0_clk),
    .X(clknet_leaf_264_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_265_clk (.A(clknet_5_24_0_clk),
    .X(clknet_leaf_265_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_266_clk (.A(clknet_5_24_0_clk),
    .X(clknet_leaf_266_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_267_clk (.A(clknet_5_24_0_clk),
    .X(clknet_leaf_267_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_268_clk (.A(clknet_5_24_0_clk),
    .X(clknet_leaf_268_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_269_clk (.A(clknet_5_24_0_clk),
    .X(clknet_leaf_269_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_1_0_0_clk (.A(clknet_0_clk),
    .X(clknet_1_0_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_1_0_1_clk (.A(clknet_1_0_0_clk),
    .X(clknet_1_0_1_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_1_1_0_clk (.A(clknet_0_clk),
    .X(clknet_1_1_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_1_1_1_clk (.A(clknet_1_1_0_clk),
    .X(clknet_1_1_1_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_2_0_0_clk (.A(clknet_1_0_1_clk),
    .X(clknet_2_0_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_2_0_1_clk (.A(clknet_2_0_0_clk),
    .X(clknet_2_0_1_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_2_1_0_clk (.A(clknet_1_0_1_clk),
    .X(clknet_2_1_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_2_1_1_clk (.A(clknet_2_1_0_clk),
    .X(clknet_2_1_1_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_2_2_0_clk (.A(clknet_1_1_1_clk),
    .X(clknet_2_2_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_2_2_1_clk (.A(clknet_2_2_0_clk),
    .X(clknet_2_2_1_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_2_3_0_clk (.A(clknet_1_1_1_clk),
    .X(clknet_2_3_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_2_3_1_clk (.A(clknet_2_3_0_clk),
    .X(clknet_2_3_1_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_3_0_0_clk (.A(clknet_2_0_1_clk),
    .X(clknet_3_0_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_3_1_0_clk (.A(clknet_2_0_1_clk),
    .X(clknet_3_1_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_3_2_0_clk (.A(clknet_2_1_1_clk),
    .X(clknet_3_2_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_3_3_0_clk (.A(clknet_2_1_1_clk),
    .X(clknet_3_3_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_3_4_0_clk (.A(clknet_2_2_1_clk),
    .X(clknet_3_4_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_3_5_0_clk (.A(clknet_2_2_1_clk),
    .X(clknet_3_5_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_3_6_0_clk (.A(clknet_2_3_1_clk),
    .X(clknet_3_6_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_3_7_0_clk (.A(clknet_2_3_1_clk),
    .X(clknet_3_7_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_0_0_clk (.A(clknet_3_0_0_clk),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_1_0_clk (.A(clknet_3_0_0_clk),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_2_0_clk (.A(clknet_3_1_0_clk),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_3_0_clk (.A(clknet_3_1_0_clk),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_4_0_clk (.A(clknet_3_2_0_clk),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_5_0_clk (.A(clknet_3_2_0_clk),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_6_0_clk (.A(clknet_3_3_0_clk),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_7_0_clk (.A(clknet_3_3_0_clk),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_8_0_clk (.A(clknet_3_4_0_clk),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_9_0_clk (.A(clknet_3_4_0_clk),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_10_0_clk (.A(clknet_3_5_0_clk),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_11_0_clk (.A(clknet_3_5_0_clk),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_12_0_clk (.A(clknet_3_6_0_clk),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_13_0_clk (.A(clknet_3_6_0_clk),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_14_0_clk (.A(clknet_3_7_0_clk),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_15_0_clk (.A(clknet_3_7_0_clk),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_0_0_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_0_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_1_0_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_1_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_2_0_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_2_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_3_0_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_3_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_4_0_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_4_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_5_0_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_5_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_6_0_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_6_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_7_0_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_7_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_8_0_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_8_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_9_0_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_9_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_10_0_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_10_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_11_0_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_11_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_12_0_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_12_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_13_0_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_13_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_14_0_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_14_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_15_0_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_15_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_16_0_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_16_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_17_0_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_17_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_18_0_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_18_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_19_0_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_19_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_20_0_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_20_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_21_0_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_21_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_22_0_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_22_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_23_0_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_23_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_24_0_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_24_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_25_0_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_25_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_26_0_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_26_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_27_0_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_27_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_28_0_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_28_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_29_0_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_29_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_30_0_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_30_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_31_0_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_31_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_0_clk (.A(clknet_5_5_0_clk),
    .X(clknet_opt_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_1_clk (.A(clknet_5_5_0_clk),
    .X(clknet_opt_1_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_2_clk (.A(clknet_5_7_0_clk),
    .X(clknet_opt_2_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_3_clk (.A(clknet_5_7_0_clk),
    .X(clknet_opt_3_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_4_clk (.A(clknet_5_12_0_clk),
    .X(clknet_opt_4_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_5_clk (.A(clknet_5_12_0_clk),
    .X(clknet_opt_5_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_6_clk (.A(clknet_5_12_0_clk),
    .X(clknet_opt_6_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_7_clk (.A(clknet_5_12_0_clk),
    .X(clknet_opt_7_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_8_clk (.A(clknet_5_12_0_clk),
    .X(clknet_opt_8_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_9_clk (.A(clknet_5_13_0_clk),
    .X(clknet_opt_9_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_10_clk (.A(clknet_5_13_0_clk),
    .X(clknet_opt_10_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_11_clk (.A(clknet_5_13_0_clk),
    .X(clknet_opt_11_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_12_clk (.A(clknet_5_13_0_clk),
    .X(clknet_opt_12_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_13_clk (.A(clknet_5_13_0_clk),
    .X(clknet_opt_13_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_14_clk (.A(clknet_5_13_0_clk),
    .X(clknet_opt_14_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_15_clk (.A(clknet_5_13_0_clk),
    .X(clknet_opt_15_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_16_clk (.A(clknet_5_13_0_clk),
    .X(clknet_opt_16_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_17_clk (.A(clknet_5_20_0_clk),
    .X(clknet_opt_17_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_18_clk (.A(clknet_5_20_0_clk),
    .X(clknet_opt_18_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_19_clk (.A(clknet_5_20_0_clk),
    .X(clknet_opt_19_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_20_clk (.A(clknet_5_20_0_clk),
    .X(clknet_opt_20_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_21_clk (.A(clknet_5_21_0_clk),
    .X(clknet_opt_21_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_22_clk (.A(clknet_5_21_0_clk),
    .X(clknet_opt_22_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_23_clk (.A(clknet_5_21_0_clk),
    .X(clknet_opt_23_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_24_clk (.A(clknet_5_22_0_clk),
    .X(clknet_opt_24_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_25_clk (.A(clknet_5_22_0_clk),
    .X(clknet_opt_25_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_26_clk (.A(clknet_5_22_0_clk),
    .X(clknet_opt_26_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_27_clk (.A(clknet_5_23_0_clk),
    .X(clknet_opt_27_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_28_clk (.A(clknet_5_23_0_clk),
    .X(clknet_opt_28_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_29_clk (.A(clknet_5_23_0_clk),
    .X(clknet_opt_29_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_30_clk (.A(clknet_5_23_0_clk),
    .X(clknet_opt_30_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_31_clk (.A(clknet_5_25_0_clk),
    .X(clknet_opt_31_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_32_clk (.A(clknet_5_27_0_clk),
    .X(clknet_opt_32_clk));
endmodule
